# Copyright (c) 1993 - 2021 ARM Limited. All Rights Reserved.
# Use of this Software is subject to the terms and conditions of the
# applicable license agreement with ARM Limited.

# PhyVGen V 8.17.0
# ARM Version r0p0
# Creation Date: Tue Apr 27 11:33:11 2021


# Memory Configuration:
# ~~~~~~~~~~~~~~~~~~~~~
#  -activity_factor 50 -atf off -back_biasing off -bits 32 -bmux off
# -bus_notation on -c4obs off -check_instname off -diodes on -drive 6 -ema on
# -eol_guardband 0 -flexible_banking 4 -flexible_slice 2 -frequency 1.0
# -instname gf12lp_1rw_lg12_w32_bit -left_bus_delim "[" -lren_bankmask off -mux
# 4 -mvt BASE -name_case upper -pipeline off -power_gating off -power_type otc
# -prefix "" -pwr_gnd_rename vddpe:VDDPE,vddce:VDDCE,vsse:VSSE -rcols 2
# -redundancy off -retention on -right_bus_delim "]" -rrows 0 -scan off -ser
# none -site_def off -top_layer m5-m10 -vmin_assist off -words 4096 -write_mask
# on -write_thru off -corners
# ffpg_sigcmin_0p88v_0p88v_m40c,sspg_sigcmax_0p72v_0p72v_125c,tt_nominal_0p80v_0p80v_25c
# 

VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO gf12lp_1rw_lg12_w32_bit
	FOREIGN gf12lp_1rw_lg12_w32_bit 0 0 ;
	SYMMETRY X Y ;
	SIZE 201.665 BY 82.176 ;
	CLASS BLOCK ;
	PIN A[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 44.197 0.18 44.267 ;
			LAYER	M2 ;
			RECT	0 44.196 0.134 44.268 ;
			LAYER	M3 ;
			RECT	0 44.196 0.134 44.268 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END A[0]

	PIN A[10]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 42.037 0.18 42.107 ;
			LAYER	M2 ;
			RECT	0 42.036 0.134 42.108 ;
			LAYER	M3 ;
			RECT	0 42.036 0.134 42.108 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END A[10]

	PIN A[11]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 43.717 0.18 43.787 ;
			LAYER	M2 ;
			RECT	0 43.716 0.134 43.788 ;
			LAYER	M3 ;
			RECT	0 43.716 0.134 43.788 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END A[11]

	PIN A[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 45.061 0.18 45.131 ;
			LAYER	M2 ;
			RECT	0 45.06 0.134 45.132 ;
			LAYER	M3 ;
			RECT	0 45.06 0.134 45.132 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END A[1]

	PIN A[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 37.525 0.18 37.595 ;
			LAYER	M2 ;
			RECT	0 37.524 0.134 37.596 ;
			LAYER	M3 ;
			RECT	0 37.524 0.134 37.596 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END A[2]

	PIN A[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 35.605 0.18 35.675 ;
			LAYER	M2 ;
			RECT	0 35.604 0.134 35.676 ;
			LAYER	M3 ;
			RECT	0 35.604 0.134 35.676 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END A[3]

	PIN A[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 35.749 0.18 35.819 ;
			LAYER	M2 ;
			RECT	0 35.748 0.134 35.82 ;
			LAYER	M3 ;
			RECT	0 35.748 0.134 35.82 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END A[4]

	PIN A[5]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 39.445 0.18 39.515 ;
			LAYER	M2 ;
			RECT	0 39.444 0.134 39.516 ;
			LAYER	M3 ;
			RECT	0 39.444 0.134 39.516 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END A[5]

	PIN A[6]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 39.253 0.18 39.323 ;
			LAYER	M2 ;
			RECT	0 39.252 0.134 39.324 ;
			LAYER	M3 ;
			RECT	0 39.252 0.134 39.324 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END A[6]

	PIN A[7]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 38.005 0.18 38.075 ;
			LAYER	M2 ;
			RECT	0 38.004 0.134 38.076 ;
			LAYER	M3 ;
			RECT	0 38.004 0.134 38.076 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END A[7]

	PIN A[8]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 40.549 0.18 40.619 ;
			LAYER	M2 ;
			RECT	0 40.548 0.134 40.62 ;
			LAYER	M3 ;
			RECT	0 40.548 0.134 40.62 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END A[8]

	PIN A[9]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 41.029 0.18 41.099 ;
			LAYER	M2 ;
			RECT	0 41.028 0.134 41.1 ;
			LAYER	M3 ;
			RECT	0 41.028 0.134 41.1 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END A[9]

	PIN CEN
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 33.973 0.18 34.043 ;
			LAYER	M2 ;
			RECT	0 33.972 0.134 34.044 ;
			LAYER	M3 ;
			RECT	0 33.972 0.134 34.044 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END CEN

	PIN CLK
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 37.333 0.18 37.403 ;
			LAYER	M2 ;
			RECT	0 37.332 0.134 37.404 ;
			LAYER	M3 ;
			RECT	0 37.332 0.134 37.404 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END CLK

	PIN D[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 0.949 0.18 1.019 ;
			LAYER	M2 ;
			RECT	0 0.948 0.134 1.02 ;
			LAYER	M3 ;
			RECT	0 0.948 0.134 1.02 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[0]

	PIN D[10]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 20.149 0.18 20.219 ;
			LAYER	M2 ;
			RECT	0 20.148 0.134 20.22 ;
			LAYER	M3 ;
			RECT	0 20.148 0.134 20.22 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[10]

	PIN D[11]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 22.069 0.18 22.139 ;
			LAYER	M2 ;
			RECT	0 22.068 0.134 22.14 ;
			LAYER	M3 ;
			RECT	0 22.068 0.134 22.14 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[11]

	PIN D[12]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 23.989 0.18 24.059 ;
			LAYER	M2 ;
			RECT	0 23.988 0.134 24.06 ;
			LAYER	M3 ;
			RECT	0 23.988 0.134 24.06 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[12]

	PIN D[13]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 25.909 0.18 25.979 ;
			LAYER	M2 ;
			RECT	0 25.908 0.134 25.98 ;
			LAYER	M3 ;
			RECT	0 25.908 0.134 25.98 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[13]

	PIN D[14]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 27.829 0.18 27.899 ;
			LAYER	M2 ;
			RECT	0 27.828 0.134 27.9 ;
			LAYER	M3 ;
			RECT	0 27.828 0.134 27.9 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[14]

	PIN D[15]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 29.749 0.18 29.819 ;
			LAYER	M2 ;
			RECT	0 29.748 0.134 29.82 ;
			LAYER	M3 ;
			RECT	0 29.748 0.134 29.82 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[15]

	PIN D[16]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 52.357 0.18 52.427 ;
			LAYER	M2 ;
			RECT	0 52.356 0.134 52.428 ;
			LAYER	M3 ;
			RECT	0 52.356 0.134 52.428 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[16]

	PIN D[17]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 54.277 0.18 54.347 ;
			LAYER	M2 ;
			RECT	0 54.276 0.134 54.348 ;
			LAYER	M3 ;
			RECT	0 54.276 0.134 54.348 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[17]

	PIN D[18]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 56.197 0.18 56.267 ;
			LAYER	M2 ;
			RECT	0 56.196 0.134 56.268 ;
			LAYER	M3 ;
			RECT	0 56.196 0.134 56.268 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[18]

	PIN D[19]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 58.117 0.18 58.187 ;
			LAYER	M2 ;
			RECT	0 58.116 0.134 58.188 ;
			LAYER	M3 ;
			RECT	0 58.116 0.134 58.188 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[19]

	PIN D[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 2.869 0.18 2.939 ;
			LAYER	M2 ;
			RECT	0 2.868 0.134 2.94 ;
			LAYER	M3 ;
			RECT	0 2.868 0.134 2.94 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[1]

	PIN D[20]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 60.037 0.18 60.107 ;
			LAYER	M2 ;
			RECT	0 60.036 0.134 60.108 ;
			LAYER	M3 ;
			RECT	0 60.036 0.134 60.108 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[20]

	PIN D[21]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 61.957 0.18 62.027 ;
			LAYER	M2 ;
			RECT	0 61.956 0.134 62.028 ;
			LAYER	M3 ;
			RECT	0 61.956 0.134 62.028 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[21]

	PIN D[22]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 63.877 0.18 63.947 ;
			LAYER	M2 ;
			RECT	0 63.876 0.134 63.948 ;
			LAYER	M3 ;
			RECT	0 63.876 0.134 63.948 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[22]

	PIN D[23]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 65.797 0.18 65.867 ;
			LAYER	M2 ;
			RECT	0 65.796 0.134 65.868 ;
			LAYER	M3 ;
			RECT	0 65.796 0.134 65.868 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[23]

	PIN D[24]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 67.717 0.18 67.787 ;
			LAYER	M2 ;
			RECT	0 67.716 0.134 67.788 ;
			LAYER	M3 ;
			RECT	0 67.716 0.134 67.788 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[24]

	PIN D[25]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 69.637 0.18 69.707 ;
			LAYER	M2 ;
			RECT	0 69.636 0.134 69.708 ;
			LAYER	M3 ;
			RECT	0 69.636 0.134 69.708 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[25]

	PIN D[26]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 71.557 0.18 71.627 ;
			LAYER	M2 ;
			RECT	0 71.556 0.134 71.628 ;
			LAYER	M3 ;
			RECT	0 71.556 0.134 71.628 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[26]

	PIN D[27]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 73.477 0.18 73.547 ;
			LAYER	M2 ;
			RECT	0 73.476 0.134 73.548 ;
			LAYER	M3 ;
			RECT	0 73.476 0.134 73.548 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[27]

	PIN D[28]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 75.397 0.18 75.467 ;
			LAYER	M2 ;
			RECT	0 75.396 0.134 75.468 ;
			LAYER	M3 ;
			RECT	0 75.396 0.134 75.468 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[28]

	PIN D[29]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 77.317 0.18 77.387 ;
			LAYER	M2 ;
			RECT	0 77.316 0.134 77.388 ;
			LAYER	M3 ;
			RECT	0 77.316 0.134 77.388 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[29]

	PIN D[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 4.789 0.18 4.859 ;
			LAYER	M2 ;
			RECT	0 4.788 0.134 4.86 ;
			LAYER	M3 ;
			RECT	0 4.788 0.134 4.86 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[2]

	PIN D[30]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 79.237 0.18 79.307 ;
			LAYER	M2 ;
			RECT	0 79.236 0.134 79.308 ;
			LAYER	M3 ;
			RECT	0 79.236 0.134 79.308 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[30]

	PIN D[31]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 81.157 0.18 81.227 ;
			LAYER	M2 ;
			RECT	0 81.156 0.134 81.228 ;
			LAYER	M3 ;
			RECT	0 81.156 0.134 81.228 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[31]

	PIN D[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 6.709 0.18 6.779 ;
			LAYER	M2 ;
			RECT	0 6.708 0.134 6.78 ;
			LAYER	M3 ;
			RECT	0 6.708 0.134 6.78 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[3]

	PIN D[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 8.629 0.18 8.699 ;
			LAYER	M2 ;
			RECT	0 8.628 0.134 8.7 ;
			LAYER	M3 ;
			RECT	0 8.628 0.134 8.7 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[4]

	PIN D[5]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 10.549 0.18 10.619 ;
			LAYER	M2 ;
			RECT	0 10.548 0.134 10.62 ;
			LAYER	M3 ;
			RECT	0 10.548 0.134 10.62 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[5]

	PIN D[6]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 12.469 0.18 12.539 ;
			LAYER	M2 ;
			RECT	0 12.468 0.134 12.54 ;
			LAYER	M3 ;
			RECT	0 12.468 0.134 12.54 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[6]

	PIN D[7]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 14.389 0.18 14.459 ;
			LAYER	M2 ;
			RECT	0 14.388 0.134 14.46 ;
			LAYER	M3 ;
			RECT	0 14.388 0.134 14.46 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[7]

	PIN D[8]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 16.309 0.18 16.379 ;
			LAYER	M2 ;
			RECT	0 16.308 0.134 16.38 ;
			LAYER	M3 ;
			RECT	0 16.308 0.134 16.38 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[8]

	PIN D[9]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 18.229 0.18 18.299 ;
			LAYER	M2 ;
			RECT	0 18.228 0.134 18.3 ;
			LAYER	M3 ;
			RECT	0 18.228 0.134 18.3 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END D[9]

	PIN EMAS
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 34.117 0.18 34.187 ;
			LAYER	M2 ;
			RECT	0 34.116 0.134 34.188 ;
			LAYER	M3 ;
			RECT	0 34.116 0.134 34.188 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END EMAS

	PIN EMAW[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 34.597 0.18 34.667 ;
			LAYER	M2 ;
			RECT	0 34.596 0.134 34.668 ;
			LAYER	M3 ;
			RECT	0 34.596 0.134 34.668 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END EMAW[0]

	PIN EMAW[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 34.309 0.18 34.379 ;
			LAYER	M2 ;
			RECT	0 34.308 0.134 34.38 ;
			LAYER	M3 ;
			RECT	0 34.308 0.134 34.38 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END EMAW[1]

	PIN EMA[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 42.229 0.18 42.299 ;
			LAYER	M2 ;
			RECT	0 42.228 0.134 42.3 ;
			LAYER	M3 ;
			RECT	0 42.228 0.134 42.3 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END EMA[0]

	PIN EMA[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 41.557 0.18 41.627 ;
			LAYER	M2 ;
			RECT	0 41.556 0.134 41.628 ;
			LAYER	M3 ;
			RECT	0 41.556 0.134 41.628 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END EMA[1]

	PIN EMA[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 39.925 0.18 39.995 ;
			LAYER	M2 ;
			RECT	0 39.924 0.134 39.996 ;
			LAYER	M3 ;
			RECT	0 39.924 0.134 39.996 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END EMA[2]

	PIN GWEN
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 35.269 0.18 35.339 ;
			LAYER	M2 ;
			RECT	0 35.268 0.134 35.34 ;
			LAYER	M3 ;
			RECT	0 35.268 0.134 35.34 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END GWEN

	PIN Q[0]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 1.432 0.18 1.502 ;
			LAYER	M2 ;
			RECT	0 1.431 0.134 1.503 ;
			LAYER	M3 ;
			RECT	0 1.431 0.134 1.503 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[0]

	PIN Q[10]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 20.632 0.18 20.702 ;
			LAYER	M2 ;
			RECT	0 20.631 0.134 20.703 ;
			LAYER	M3 ;
			RECT	0 20.631 0.134 20.703 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[10]

	PIN Q[11]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 22.552 0.18 22.622 ;
			LAYER	M2 ;
			RECT	0 22.551 0.134 22.623 ;
			LAYER	M3 ;
			RECT	0 22.551 0.134 22.623 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[11]

	PIN Q[12]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 24.472 0.18 24.542 ;
			LAYER	M2 ;
			RECT	0 24.471 0.134 24.543 ;
			LAYER	M3 ;
			RECT	0 24.471 0.134 24.543 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[12]

	PIN Q[13]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 26.392 0.18 26.462 ;
			LAYER	M2 ;
			RECT	0 26.391 0.134 26.463 ;
			LAYER	M3 ;
			RECT	0 26.391 0.134 26.463 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[13]

	PIN Q[14]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 28.312 0.18 28.382 ;
			LAYER	M2 ;
			RECT	0 28.311 0.134 28.383 ;
			LAYER	M3 ;
			RECT	0 28.311 0.134 28.383 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[14]

	PIN Q[15]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 30.232 0.18 30.302 ;
			LAYER	M2 ;
			RECT	0 30.231 0.134 30.303 ;
			LAYER	M3 ;
			RECT	0 30.231 0.134 30.303 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[15]

	PIN Q[16]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 51.874 0.18 51.944 ;
			LAYER	M2 ;
			RECT	0 51.873 0.134 51.945 ;
			LAYER	M3 ;
			RECT	0 51.873 0.134 51.945 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[16]

	PIN Q[17]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 53.794 0.18 53.864 ;
			LAYER	M2 ;
			RECT	0 53.793 0.134 53.865 ;
			LAYER	M3 ;
			RECT	0 53.793 0.134 53.865 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[17]

	PIN Q[18]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 55.714 0.18 55.784 ;
			LAYER	M2 ;
			RECT	0 55.713 0.134 55.785 ;
			LAYER	M3 ;
			RECT	0 55.713 0.134 55.785 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[18]

	PIN Q[19]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 57.634 0.18 57.704 ;
			LAYER	M2 ;
			RECT	0 57.633 0.134 57.705 ;
			LAYER	M3 ;
			RECT	0 57.633 0.134 57.705 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[19]

	PIN Q[1]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 3.352 0.18 3.422 ;
			LAYER	M2 ;
			RECT	0 3.351 0.134 3.423 ;
			LAYER	M3 ;
			RECT	0 3.351 0.134 3.423 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[1]

	PIN Q[20]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 59.554 0.18 59.624 ;
			LAYER	M2 ;
			RECT	0 59.553 0.134 59.625 ;
			LAYER	M3 ;
			RECT	0 59.553 0.134 59.625 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[20]

	PIN Q[21]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 61.474 0.18 61.544 ;
			LAYER	M2 ;
			RECT	0 61.473 0.134 61.545 ;
			LAYER	M3 ;
			RECT	0 61.473 0.134 61.545 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[21]

	PIN Q[22]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 63.394 0.18 63.464 ;
			LAYER	M2 ;
			RECT	0 63.393 0.134 63.465 ;
			LAYER	M3 ;
			RECT	0 63.393 0.134 63.465 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[22]

	PIN Q[23]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 65.314 0.18 65.384 ;
			LAYER	M2 ;
			RECT	0 65.313 0.134 65.385 ;
			LAYER	M3 ;
			RECT	0 65.313 0.134 65.385 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[23]

	PIN Q[24]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 67.234 0.18 67.304 ;
			LAYER	M2 ;
			RECT	0 67.233 0.134 67.305 ;
			LAYER	M3 ;
			RECT	0 67.233 0.134 67.305 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[24]

	PIN Q[25]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 69.154 0.18 69.224 ;
			LAYER	M2 ;
			RECT	0 69.153 0.134 69.225 ;
			LAYER	M3 ;
			RECT	0 69.153 0.134 69.225 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[25]

	PIN Q[26]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 71.074 0.18 71.144 ;
			LAYER	M2 ;
			RECT	0 71.073 0.134 71.145 ;
			LAYER	M3 ;
			RECT	0 71.073 0.134 71.145 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[26]

	PIN Q[27]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 72.994 0.18 73.064 ;
			LAYER	M2 ;
			RECT	0 72.993 0.134 73.065 ;
			LAYER	M3 ;
			RECT	0 72.993 0.134 73.065 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[27]

	PIN Q[28]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 74.914 0.18 74.984 ;
			LAYER	M2 ;
			RECT	0 74.913 0.134 74.985 ;
			LAYER	M3 ;
			RECT	0 74.913 0.134 74.985 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[28]

	PIN Q[29]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 76.834 0.18 76.904 ;
			LAYER	M2 ;
			RECT	0 76.833 0.134 76.905 ;
			LAYER	M3 ;
			RECT	0 76.833 0.134 76.905 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[29]

	PIN Q[2]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 5.272 0.18 5.342 ;
			LAYER	M2 ;
			RECT	0 5.271 0.134 5.343 ;
			LAYER	M3 ;
			RECT	0 5.271 0.134 5.343 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[2]

	PIN Q[30]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 78.754 0.18 78.824 ;
			LAYER	M2 ;
			RECT	0 78.753 0.134 78.825 ;
			LAYER	M3 ;
			RECT	0 78.753 0.134 78.825 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[30]

	PIN Q[31]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 80.674 0.18 80.744 ;
			LAYER	M2 ;
			RECT	0 80.673 0.134 80.745 ;
			LAYER	M3 ;
			RECT	0 80.673 0.134 80.745 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[31]

	PIN Q[3]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 7.192 0.18 7.262 ;
			LAYER	M2 ;
			RECT	0 7.191 0.134 7.263 ;
			LAYER	M3 ;
			RECT	0 7.191 0.134 7.263 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[3]

	PIN Q[4]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 9.112 0.18 9.182 ;
			LAYER	M2 ;
			RECT	0 9.111 0.134 9.183 ;
			LAYER	M3 ;
			RECT	0 9.111 0.134 9.183 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[4]

	PIN Q[5]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 11.032 0.18 11.102 ;
			LAYER	M2 ;
			RECT	0 11.031 0.134 11.103 ;
			LAYER	M3 ;
			RECT	0 11.031 0.134 11.103 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[5]

	PIN Q[6]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 12.952 0.18 13.022 ;
			LAYER	M2 ;
			RECT	0 12.951 0.134 13.023 ;
			LAYER	M3 ;
			RECT	0 12.951 0.134 13.023 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[6]

	PIN Q[7]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 14.872 0.18 14.942 ;
			LAYER	M2 ;
			RECT	0 14.871 0.134 14.943 ;
			LAYER	M3 ;
			RECT	0 14.871 0.134 14.943 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[7]

	PIN Q[8]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 16.792 0.18 16.862 ;
			LAYER	M2 ;
			RECT	0 16.791 0.134 16.863 ;
			LAYER	M3 ;
			RECT	0 16.791 0.134 16.863 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[8]

	PIN Q[9]
		USE SIGNAL ;
		DIRECTION OUTPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 18.712 0.18 18.782 ;
			LAYER	M2 ;
			RECT	0 18.711 0.134 18.783 ;
			LAYER	M3 ;
			RECT	0 18.711 0.134 18.783 ;
		END

		ANTENNADIFFAREA 0.00252 ;
	END Q[9]

	PIN RET1N
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 47.605 0.18 47.675 ;
			LAYER	M2 ;
			RECT	0 47.604 0.134 47.676 ;
			LAYER	M3 ;
			RECT	0 47.604 0.134 47.676 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END RET1N

	PIN STOV
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 35.125 0.18 35.195 ;
			LAYER	M2 ;
			RECT	0 35.124 0.134 35.196 ;
			LAYER	M3 ;
			RECT	0 35.124 0.134 35.196 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END STOV

	PIN VDDCE
		USE POWER ;
		DIRECTION INOUT ;
		PORT
			LAYER	C4 ;
			RECT	0.294 80.816 201.665 80.926 ;
			LAYER	J3 ;
			RECT	5.514 80.839 5.578 80.903 ;
			RECT	5.675 80.839 5.707 80.903 ;
			RECT	49.691 80.839 49.723 80.903 ;
			RECT	49.82 80.839 49.884 80.903 ;
			RECT	58.32 80.839 58.384 80.903 ;
			RECT	58.481 80.839 58.513 80.903 ;
			RECT	102.497 80.839 102.529 80.903 ;
			RECT	102.626 80.839 102.69 80.903 ;
			RECT	103.512 80.839 103.576 80.903 ;
			RECT	103.673 80.839 103.705 80.903 ;
			RECT	147.689 80.839 147.721 80.903 ;
			RECT	147.818 80.839 147.882 80.903 ;
			RECT	156.318 80.839 156.382 80.903 ;
			RECT	156.479 80.839 156.511 80.903 ;
			RECT	200.495 80.839 200.527 80.903 ;
			RECT	200.624 80.839 200.688 80.903 ;
			RECT	201.14 80.855 201.204 80.887 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 76.976 201.665 77.086 ;
			LAYER	J3 ;
			RECT	5.514 76.999 5.578 77.063 ;
			RECT	5.675 76.999 5.707 77.063 ;
			RECT	49.691 76.999 49.723 77.063 ;
			RECT	49.82 76.999 49.884 77.063 ;
			RECT	58.32 76.999 58.384 77.063 ;
			RECT	58.481 76.999 58.513 77.063 ;
			RECT	102.497 76.999 102.529 77.063 ;
			RECT	102.626 76.999 102.69 77.063 ;
			RECT	103.512 76.999 103.576 77.063 ;
			RECT	103.673 76.999 103.705 77.063 ;
			RECT	147.689 76.999 147.721 77.063 ;
			RECT	147.818 76.999 147.882 77.063 ;
			RECT	156.318 76.999 156.382 77.063 ;
			RECT	156.479 76.999 156.511 77.063 ;
			RECT	200.495 76.999 200.527 77.063 ;
			RECT	200.624 76.999 200.688 77.063 ;
			RECT	201.14 77.015 201.204 77.047 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 30.05 201.665 30.16 ;
			LAYER	J3 ;
			RECT	5.514 30.073 5.578 30.137 ;
			RECT	5.675 30.073 5.707 30.137 ;
			RECT	49.691 30.073 49.723 30.137 ;
			RECT	49.82 30.073 49.884 30.137 ;
			RECT	58.32 30.073 58.384 30.137 ;
			RECT	58.481 30.073 58.513 30.137 ;
			RECT	102.497 30.073 102.529 30.137 ;
			RECT	102.626 30.073 102.69 30.137 ;
			RECT	103.512 30.073 103.576 30.137 ;
			RECT	103.673 30.073 103.705 30.137 ;
			RECT	147.689 30.073 147.721 30.137 ;
			RECT	147.818 30.073 147.882 30.137 ;
			RECT	156.318 30.073 156.382 30.137 ;
			RECT	156.479 30.073 156.511 30.137 ;
			RECT	200.495 30.073 200.527 30.137 ;
			RECT	200.624 30.073 200.688 30.137 ;
			RECT	201.14 30.089 201.204 30.121 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 28.13 201.665 28.24 ;
			LAYER	J3 ;
			RECT	5.514 28.153 5.578 28.217 ;
			RECT	5.675 28.153 5.707 28.217 ;
			RECT	49.691 28.153 49.723 28.217 ;
			RECT	49.82 28.153 49.884 28.217 ;
			RECT	58.32 28.153 58.384 28.217 ;
			RECT	58.481 28.153 58.513 28.217 ;
			RECT	102.497 28.153 102.529 28.217 ;
			RECT	102.626 28.153 102.69 28.217 ;
			RECT	103.512 28.153 103.576 28.217 ;
			RECT	103.673 28.153 103.705 28.217 ;
			RECT	147.689 28.153 147.721 28.217 ;
			RECT	147.818 28.153 147.882 28.217 ;
			RECT	156.318 28.153 156.382 28.217 ;
			RECT	156.479 28.153 156.511 28.217 ;
			RECT	200.495 28.153 200.527 28.217 ;
			RECT	200.624 28.153 200.688 28.217 ;
			RECT	201.14 28.169 201.204 28.201 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 26.21 201.665 26.32 ;
			LAYER	J3 ;
			RECT	5.514 26.233 5.578 26.297 ;
			RECT	5.675 26.233 5.707 26.297 ;
			RECT	49.691 26.233 49.723 26.297 ;
			RECT	49.82 26.233 49.884 26.297 ;
			RECT	58.32 26.233 58.384 26.297 ;
			RECT	58.481 26.233 58.513 26.297 ;
			RECT	102.497 26.233 102.529 26.297 ;
			RECT	102.626 26.233 102.69 26.297 ;
			RECT	103.512 26.233 103.576 26.297 ;
			RECT	103.673 26.233 103.705 26.297 ;
			RECT	147.689 26.233 147.721 26.297 ;
			RECT	147.818 26.233 147.882 26.297 ;
			RECT	156.318 26.233 156.382 26.297 ;
			RECT	156.479 26.233 156.511 26.297 ;
			RECT	200.495 26.233 200.527 26.297 ;
			RECT	200.624 26.233 200.688 26.297 ;
			RECT	201.14 26.249 201.204 26.281 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 24.29 201.665 24.4 ;
			LAYER	J3 ;
			RECT	5.514 24.313 5.578 24.377 ;
			RECT	5.675 24.313 5.707 24.377 ;
			RECT	49.691 24.313 49.723 24.377 ;
			RECT	49.82 24.313 49.884 24.377 ;
			RECT	58.32 24.313 58.384 24.377 ;
			RECT	58.481 24.313 58.513 24.377 ;
			RECT	102.497 24.313 102.529 24.377 ;
			RECT	102.626 24.313 102.69 24.377 ;
			RECT	103.512 24.313 103.576 24.377 ;
			RECT	103.673 24.313 103.705 24.377 ;
			RECT	147.689 24.313 147.721 24.377 ;
			RECT	147.818 24.313 147.882 24.377 ;
			RECT	156.318 24.313 156.382 24.377 ;
			RECT	156.479 24.313 156.511 24.377 ;
			RECT	200.495 24.313 200.527 24.377 ;
			RECT	200.624 24.313 200.688 24.377 ;
			RECT	201.14 24.329 201.204 24.361 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 22.37 201.665 22.48 ;
			LAYER	J3 ;
			RECT	5.514 22.393 5.578 22.457 ;
			RECT	5.675 22.393 5.707 22.457 ;
			RECT	49.691 22.393 49.723 22.457 ;
			RECT	49.82 22.393 49.884 22.457 ;
			RECT	58.32 22.393 58.384 22.457 ;
			RECT	58.481 22.393 58.513 22.457 ;
			RECT	102.497 22.393 102.529 22.457 ;
			RECT	102.626 22.393 102.69 22.457 ;
			RECT	103.512 22.393 103.576 22.457 ;
			RECT	103.673 22.393 103.705 22.457 ;
			RECT	147.689 22.393 147.721 22.457 ;
			RECT	147.818 22.393 147.882 22.457 ;
			RECT	156.318 22.393 156.382 22.457 ;
			RECT	156.479 22.393 156.511 22.457 ;
			RECT	200.495 22.393 200.527 22.457 ;
			RECT	200.624 22.393 200.688 22.457 ;
			RECT	201.14 22.409 201.204 22.441 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 20.45 201.665 20.56 ;
			LAYER	J3 ;
			RECT	5.514 20.473 5.578 20.537 ;
			RECT	5.675 20.473 5.707 20.537 ;
			RECT	49.691 20.473 49.723 20.537 ;
			RECT	49.82 20.473 49.884 20.537 ;
			RECT	58.32 20.473 58.384 20.537 ;
			RECT	58.481 20.473 58.513 20.537 ;
			RECT	102.497 20.473 102.529 20.537 ;
			RECT	102.626 20.473 102.69 20.537 ;
			RECT	103.512 20.473 103.576 20.537 ;
			RECT	103.673 20.473 103.705 20.537 ;
			RECT	147.689 20.473 147.721 20.537 ;
			RECT	147.818 20.473 147.882 20.537 ;
			RECT	156.318 20.473 156.382 20.537 ;
			RECT	156.479 20.473 156.511 20.537 ;
			RECT	200.495 20.473 200.527 20.537 ;
			RECT	200.624 20.473 200.688 20.537 ;
			RECT	201.14 20.489 201.204 20.521 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 18.53 201.665 18.64 ;
			LAYER	J3 ;
			RECT	5.514 18.553 5.578 18.617 ;
			RECT	5.675 18.553 5.707 18.617 ;
			RECT	49.691 18.553 49.723 18.617 ;
			RECT	49.82 18.553 49.884 18.617 ;
			RECT	58.32 18.553 58.384 18.617 ;
			RECT	58.481 18.553 58.513 18.617 ;
			RECT	102.497 18.553 102.529 18.617 ;
			RECT	102.626 18.553 102.69 18.617 ;
			RECT	103.512 18.553 103.576 18.617 ;
			RECT	103.673 18.553 103.705 18.617 ;
			RECT	147.689 18.553 147.721 18.617 ;
			RECT	147.818 18.553 147.882 18.617 ;
			RECT	156.318 18.553 156.382 18.617 ;
			RECT	156.479 18.553 156.511 18.617 ;
			RECT	200.495 18.553 200.527 18.617 ;
			RECT	200.624 18.553 200.688 18.617 ;
			RECT	201.14 18.569 201.204 18.601 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 16.61 201.665 16.72 ;
			LAYER	J3 ;
			RECT	5.514 16.633 5.578 16.697 ;
			RECT	5.675 16.633 5.707 16.697 ;
			RECT	49.691 16.633 49.723 16.697 ;
			RECT	49.82 16.633 49.884 16.697 ;
			RECT	58.32 16.633 58.384 16.697 ;
			RECT	58.481 16.633 58.513 16.697 ;
			RECT	102.497 16.633 102.529 16.697 ;
			RECT	102.626 16.633 102.69 16.697 ;
			RECT	103.512 16.633 103.576 16.697 ;
			RECT	103.673 16.633 103.705 16.697 ;
			RECT	147.689 16.633 147.721 16.697 ;
			RECT	147.818 16.633 147.882 16.697 ;
			RECT	156.318 16.633 156.382 16.697 ;
			RECT	156.479 16.633 156.511 16.697 ;
			RECT	200.495 16.633 200.527 16.697 ;
			RECT	200.624 16.633 200.688 16.697 ;
			RECT	201.14 16.649 201.204 16.681 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 14.69 201.665 14.8 ;
			LAYER	J3 ;
			RECT	5.514 14.713 5.578 14.777 ;
			RECT	5.675 14.713 5.707 14.777 ;
			RECT	49.691 14.713 49.723 14.777 ;
			RECT	49.82 14.713 49.884 14.777 ;
			RECT	58.32 14.713 58.384 14.777 ;
			RECT	58.481 14.713 58.513 14.777 ;
			RECT	102.497 14.713 102.529 14.777 ;
			RECT	102.626 14.713 102.69 14.777 ;
			RECT	103.512 14.713 103.576 14.777 ;
			RECT	103.673 14.713 103.705 14.777 ;
			RECT	147.689 14.713 147.721 14.777 ;
			RECT	147.818 14.713 147.882 14.777 ;
			RECT	156.318 14.713 156.382 14.777 ;
			RECT	156.479 14.713 156.511 14.777 ;
			RECT	200.495 14.713 200.527 14.777 ;
			RECT	200.624 14.713 200.688 14.777 ;
			RECT	201.14 14.729 201.204 14.761 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 12.77 201.665 12.88 ;
			LAYER	J3 ;
			RECT	5.514 12.793 5.578 12.857 ;
			RECT	5.675 12.793 5.707 12.857 ;
			RECT	49.691 12.793 49.723 12.857 ;
			RECT	49.82 12.793 49.884 12.857 ;
			RECT	58.32 12.793 58.384 12.857 ;
			RECT	58.481 12.793 58.513 12.857 ;
			RECT	102.497 12.793 102.529 12.857 ;
			RECT	102.626 12.793 102.69 12.857 ;
			RECT	103.512 12.793 103.576 12.857 ;
			RECT	103.673 12.793 103.705 12.857 ;
			RECT	147.689 12.793 147.721 12.857 ;
			RECT	147.818 12.793 147.882 12.857 ;
			RECT	156.318 12.793 156.382 12.857 ;
			RECT	156.479 12.793 156.511 12.857 ;
			RECT	200.495 12.793 200.527 12.857 ;
			RECT	200.624 12.793 200.688 12.857 ;
			RECT	201.14 12.809 201.204 12.841 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 75.056 201.665 75.166 ;
			LAYER	J3 ;
			RECT	5.514 75.079 5.578 75.143 ;
			RECT	5.675 75.079 5.707 75.143 ;
			RECT	49.691 75.079 49.723 75.143 ;
			RECT	49.82 75.079 49.884 75.143 ;
			RECT	58.32 75.079 58.384 75.143 ;
			RECT	58.481 75.079 58.513 75.143 ;
			RECT	102.497 75.079 102.529 75.143 ;
			RECT	102.626 75.079 102.69 75.143 ;
			RECT	103.512 75.079 103.576 75.143 ;
			RECT	103.673 75.079 103.705 75.143 ;
			RECT	147.689 75.079 147.721 75.143 ;
			RECT	147.818 75.079 147.882 75.143 ;
			RECT	156.318 75.079 156.382 75.143 ;
			RECT	156.479 75.079 156.511 75.143 ;
			RECT	200.495 75.079 200.527 75.143 ;
			RECT	200.624 75.079 200.688 75.143 ;
			RECT	201.14 75.095 201.204 75.127 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 10.85 201.665 10.96 ;
			LAYER	J3 ;
			RECT	5.514 10.873 5.578 10.937 ;
			RECT	5.675 10.873 5.707 10.937 ;
			RECT	49.691 10.873 49.723 10.937 ;
			RECT	49.82 10.873 49.884 10.937 ;
			RECT	58.32 10.873 58.384 10.937 ;
			RECT	58.481 10.873 58.513 10.937 ;
			RECT	102.497 10.873 102.529 10.937 ;
			RECT	102.626 10.873 102.69 10.937 ;
			RECT	103.512 10.873 103.576 10.937 ;
			RECT	103.673 10.873 103.705 10.937 ;
			RECT	147.689 10.873 147.721 10.937 ;
			RECT	147.818 10.873 147.882 10.937 ;
			RECT	156.318 10.873 156.382 10.937 ;
			RECT	156.479 10.873 156.511 10.937 ;
			RECT	200.495 10.873 200.527 10.937 ;
			RECT	200.624 10.873 200.688 10.937 ;
			RECT	201.14 10.889 201.204 10.921 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 8.93 201.665 9.04 ;
			LAYER	J3 ;
			RECT	5.514 8.953 5.578 9.017 ;
			RECT	5.675 8.953 5.707 9.017 ;
			RECT	49.691 8.953 49.723 9.017 ;
			RECT	49.82 8.953 49.884 9.017 ;
			RECT	58.32 8.953 58.384 9.017 ;
			RECT	58.481 8.953 58.513 9.017 ;
			RECT	102.497 8.953 102.529 9.017 ;
			RECT	102.626 8.953 102.69 9.017 ;
			RECT	103.512 8.953 103.576 9.017 ;
			RECT	103.673 8.953 103.705 9.017 ;
			RECT	147.689 8.953 147.721 9.017 ;
			RECT	147.818 8.953 147.882 9.017 ;
			RECT	156.318 8.953 156.382 9.017 ;
			RECT	156.479 8.953 156.511 9.017 ;
			RECT	200.495 8.953 200.527 9.017 ;
			RECT	200.624 8.953 200.688 9.017 ;
			RECT	201.14 8.969 201.204 9.001 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 7.01 201.665 7.12 ;
			LAYER	J3 ;
			RECT	5.514 7.033 5.578 7.097 ;
			RECT	5.675 7.033 5.707 7.097 ;
			RECT	49.691 7.033 49.723 7.097 ;
			RECT	49.82 7.033 49.884 7.097 ;
			RECT	58.32 7.033 58.384 7.097 ;
			RECT	58.481 7.033 58.513 7.097 ;
			RECT	102.497 7.033 102.529 7.097 ;
			RECT	102.626 7.033 102.69 7.097 ;
			RECT	103.512 7.033 103.576 7.097 ;
			RECT	103.673 7.033 103.705 7.097 ;
			RECT	147.689 7.033 147.721 7.097 ;
			RECT	147.818 7.033 147.882 7.097 ;
			RECT	156.318 7.033 156.382 7.097 ;
			RECT	156.479 7.033 156.511 7.097 ;
			RECT	200.495 7.033 200.527 7.097 ;
			RECT	200.624 7.033 200.688 7.097 ;
			RECT	201.14 7.049 201.204 7.081 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 5.09 201.665 5.2 ;
			LAYER	J3 ;
			RECT	5.514 5.113 5.578 5.177 ;
			RECT	5.675 5.113 5.707 5.177 ;
			RECT	49.691 5.113 49.723 5.177 ;
			RECT	49.82 5.113 49.884 5.177 ;
			RECT	58.32 5.113 58.384 5.177 ;
			RECT	58.481 5.113 58.513 5.177 ;
			RECT	102.497 5.113 102.529 5.177 ;
			RECT	102.626 5.113 102.69 5.177 ;
			RECT	103.512 5.113 103.576 5.177 ;
			RECT	103.673 5.113 103.705 5.177 ;
			RECT	147.689 5.113 147.721 5.177 ;
			RECT	147.818 5.113 147.882 5.177 ;
			RECT	156.318 5.113 156.382 5.177 ;
			RECT	156.479 5.113 156.511 5.177 ;
			RECT	200.495 5.113 200.527 5.177 ;
			RECT	200.624 5.113 200.688 5.177 ;
			RECT	201.14 5.129 201.204 5.161 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 3.17 201.665 3.28 ;
			LAYER	J3 ;
			RECT	5.514 3.193 5.578 3.257 ;
			RECT	5.675 3.193 5.707 3.257 ;
			RECT	49.691 3.193 49.723 3.257 ;
			RECT	49.82 3.193 49.884 3.257 ;
			RECT	58.32 3.193 58.384 3.257 ;
			RECT	58.481 3.193 58.513 3.257 ;
			RECT	102.497 3.193 102.529 3.257 ;
			RECT	102.626 3.193 102.69 3.257 ;
			RECT	103.512 3.193 103.576 3.257 ;
			RECT	103.673 3.193 103.705 3.257 ;
			RECT	147.689 3.193 147.721 3.257 ;
			RECT	147.818 3.193 147.882 3.257 ;
			RECT	156.318 3.193 156.382 3.257 ;
			RECT	156.479 3.193 156.511 3.257 ;
			RECT	200.495 3.193 200.527 3.257 ;
			RECT	200.624 3.193 200.688 3.257 ;
			RECT	201.14 3.209 201.204 3.241 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 1.25 201.665 1.36 ;
			LAYER	J3 ;
			RECT	5.514 1.273 5.578 1.337 ;
			RECT	5.675 1.273 5.707 1.337 ;
			RECT	49.691 1.273 49.723 1.337 ;
			RECT	49.82 1.273 49.884 1.337 ;
			RECT	58.32 1.273 58.384 1.337 ;
			RECT	58.481 1.273 58.513 1.337 ;
			RECT	102.497 1.273 102.529 1.337 ;
			RECT	102.626 1.273 102.69 1.337 ;
			RECT	103.512 1.273 103.576 1.337 ;
			RECT	103.673 1.273 103.705 1.337 ;
			RECT	147.689 1.273 147.721 1.337 ;
			RECT	147.818 1.273 147.882 1.337 ;
			RECT	156.318 1.273 156.382 1.337 ;
			RECT	156.479 1.273 156.511 1.337 ;
			RECT	200.495 1.273 200.527 1.337 ;
			RECT	200.624 1.273 200.688 1.337 ;
			RECT	201.14 1.289 201.204 1.321 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 73.136 201.665 73.246 ;
			LAYER	J3 ;
			RECT	5.514 73.159 5.578 73.223 ;
			RECT	5.675 73.159 5.707 73.223 ;
			RECT	49.691 73.159 49.723 73.223 ;
			RECT	49.82 73.159 49.884 73.223 ;
			RECT	58.32 73.159 58.384 73.223 ;
			RECT	58.481 73.159 58.513 73.223 ;
			RECT	102.497 73.159 102.529 73.223 ;
			RECT	102.626 73.159 102.69 73.223 ;
			RECT	103.512 73.159 103.576 73.223 ;
			RECT	103.673 73.159 103.705 73.223 ;
			RECT	147.689 73.159 147.721 73.223 ;
			RECT	147.818 73.159 147.882 73.223 ;
			RECT	156.318 73.159 156.382 73.223 ;
			RECT	156.479 73.159 156.511 73.223 ;
			RECT	200.495 73.159 200.527 73.223 ;
			RECT	200.624 73.159 200.688 73.223 ;
			RECT	201.14 73.175 201.204 73.207 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 71.216 201.665 71.326 ;
			LAYER	J3 ;
			RECT	5.514 71.239 5.578 71.303 ;
			RECT	5.675 71.239 5.707 71.303 ;
			RECT	49.691 71.239 49.723 71.303 ;
			RECT	49.82 71.239 49.884 71.303 ;
			RECT	58.32 71.239 58.384 71.303 ;
			RECT	58.481 71.239 58.513 71.303 ;
			RECT	102.497 71.239 102.529 71.303 ;
			RECT	102.626 71.239 102.69 71.303 ;
			RECT	103.512 71.239 103.576 71.303 ;
			RECT	103.673 71.239 103.705 71.303 ;
			RECT	147.689 71.239 147.721 71.303 ;
			RECT	147.818 71.239 147.882 71.303 ;
			RECT	156.318 71.239 156.382 71.303 ;
			RECT	156.479 71.239 156.511 71.303 ;
			RECT	200.495 71.239 200.527 71.303 ;
			RECT	200.624 71.239 200.688 71.303 ;
			RECT	201.14 71.255 201.204 71.287 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 69.296 201.665 69.406 ;
			LAYER	J3 ;
			RECT	5.514 69.319 5.578 69.383 ;
			RECT	5.675 69.319 5.707 69.383 ;
			RECT	49.691 69.319 49.723 69.383 ;
			RECT	49.82 69.319 49.884 69.383 ;
			RECT	58.32 69.319 58.384 69.383 ;
			RECT	58.481 69.319 58.513 69.383 ;
			RECT	102.497 69.319 102.529 69.383 ;
			RECT	102.626 69.319 102.69 69.383 ;
			RECT	103.512 69.319 103.576 69.383 ;
			RECT	103.673 69.319 103.705 69.383 ;
			RECT	147.689 69.319 147.721 69.383 ;
			RECT	147.818 69.319 147.882 69.383 ;
			RECT	156.318 69.319 156.382 69.383 ;
			RECT	156.479 69.319 156.511 69.383 ;
			RECT	200.495 69.319 200.527 69.383 ;
			RECT	200.624 69.319 200.688 69.383 ;
			RECT	201.14 69.335 201.204 69.367 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 67.376 201.665 67.486 ;
			LAYER	J3 ;
			RECT	5.514 67.399 5.578 67.463 ;
			RECT	5.675 67.399 5.707 67.463 ;
			RECT	49.691 67.399 49.723 67.463 ;
			RECT	49.82 67.399 49.884 67.463 ;
			RECT	58.32 67.399 58.384 67.463 ;
			RECT	58.481 67.399 58.513 67.463 ;
			RECT	102.497 67.399 102.529 67.463 ;
			RECT	102.626 67.399 102.69 67.463 ;
			RECT	103.512 67.399 103.576 67.463 ;
			RECT	103.673 67.399 103.705 67.463 ;
			RECT	147.689 67.399 147.721 67.463 ;
			RECT	147.818 67.399 147.882 67.463 ;
			RECT	156.318 67.399 156.382 67.463 ;
			RECT	156.479 67.399 156.511 67.463 ;
			RECT	200.495 67.399 200.527 67.463 ;
			RECT	200.624 67.399 200.688 67.463 ;
			RECT	201.14 67.415 201.204 67.447 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 65.456 201.665 65.566 ;
			LAYER	J3 ;
			RECT	5.514 65.479 5.578 65.543 ;
			RECT	5.675 65.479 5.707 65.543 ;
			RECT	49.691 65.479 49.723 65.543 ;
			RECT	49.82 65.479 49.884 65.543 ;
			RECT	58.32 65.479 58.384 65.543 ;
			RECT	58.481 65.479 58.513 65.543 ;
			RECT	102.497 65.479 102.529 65.543 ;
			RECT	102.626 65.479 102.69 65.543 ;
			RECT	103.512 65.479 103.576 65.543 ;
			RECT	103.673 65.479 103.705 65.543 ;
			RECT	147.689 65.479 147.721 65.543 ;
			RECT	147.818 65.479 147.882 65.543 ;
			RECT	156.318 65.479 156.382 65.543 ;
			RECT	156.479 65.479 156.511 65.543 ;
			RECT	200.495 65.479 200.527 65.543 ;
			RECT	200.624 65.479 200.688 65.543 ;
			RECT	201.14 65.495 201.204 65.527 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 63.536 201.665 63.646 ;
			LAYER	J3 ;
			RECT	5.514 63.559 5.578 63.623 ;
			RECT	5.675 63.559 5.707 63.623 ;
			RECT	49.691 63.559 49.723 63.623 ;
			RECT	49.82 63.559 49.884 63.623 ;
			RECT	58.32 63.559 58.384 63.623 ;
			RECT	58.481 63.559 58.513 63.623 ;
			RECT	102.497 63.559 102.529 63.623 ;
			RECT	102.626 63.559 102.69 63.623 ;
			RECT	103.512 63.559 103.576 63.623 ;
			RECT	103.673 63.559 103.705 63.623 ;
			RECT	147.689 63.559 147.721 63.623 ;
			RECT	147.818 63.559 147.882 63.623 ;
			RECT	156.318 63.559 156.382 63.623 ;
			RECT	156.479 63.559 156.511 63.623 ;
			RECT	200.495 63.559 200.527 63.623 ;
			RECT	200.624 63.559 200.688 63.623 ;
			RECT	201.14 63.575 201.204 63.607 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 61.616 201.665 61.726 ;
			LAYER	J3 ;
			RECT	5.514 61.639 5.578 61.703 ;
			RECT	5.675 61.639 5.707 61.703 ;
			RECT	49.691 61.639 49.723 61.703 ;
			RECT	49.82 61.639 49.884 61.703 ;
			RECT	58.32 61.639 58.384 61.703 ;
			RECT	58.481 61.639 58.513 61.703 ;
			RECT	102.497 61.639 102.529 61.703 ;
			RECT	102.626 61.639 102.69 61.703 ;
			RECT	103.512 61.639 103.576 61.703 ;
			RECT	103.673 61.639 103.705 61.703 ;
			RECT	147.689 61.639 147.721 61.703 ;
			RECT	147.818 61.639 147.882 61.703 ;
			RECT	156.318 61.639 156.382 61.703 ;
			RECT	156.479 61.639 156.511 61.703 ;
			RECT	200.495 61.639 200.527 61.703 ;
			RECT	200.624 61.639 200.688 61.703 ;
			RECT	201.14 61.655 201.204 61.687 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 59.696 201.665 59.806 ;
			LAYER	J3 ;
			RECT	5.514 59.719 5.578 59.783 ;
			RECT	5.675 59.719 5.707 59.783 ;
			RECT	49.691 59.719 49.723 59.783 ;
			RECT	49.82 59.719 49.884 59.783 ;
			RECT	58.32 59.719 58.384 59.783 ;
			RECT	58.481 59.719 58.513 59.783 ;
			RECT	102.497 59.719 102.529 59.783 ;
			RECT	102.626 59.719 102.69 59.783 ;
			RECT	103.512 59.719 103.576 59.783 ;
			RECT	103.673 59.719 103.705 59.783 ;
			RECT	147.689 59.719 147.721 59.783 ;
			RECT	147.818 59.719 147.882 59.783 ;
			RECT	156.318 59.719 156.382 59.783 ;
			RECT	156.479 59.719 156.511 59.783 ;
			RECT	200.495 59.719 200.527 59.783 ;
			RECT	200.624 59.719 200.688 59.783 ;
			RECT	201.14 59.735 201.204 59.767 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 57.776 201.665 57.886 ;
			LAYER	J3 ;
			RECT	5.514 57.799 5.578 57.863 ;
			RECT	5.675 57.799 5.707 57.863 ;
			RECT	49.691 57.799 49.723 57.863 ;
			RECT	49.82 57.799 49.884 57.863 ;
			RECT	58.32 57.799 58.384 57.863 ;
			RECT	58.481 57.799 58.513 57.863 ;
			RECT	102.497 57.799 102.529 57.863 ;
			RECT	102.626 57.799 102.69 57.863 ;
			RECT	103.512 57.799 103.576 57.863 ;
			RECT	103.673 57.799 103.705 57.863 ;
			RECT	147.689 57.799 147.721 57.863 ;
			RECT	147.818 57.799 147.882 57.863 ;
			RECT	156.318 57.799 156.382 57.863 ;
			RECT	156.479 57.799 156.511 57.863 ;
			RECT	200.495 57.799 200.527 57.863 ;
			RECT	200.624 57.799 200.688 57.863 ;
			RECT	201.14 57.815 201.204 57.847 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 55.856 201.665 55.966 ;
			LAYER	J3 ;
			RECT	5.514 55.879 5.578 55.943 ;
			RECT	5.675 55.879 5.707 55.943 ;
			RECT	49.691 55.879 49.723 55.943 ;
			RECT	49.82 55.879 49.884 55.943 ;
			RECT	58.32 55.879 58.384 55.943 ;
			RECT	58.481 55.879 58.513 55.943 ;
			RECT	102.497 55.879 102.529 55.943 ;
			RECT	102.626 55.879 102.69 55.943 ;
			RECT	103.512 55.879 103.576 55.943 ;
			RECT	103.673 55.879 103.705 55.943 ;
			RECT	147.689 55.879 147.721 55.943 ;
			RECT	147.818 55.879 147.882 55.943 ;
			RECT	156.318 55.879 156.382 55.943 ;
			RECT	156.479 55.879 156.511 55.943 ;
			RECT	200.495 55.879 200.527 55.943 ;
			RECT	200.624 55.879 200.688 55.943 ;
			RECT	201.14 55.895 201.204 55.927 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 53.936 201.665 54.046 ;
			LAYER	J3 ;
			RECT	5.514 53.959 5.578 54.023 ;
			RECT	5.675 53.959 5.707 54.023 ;
			RECT	49.691 53.959 49.723 54.023 ;
			RECT	49.82 53.959 49.884 54.023 ;
			RECT	58.32 53.959 58.384 54.023 ;
			RECT	58.481 53.959 58.513 54.023 ;
			RECT	102.497 53.959 102.529 54.023 ;
			RECT	102.626 53.959 102.69 54.023 ;
			RECT	103.512 53.959 103.576 54.023 ;
			RECT	103.673 53.959 103.705 54.023 ;
			RECT	147.689 53.959 147.721 54.023 ;
			RECT	147.818 53.959 147.882 54.023 ;
			RECT	156.318 53.959 156.382 54.023 ;
			RECT	156.479 53.959 156.511 54.023 ;
			RECT	200.495 53.959 200.527 54.023 ;
			RECT	200.624 53.959 200.688 54.023 ;
			RECT	201.14 53.975 201.204 54.007 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 52.016 201.665 52.126 ;
			LAYER	J3 ;
			RECT	5.514 52.039 5.578 52.103 ;
			RECT	5.675 52.039 5.707 52.103 ;
			RECT	49.691 52.039 49.723 52.103 ;
			RECT	49.82 52.039 49.884 52.103 ;
			RECT	58.32 52.039 58.384 52.103 ;
			RECT	58.481 52.039 58.513 52.103 ;
			RECT	102.497 52.039 102.529 52.103 ;
			RECT	102.626 52.039 102.69 52.103 ;
			RECT	103.512 52.039 103.576 52.103 ;
			RECT	103.673 52.039 103.705 52.103 ;
			RECT	147.689 52.039 147.721 52.103 ;
			RECT	147.818 52.039 147.882 52.103 ;
			RECT	156.318 52.039 156.382 52.103 ;
			RECT	156.479 52.039 156.511 52.103 ;
			RECT	200.495 52.039 200.527 52.103 ;
			RECT	200.624 52.039 200.688 52.103 ;
			RECT	201.14 52.055 201.204 52.087 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 78.896 201.665 79.006 ;
			LAYER	J3 ;
			RECT	5.514 78.919 5.578 78.983 ;
			RECT	5.675 78.919 5.707 78.983 ;
			RECT	49.691 78.919 49.723 78.983 ;
			RECT	49.82 78.919 49.884 78.983 ;
			RECT	58.32 78.919 58.384 78.983 ;
			RECT	58.481 78.919 58.513 78.983 ;
			RECT	102.497 78.919 102.529 78.983 ;
			RECT	102.626 78.919 102.69 78.983 ;
			RECT	103.512 78.919 103.576 78.983 ;
			RECT	103.673 78.919 103.705 78.983 ;
			RECT	147.689 78.919 147.721 78.983 ;
			RECT	147.818 78.919 147.882 78.983 ;
			RECT	156.318 78.919 156.382 78.983 ;
			RECT	156.479 78.919 156.511 78.983 ;
			RECT	200.495 78.919 200.527 78.983 ;
			RECT	200.624 78.919 200.688 78.983 ;
			RECT	201.14 78.935 201.204 78.967 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 35.362 201.665 35.482 ;
			LAYER	J3 ;
			RECT	4.982 35.39 5.014 35.454 ;
			RECT	5.514 35.39 5.578 35.454 ;
			RECT	5.848 35.39 5.88 35.454 ;
			RECT	6.379 35.39 6.411 35.454 ;
			RECT	6.715 35.39 6.747 35.454 ;
			RECT	7.051 35.39 7.083 35.454 ;
			RECT	7.387 35.39 7.419 35.454 ;
			RECT	7.723 35.39 7.755 35.454 ;
			RECT	8.059 35.39 8.091 35.454 ;
			RECT	8.395 35.39 8.427 35.454 ;
			RECT	8.731 35.39 8.763 35.454 ;
			RECT	9.067 35.39 9.099 35.454 ;
			RECT	9.403 35.39 9.435 35.454 ;
			RECT	9.739 35.39 9.771 35.454 ;
			RECT	10.075 35.39 10.107 35.454 ;
			RECT	10.411 35.39 10.443 35.454 ;
			RECT	10.747 35.39 10.779 35.454 ;
			RECT	11.083 35.39 11.115 35.454 ;
			RECT	11.419 35.39 11.451 35.454 ;
			RECT	11.755 35.39 11.787 35.454 ;
			RECT	12.091 35.39 12.123 35.454 ;
			RECT	12.427 35.39 12.459 35.454 ;
			RECT	12.763 35.39 12.795 35.454 ;
			RECT	13.099 35.39 13.131 35.454 ;
			RECT	13.435 35.39 13.467 35.454 ;
			RECT	13.771 35.39 13.803 35.454 ;
			RECT	14.107 35.39 14.139 35.454 ;
			RECT	14.443 35.39 14.475 35.454 ;
			RECT	14.779 35.39 14.811 35.454 ;
			RECT	15.115 35.39 15.147 35.454 ;
			RECT	15.451 35.39 15.483 35.454 ;
			RECT	15.787 35.39 15.819 35.454 ;
			RECT	16.123 35.39 16.155 35.454 ;
			RECT	16.459 35.39 16.491 35.454 ;
			RECT	16.795 35.39 16.827 35.454 ;
			RECT	17.131 35.39 17.163 35.454 ;
			RECT	17.467 35.39 17.499 35.454 ;
			RECT	17.803 35.39 17.835 35.454 ;
			RECT	18.139 35.39 18.171 35.454 ;
			RECT	18.475 35.39 18.507 35.454 ;
			RECT	18.811 35.39 18.843 35.454 ;
			RECT	19.147 35.39 19.179 35.454 ;
			RECT	19.483 35.39 19.515 35.454 ;
			RECT	19.819 35.39 19.851 35.454 ;
			RECT	20.155 35.39 20.187 35.454 ;
			RECT	20.491 35.39 20.523 35.454 ;
			RECT	20.827 35.39 20.859 35.454 ;
			RECT	21.163 35.39 21.195 35.454 ;
			RECT	21.499 35.39 21.531 35.454 ;
			RECT	21.835 35.39 21.867 35.454 ;
			RECT	22.171 35.39 22.203 35.454 ;
			RECT	22.507 35.39 22.539 35.454 ;
			RECT	22.843 35.39 22.875 35.454 ;
			RECT	23.179 35.39 23.211 35.454 ;
			RECT	23.515 35.39 23.547 35.454 ;
			RECT	23.851 35.39 23.883 35.454 ;
			RECT	24.187 35.39 24.219 35.454 ;
			RECT	24.523 35.39 24.555 35.454 ;
			RECT	24.859 35.39 24.891 35.454 ;
			RECT	25.195 35.39 25.227 35.454 ;
			RECT	25.531 35.39 25.563 35.454 ;
			RECT	25.867 35.39 25.899 35.454 ;
			RECT	26.203 35.39 26.235 35.454 ;
			RECT	26.539 35.39 26.571 35.454 ;
			RECT	26.875 35.39 26.907 35.454 ;
			RECT	27.211 35.39 27.243 35.454 ;
			RECT	27.547 35.39 27.579 35.454 ;
			RECT	27.878 35.39 27.91 35.454 ;
			RECT	28.214 35.39 28.246 35.454 ;
			RECT	28.55 35.39 28.582 35.454 ;
			RECT	28.886 35.39 28.918 35.454 ;
			RECT	29.222 35.39 29.254 35.454 ;
			RECT	29.558 35.39 29.59 35.454 ;
			RECT	29.894 35.39 29.926 35.454 ;
			RECT	30.23 35.39 30.262 35.454 ;
			RECT	30.566 35.39 30.598 35.454 ;
			RECT	30.902 35.39 30.934 35.454 ;
			RECT	31.238 35.39 31.27 35.454 ;
			RECT	31.574 35.39 31.606 35.454 ;
			RECT	31.91 35.39 31.942 35.454 ;
			RECT	32.246 35.39 32.278 35.454 ;
			RECT	32.582 35.39 32.614 35.454 ;
			RECT	32.918 35.39 32.95 35.454 ;
			RECT	33.254 35.39 33.286 35.454 ;
			RECT	33.59 35.39 33.622 35.454 ;
			RECT	33.926 35.39 33.958 35.454 ;
			RECT	34.262 35.39 34.294 35.454 ;
			RECT	34.598 35.39 34.63 35.454 ;
			RECT	34.934 35.39 34.966 35.454 ;
			RECT	35.27 35.39 35.302 35.454 ;
			RECT	35.606 35.39 35.638 35.454 ;
			RECT	35.942 35.39 35.974 35.454 ;
			RECT	36.278 35.39 36.31 35.454 ;
			RECT	36.614 35.39 36.646 35.454 ;
			RECT	36.95 35.39 36.982 35.454 ;
			RECT	37.286 35.39 37.318 35.454 ;
			RECT	37.622 35.39 37.654 35.454 ;
			RECT	37.958 35.39 37.99 35.454 ;
			RECT	38.294 35.39 38.326 35.454 ;
			RECT	38.63 35.39 38.662 35.454 ;
			RECT	38.966 35.39 38.998 35.454 ;
			RECT	39.302 35.39 39.334 35.454 ;
			RECT	39.638 35.39 39.67 35.454 ;
			RECT	39.974 35.39 40.006 35.454 ;
			RECT	40.31 35.39 40.342 35.454 ;
			RECT	40.646 35.39 40.678 35.454 ;
			RECT	40.982 35.39 41.014 35.454 ;
			RECT	41.318 35.39 41.35 35.454 ;
			RECT	41.654 35.39 41.686 35.454 ;
			RECT	41.99 35.39 42.022 35.454 ;
			RECT	42.326 35.39 42.358 35.454 ;
			RECT	42.662 35.39 42.694 35.454 ;
			RECT	42.998 35.39 43.03 35.454 ;
			RECT	43.334 35.39 43.366 35.454 ;
			RECT	43.67 35.39 43.702 35.454 ;
			RECT	44.342 35.39 44.374 35.454 ;
			RECT	44.678 35.39 44.71 35.454 ;
			RECT	45.014 35.39 45.046 35.454 ;
			RECT	45.35 35.39 45.382 35.454 ;
			RECT	45.686 35.39 45.718 35.454 ;
			RECT	46.022 35.39 46.054 35.454 ;
			RECT	46.358 35.39 46.39 35.454 ;
			RECT	46.694 35.39 46.726 35.454 ;
			RECT	47.03 35.39 47.062 35.454 ;
			RECT	47.366 35.39 47.398 35.454 ;
			RECT	47.702 35.39 47.734 35.454 ;
			RECT	48.038 35.39 48.07 35.454 ;
			RECT	48.374 35.39 48.406 35.454 ;
			RECT	48.71 35.39 48.742 35.454 ;
			RECT	49.046 35.39 49.078 35.454 ;
			RECT	49.227 35.39 49.259 35.454 ;
			RECT	49.994 35.39 50.026 35.454 ;
			RECT	50.266 35.39 50.298 35.454 ;
			RECT	52.15 35.39 52.182 35.454 ;
			RECT	58.178 35.39 58.21 35.454 ;
			RECT	58.945 35.39 58.977 35.454 ;
			RECT	59.126 35.39 59.158 35.454 ;
			RECT	59.462 35.39 59.494 35.454 ;
			RECT	59.798 35.39 59.83 35.454 ;
			RECT	60.134 35.39 60.166 35.454 ;
			RECT	60.47 35.39 60.502 35.454 ;
			RECT	60.806 35.39 60.838 35.454 ;
			RECT	61.142 35.39 61.174 35.454 ;
			RECT	61.478 35.39 61.51 35.454 ;
			RECT	61.814 35.39 61.846 35.454 ;
			RECT	62.15 35.39 62.182 35.454 ;
			RECT	62.486 35.39 62.518 35.454 ;
			RECT	62.822 35.39 62.854 35.454 ;
			RECT	63.158 35.39 63.19 35.454 ;
			RECT	63.494 35.39 63.526 35.454 ;
			RECT	63.83 35.39 63.862 35.454 ;
			RECT	64.502 35.39 64.534 35.454 ;
			RECT	64.838 35.39 64.87 35.454 ;
			RECT	65.174 35.39 65.206 35.454 ;
			RECT	65.51 35.39 65.542 35.454 ;
			RECT	65.846 35.39 65.878 35.454 ;
			RECT	66.182 35.39 66.214 35.454 ;
			RECT	66.518 35.39 66.55 35.454 ;
			RECT	66.854 35.39 66.886 35.454 ;
			RECT	67.19 35.39 67.222 35.454 ;
			RECT	67.526 35.39 67.558 35.454 ;
			RECT	67.862 35.39 67.894 35.454 ;
			RECT	68.198 35.39 68.23 35.454 ;
			RECT	68.534 35.39 68.566 35.454 ;
			RECT	68.87 35.39 68.902 35.454 ;
			RECT	69.206 35.39 69.238 35.454 ;
			RECT	69.542 35.39 69.574 35.454 ;
			RECT	69.878 35.39 69.91 35.454 ;
			RECT	70.214 35.39 70.246 35.454 ;
			RECT	70.55 35.39 70.582 35.454 ;
			RECT	70.886 35.39 70.918 35.454 ;
			RECT	71.222 35.39 71.254 35.454 ;
			RECT	71.558 35.39 71.59 35.454 ;
			RECT	71.894 35.39 71.926 35.454 ;
			RECT	72.23 35.39 72.262 35.454 ;
			RECT	72.566 35.39 72.598 35.454 ;
			RECT	72.902 35.39 72.934 35.454 ;
			RECT	73.238 35.39 73.27 35.454 ;
			RECT	73.574 35.39 73.606 35.454 ;
			RECT	73.91 35.39 73.942 35.454 ;
			RECT	74.246 35.39 74.278 35.454 ;
			RECT	74.582 35.39 74.614 35.454 ;
			RECT	74.918 35.39 74.95 35.454 ;
			RECT	75.254 35.39 75.286 35.454 ;
			RECT	75.59 35.39 75.622 35.454 ;
			RECT	75.926 35.39 75.958 35.454 ;
			RECT	76.262 35.39 76.294 35.454 ;
			RECT	76.598 35.39 76.63 35.454 ;
			RECT	76.934 35.39 76.966 35.454 ;
			RECT	77.27 35.39 77.302 35.454 ;
			RECT	77.606 35.39 77.638 35.454 ;
			RECT	77.942 35.39 77.974 35.454 ;
			RECT	78.278 35.39 78.31 35.454 ;
			RECT	78.614 35.39 78.646 35.454 ;
			RECT	78.95 35.39 78.982 35.454 ;
			RECT	79.286 35.39 79.318 35.454 ;
			RECT	79.622 35.39 79.654 35.454 ;
			RECT	79.958 35.39 79.99 35.454 ;
			RECT	80.294 35.39 80.326 35.454 ;
			RECT	80.625 35.39 80.657 35.454 ;
			RECT	80.961 35.39 80.993 35.454 ;
			RECT	81.297 35.39 81.329 35.454 ;
			RECT	81.633 35.39 81.665 35.454 ;
			RECT	81.969 35.39 82.001 35.454 ;
			RECT	82.305 35.39 82.337 35.454 ;
			RECT	82.641 35.39 82.673 35.454 ;
			RECT	82.977 35.39 83.009 35.454 ;
			RECT	83.313 35.39 83.345 35.454 ;
			RECT	83.649 35.39 83.681 35.454 ;
			RECT	83.985 35.39 84.017 35.454 ;
			RECT	84.321 35.39 84.353 35.454 ;
			RECT	84.657 35.39 84.689 35.454 ;
			RECT	84.993 35.39 85.025 35.454 ;
			RECT	85.329 35.39 85.361 35.454 ;
			RECT	85.665 35.39 85.697 35.454 ;
			RECT	86.001 35.39 86.033 35.454 ;
			RECT	86.337 35.39 86.369 35.454 ;
			RECT	86.673 35.39 86.705 35.454 ;
			RECT	87.009 35.39 87.041 35.454 ;
			RECT	87.345 35.39 87.377 35.454 ;
			RECT	87.681 35.39 87.713 35.454 ;
			RECT	88.017 35.39 88.049 35.454 ;
			RECT	88.353 35.39 88.385 35.454 ;
			RECT	88.689 35.39 88.721 35.454 ;
			RECT	89.025 35.39 89.057 35.454 ;
			RECT	89.361 35.39 89.393 35.454 ;
			RECT	89.697 35.39 89.729 35.454 ;
			RECT	90.033 35.39 90.065 35.454 ;
			RECT	90.369 35.39 90.401 35.454 ;
			RECT	90.705 35.39 90.737 35.454 ;
			RECT	91.041 35.39 91.073 35.454 ;
			RECT	91.377 35.39 91.409 35.454 ;
			RECT	91.713 35.39 91.745 35.454 ;
			RECT	92.049 35.39 92.081 35.454 ;
			RECT	92.385 35.39 92.417 35.454 ;
			RECT	92.721 35.39 92.753 35.454 ;
			RECT	93.057 35.39 93.089 35.454 ;
			RECT	93.393 35.39 93.425 35.454 ;
			RECT	93.729 35.39 93.761 35.454 ;
			RECT	94.065 35.39 94.097 35.454 ;
			RECT	94.401 35.39 94.433 35.454 ;
			RECT	94.737 35.39 94.769 35.454 ;
			RECT	95.073 35.39 95.105 35.454 ;
			RECT	95.409 35.39 95.441 35.454 ;
			RECT	95.745 35.39 95.777 35.454 ;
			RECT	96.081 35.39 96.113 35.454 ;
			RECT	96.417 35.39 96.449 35.454 ;
			RECT	96.753 35.39 96.785 35.454 ;
			RECT	97.089 35.39 97.121 35.454 ;
			RECT	97.425 35.39 97.457 35.454 ;
			RECT	97.761 35.39 97.793 35.454 ;
			RECT	98.097 35.39 98.129 35.454 ;
			RECT	98.433 35.39 98.465 35.454 ;
			RECT	98.769 35.39 98.801 35.454 ;
			RECT	99.105 35.39 99.137 35.454 ;
			RECT	99.441 35.39 99.473 35.454 ;
			RECT	99.777 35.39 99.809 35.454 ;
			RECT	100.113 35.39 100.145 35.454 ;
			RECT	100.449 35.39 100.481 35.454 ;
			RECT	100.785 35.39 100.817 35.454 ;
			RECT	101.121 35.39 101.153 35.454 ;
			RECT	101.457 35.39 101.489 35.454 ;
			RECT	101.793 35.39 101.825 35.454 ;
			RECT	102.324 35.39 102.356 35.454 ;
			RECT	102.626 35.39 102.69 35.454 ;
			RECT	103.512 35.39 103.576 35.454 ;
			RECT	103.846 35.39 103.878 35.454 ;
			RECT	104.377 35.39 104.409 35.454 ;
			RECT	104.713 35.39 104.745 35.454 ;
			RECT	105.049 35.39 105.081 35.454 ;
			RECT	105.385 35.39 105.417 35.454 ;
			RECT	105.721 35.39 105.753 35.454 ;
			RECT	106.057 35.39 106.089 35.454 ;
			RECT	106.393 35.39 106.425 35.454 ;
			RECT	106.729 35.39 106.761 35.454 ;
			RECT	107.065 35.39 107.097 35.454 ;
			RECT	107.401 35.39 107.433 35.454 ;
			RECT	107.737 35.39 107.769 35.454 ;
			RECT	108.073 35.39 108.105 35.454 ;
			RECT	108.409 35.39 108.441 35.454 ;
			RECT	108.745 35.39 108.777 35.454 ;
			RECT	109.081 35.39 109.113 35.454 ;
			RECT	109.417 35.39 109.449 35.454 ;
			RECT	109.753 35.39 109.785 35.454 ;
			RECT	110.089 35.39 110.121 35.454 ;
			RECT	110.425 35.39 110.457 35.454 ;
			RECT	110.761 35.39 110.793 35.454 ;
			RECT	111.097 35.39 111.129 35.454 ;
			RECT	111.433 35.39 111.465 35.454 ;
			RECT	111.769 35.39 111.801 35.454 ;
			RECT	112.105 35.39 112.137 35.454 ;
			RECT	112.441 35.39 112.473 35.454 ;
			RECT	112.777 35.39 112.809 35.454 ;
			RECT	113.113 35.39 113.145 35.454 ;
			RECT	113.449 35.39 113.481 35.454 ;
			RECT	113.785 35.39 113.817 35.454 ;
			RECT	114.121 35.39 114.153 35.454 ;
			RECT	114.457 35.39 114.489 35.454 ;
			RECT	114.793 35.39 114.825 35.454 ;
			RECT	115.129 35.39 115.161 35.454 ;
			RECT	115.465 35.39 115.497 35.454 ;
			RECT	115.801 35.39 115.833 35.454 ;
			RECT	116.137 35.39 116.169 35.454 ;
			RECT	116.473 35.39 116.505 35.454 ;
			RECT	116.809 35.39 116.841 35.454 ;
			RECT	117.145 35.39 117.177 35.454 ;
			RECT	117.481 35.39 117.513 35.454 ;
			RECT	117.817 35.39 117.849 35.454 ;
			RECT	118.153 35.39 118.185 35.454 ;
			RECT	118.489 35.39 118.521 35.454 ;
			RECT	118.825 35.39 118.857 35.454 ;
			RECT	119.161 35.39 119.193 35.454 ;
			RECT	119.497 35.39 119.529 35.454 ;
			RECT	119.833 35.39 119.865 35.454 ;
			RECT	120.169 35.39 120.201 35.454 ;
			RECT	120.505 35.39 120.537 35.454 ;
			RECT	120.841 35.39 120.873 35.454 ;
			RECT	121.177 35.39 121.209 35.454 ;
			RECT	121.513 35.39 121.545 35.454 ;
			RECT	121.849 35.39 121.881 35.454 ;
			RECT	122.185 35.39 122.217 35.454 ;
			RECT	122.521 35.39 122.553 35.454 ;
			RECT	122.857 35.39 122.889 35.454 ;
			RECT	123.193 35.39 123.225 35.454 ;
			RECT	123.529 35.39 123.561 35.454 ;
			RECT	123.865 35.39 123.897 35.454 ;
			RECT	124.201 35.39 124.233 35.454 ;
			RECT	124.537 35.39 124.569 35.454 ;
			RECT	124.873 35.39 124.905 35.454 ;
			RECT	125.209 35.39 125.241 35.454 ;
			RECT	125.545 35.39 125.577 35.454 ;
			RECT	125.876 35.39 125.908 35.454 ;
			RECT	126.212 35.39 126.244 35.454 ;
			RECT	126.548 35.39 126.58 35.454 ;
			RECT	126.884 35.39 126.916 35.454 ;
			RECT	127.22 35.39 127.252 35.454 ;
			RECT	127.556 35.39 127.588 35.454 ;
			RECT	127.892 35.39 127.924 35.454 ;
			RECT	128.228 35.39 128.26 35.454 ;
			RECT	128.564 35.39 128.596 35.454 ;
			RECT	128.9 35.39 128.932 35.454 ;
			RECT	129.236 35.39 129.268 35.454 ;
			RECT	129.572 35.39 129.604 35.454 ;
			RECT	129.908 35.39 129.94 35.454 ;
			RECT	130.244 35.39 130.276 35.454 ;
			RECT	130.58 35.39 130.612 35.454 ;
			RECT	130.916 35.39 130.948 35.454 ;
			RECT	131.252 35.39 131.284 35.454 ;
			RECT	131.588 35.39 131.62 35.454 ;
			RECT	131.924 35.39 131.956 35.454 ;
			RECT	132.26 35.39 132.292 35.454 ;
			RECT	132.596 35.39 132.628 35.454 ;
			RECT	132.932 35.39 132.964 35.454 ;
			RECT	133.268 35.39 133.3 35.454 ;
			RECT	133.604 35.39 133.636 35.454 ;
			RECT	133.94 35.39 133.972 35.454 ;
			RECT	134.276 35.39 134.308 35.454 ;
			RECT	134.612 35.39 134.644 35.454 ;
			RECT	134.948 35.39 134.98 35.454 ;
			RECT	135.284 35.39 135.316 35.454 ;
			RECT	135.62 35.39 135.652 35.454 ;
			RECT	135.956 35.39 135.988 35.454 ;
			RECT	136.292 35.39 136.324 35.454 ;
			RECT	136.628 35.39 136.66 35.454 ;
			RECT	136.964 35.39 136.996 35.454 ;
			RECT	137.3 35.39 137.332 35.454 ;
			RECT	137.636 35.39 137.668 35.454 ;
			RECT	137.972 35.39 138.004 35.454 ;
			RECT	138.308 35.39 138.34 35.454 ;
			RECT	138.644 35.39 138.676 35.454 ;
			RECT	138.98 35.39 139.012 35.454 ;
			RECT	139.316 35.39 139.348 35.454 ;
			RECT	139.652 35.39 139.684 35.454 ;
			RECT	139.988 35.39 140.02 35.454 ;
			RECT	140.324 35.39 140.356 35.454 ;
			RECT	140.66 35.39 140.692 35.454 ;
			RECT	140.996 35.39 141.028 35.454 ;
			RECT	141.332 35.39 141.364 35.454 ;
			RECT	141.668 35.39 141.7 35.454 ;
			RECT	142.34 35.39 142.372 35.454 ;
			RECT	142.676 35.39 142.708 35.454 ;
			RECT	143.012 35.39 143.044 35.454 ;
			RECT	143.348 35.39 143.38 35.454 ;
			RECT	143.684 35.39 143.716 35.454 ;
			RECT	144.02 35.39 144.052 35.454 ;
			RECT	144.356 35.39 144.388 35.454 ;
			RECT	144.692 35.39 144.724 35.454 ;
			RECT	145.028 35.39 145.06 35.454 ;
			RECT	145.364 35.39 145.396 35.454 ;
			RECT	145.7 35.39 145.732 35.454 ;
			RECT	146.036 35.39 146.068 35.454 ;
			RECT	146.372 35.39 146.404 35.454 ;
			RECT	146.708 35.39 146.74 35.454 ;
			RECT	147.044 35.39 147.076 35.454 ;
			RECT	147.225 35.39 147.257 35.454 ;
			RECT	147.992 35.39 148.024 35.454 ;
			RECT	148.264 35.39 148.296 35.454 ;
			RECT	150.148 35.39 150.18 35.454 ;
			RECT	156.176 35.39 156.208 35.454 ;
			RECT	156.943 35.39 156.975 35.454 ;
			RECT	157.124 35.39 157.156 35.454 ;
			RECT	157.46 35.39 157.492 35.454 ;
			RECT	157.796 35.39 157.828 35.454 ;
			RECT	158.132 35.39 158.164 35.454 ;
			RECT	158.468 35.39 158.5 35.454 ;
			RECT	158.804 35.39 158.836 35.454 ;
			RECT	159.14 35.39 159.172 35.454 ;
			RECT	159.476 35.39 159.508 35.454 ;
			RECT	159.812 35.39 159.844 35.454 ;
			RECT	160.148 35.39 160.18 35.454 ;
			RECT	160.484 35.39 160.516 35.454 ;
			RECT	160.82 35.39 160.852 35.454 ;
			RECT	161.156 35.39 161.188 35.454 ;
			RECT	161.492 35.39 161.524 35.454 ;
			RECT	161.828 35.39 161.86 35.454 ;
			RECT	162.5 35.39 162.532 35.454 ;
			RECT	162.836 35.39 162.868 35.454 ;
			RECT	163.172 35.39 163.204 35.454 ;
			RECT	163.508 35.39 163.54 35.454 ;
			RECT	163.844 35.39 163.876 35.454 ;
			RECT	164.18 35.39 164.212 35.454 ;
			RECT	164.516 35.39 164.548 35.454 ;
			RECT	164.852 35.39 164.884 35.454 ;
			RECT	165.188 35.39 165.22 35.454 ;
			RECT	165.524 35.39 165.556 35.454 ;
			RECT	165.86 35.39 165.892 35.454 ;
			RECT	166.196 35.39 166.228 35.454 ;
			RECT	166.532 35.39 166.564 35.454 ;
			RECT	166.868 35.39 166.9 35.454 ;
			RECT	167.204 35.39 167.236 35.454 ;
			RECT	167.54 35.39 167.572 35.454 ;
			RECT	167.876 35.39 167.908 35.454 ;
			RECT	168.212 35.39 168.244 35.454 ;
			RECT	168.548 35.39 168.58 35.454 ;
			RECT	168.884 35.39 168.916 35.454 ;
			RECT	169.22 35.39 169.252 35.454 ;
			RECT	169.556 35.39 169.588 35.454 ;
			RECT	169.892 35.39 169.924 35.454 ;
			RECT	170.228 35.39 170.26 35.454 ;
			RECT	170.564 35.39 170.596 35.454 ;
			RECT	170.9 35.39 170.932 35.454 ;
			RECT	171.236 35.39 171.268 35.454 ;
			RECT	171.572 35.39 171.604 35.454 ;
			RECT	171.908 35.39 171.94 35.454 ;
			RECT	172.244 35.39 172.276 35.454 ;
			RECT	172.58 35.39 172.612 35.454 ;
			RECT	172.916 35.39 172.948 35.454 ;
			RECT	173.252 35.39 173.284 35.454 ;
			RECT	173.588 35.39 173.62 35.454 ;
			RECT	173.924 35.39 173.956 35.454 ;
			RECT	174.26 35.39 174.292 35.454 ;
			RECT	174.596 35.39 174.628 35.454 ;
			RECT	174.932 35.39 174.964 35.454 ;
			RECT	175.268 35.39 175.3 35.454 ;
			RECT	175.604 35.39 175.636 35.454 ;
			RECT	175.94 35.39 175.972 35.454 ;
			RECT	176.276 35.39 176.308 35.454 ;
			RECT	176.612 35.39 176.644 35.454 ;
			RECT	176.948 35.39 176.98 35.454 ;
			RECT	177.284 35.39 177.316 35.454 ;
			RECT	177.62 35.39 177.652 35.454 ;
			RECT	177.956 35.39 177.988 35.454 ;
			RECT	178.292 35.39 178.324 35.454 ;
			RECT	178.623 35.39 178.655 35.454 ;
			RECT	178.959 35.39 178.991 35.454 ;
			RECT	179.295 35.39 179.327 35.454 ;
			RECT	179.631 35.39 179.663 35.454 ;
			RECT	179.967 35.39 179.999 35.454 ;
			RECT	180.303 35.39 180.335 35.454 ;
			RECT	180.639 35.39 180.671 35.454 ;
			RECT	180.975 35.39 181.007 35.454 ;
			RECT	181.311 35.39 181.343 35.454 ;
			RECT	181.647 35.39 181.679 35.454 ;
			RECT	181.983 35.39 182.015 35.454 ;
			RECT	182.319 35.39 182.351 35.454 ;
			RECT	182.655 35.39 182.687 35.454 ;
			RECT	182.991 35.39 183.023 35.454 ;
			RECT	183.327 35.39 183.359 35.454 ;
			RECT	183.663 35.39 183.695 35.454 ;
			RECT	183.999 35.39 184.031 35.454 ;
			RECT	184.335 35.39 184.367 35.454 ;
			RECT	184.671 35.39 184.703 35.454 ;
			RECT	185.007 35.39 185.039 35.454 ;
			RECT	185.343 35.39 185.375 35.454 ;
			RECT	185.679 35.39 185.711 35.454 ;
			RECT	186.015 35.39 186.047 35.454 ;
			RECT	186.351 35.39 186.383 35.454 ;
			RECT	186.687 35.39 186.719 35.454 ;
			RECT	187.023 35.39 187.055 35.454 ;
			RECT	187.359 35.39 187.391 35.454 ;
			RECT	187.695 35.39 187.727 35.454 ;
			RECT	188.031 35.39 188.063 35.454 ;
			RECT	188.367 35.39 188.399 35.454 ;
			RECT	188.703 35.39 188.735 35.454 ;
			RECT	189.039 35.39 189.071 35.454 ;
			RECT	189.375 35.39 189.407 35.454 ;
			RECT	189.711 35.39 189.743 35.454 ;
			RECT	190.047 35.39 190.079 35.454 ;
			RECT	190.383 35.39 190.415 35.454 ;
			RECT	190.719 35.39 190.751 35.454 ;
			RECT	191.055 35.39 191.087 35.454 ;
			RECT	191.391 35.39 191.423 35.454 ;
			RECT	191.727 35.39 191.759 35.454 ;
			RECT	192.063 35.39 192.095 35.454 ;
			RECT	192.399 35.39 192.431 35.454 ;
			RECT	192.735 35.39 192.767 35.454 ;
			RECT	193.071 35.39 193.103 35.454 ;
			RECT	193.407 35.39 193.439 35.454 ;
			RECT	193.743 35.39 193.775 35.454 ;
			RECT	194.079 35.39 194.111 35.454 ;
			RECT	194.415 35.39 194.447 35.454 ;
			RECT	194.751 35.39 194.783 35.454 ;
			RECT	195.087 35.39 195.119 35.454 ;
			RECT	195.423 35.39 195.455 35.454 ;
			RECT	195.759 35.39 195.791 35.454 ;
			RECT	196.095 35.39 196.127 35.454 ;
			RECT	196.431 35.39 196.463 35.454 ;
			RECT	196.767 35.39 196.799 35.454 ;
			RECT	197.103 35.39 197.135 35.454 ;
			RECT	197.439 35.39 197.471 35.454 ;
			RECT	197.775 35.39 197.807 35.454 ;
			RECT	198.111 35.39 198.143 35.454 ;
			RECT	198.447 35.39 198.479 35.454 ;
			RECT	198.783 35.39 198.815 35.454 ;
			RECT	199.119 35.39 199.151 35.454 ;
			RECT	199.455 35.39 199.487 35.454 ;
			RECT	199.791 35.39 199.823 35.454 ;
			RECT	200.322 35.39 200.354 35.454 ;
			RECT	200.624 35.39 200.688 35.454 ;
			RECT	201.14 35.39 201.204 35.454 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 36.845 201.665 36.965 ;
			LAYER	J3 ;
			RECT	5.848 36.873 5.88 36.937 ;
			RECT	6.379 36.873 6.411 36.937 ;
			RECT	6.715 36.873 6.747 36.937 ;
			RECT	7.051 36.873 7.083 36.937 ;
			RECT	7.387 36.873 7.419 36.937 ;
			RECT	7.723 36.873 7.755 36.937 ;
			RECT	8.059 36.873 8.091 36.937 ;
			RECT	8.395 36.873 8.427 36.937 ;
			RECT	8.731 36.873 8.763 36.937 ;
			RECT	9.067 36.873 9.099 36.937 ;
			RECT	9.403 36.873 9.435 36.937 ;
			RECT	9.739 36.873 9.771 36.937 ;
			RECT	10.075 36.873 10.107 36.937 ;
			RECT	10.411 36.873 10.443 36.937 ;
			RECT	10.747 36.873 10.779 36.937 ;
			RECT	11.083 36.873 11.115 36.937 ;
			RECT	11.419 36.873 11.451 36.937 ;
			RECT	11.755 36.873 11.787 36.937 ;
			RECT	12.091 36.873 12.123 36.937 ;
			RECT	12.427 36.873 12.459 36.937 ;
			RECT	12.763 36.873 12.795 36.937 ;
			RECT	13.099 36.873 13.131 36.937 ;
			RECT	13.435 36.873 13.467 36.937 ;
			RECT	13.771 36.873 13.803 36.937 ;
			RECT	14.107 36.873 14.139 36.937 ;
			RECT	14.443 36.873 14.475 36.937 ;
			RECT	14.779 36.873 14.811 36.937 ;
			RECT	15.115 36.873 15.147 36.937 ;
			RECT	15.451 36.873 15.483 36.937 ;
			RECT	15.787 36.873 15.819 36.937 ;
			RECT	16.123 36.873 16.155 36.937 ;
			RECT	16.459 36.873 16.491 36.937 ;
			RECT	16.795 36.873 16.827 36.937 ;
			RECT	17.131 36.873 17.163 36.937 ;
			RECT	17.467 36.873 17.499 36.937 ;
			RECT	17.803 36.873 17.835 36.937 ;
			RECT	18.139 36.873 18.171 36.937 ;
			RECT	18.475 36.873 18.507 36.937 ;
			RECT	18.811 36.873 18.843 36.937 ;
			RECT	19.147 36.873 19.179 36.937 ;
			RECT	19.483 36.873 19.515 36.937 ;
			RECT	19.819 36.873 19.851 36.937 ;
			RECT	20.155 36.873 20.187 36.937 ;
			RECT	20.491 36.873 20.523 36.937 ;
			RECT	20.827 36.873 20.859 36.937 ;
			RECT	21.163 36.873 21.195 36.937 ;
			RECT	21.499 36.873 21.531 36.937 ;
			RECT	21.835 36.873 21.867 36.937 ;
			RECT	22.171 36.873 22.203 36.937 ;
			RECT	22.507 36.873 22.539 36.937 ;
			RECT	22.843 36.873 22.875 36.937 ;
			RECT	23.179 36.873 23.211 36.937 ;
			RECT	23.515 36.873 23.547 36.937 ;
			RECT	23.851 36.873 23.883 36.937 ;
			RECT	24.187 36.873 24.219 36.937 ;
			RECT	24.523 36.873 24.555 36.937 ;
			RECT	24.859 36.873 24.891 36.937 ;
			RECT	25.195 36.873 25.227 36.937 ;
			RECT	25.531 36.873 25.563 36.937 ;
			RECT	25.867 36.873 25.899 36.937 ;
			RECT	26.203 36.873 26.235 36.937 ;
			RECT	26.539 36.873 26.571 36.937 ;
			RECT	26.875 36.873 26.907 36.937 ;
			RECT	27.211 36.873 27.243 36.937 ;
			RECT	27.547 36.873 27.579 36.937 ;
			RECT	27.878 36.873 27.91 36.937 ;
			RECT	28.214 36.873 28.246 36.937 ;
			RECT	28.55 36.873 28.582 36.937 ;
			RECT	28.886 36.873 28.918 36.937 ;
			RECT	29.222 36.873 29.254 36.937 ;
			RECT	29.558 36.873 29.59 36.937 ;
			RECT	29.894 36.873 29.926 36.937 ;
			RECT	30.23 36.873 30.262 36.937 ;
			RECT	30.566 36.873 30.598 36.937 ;
			RECT	30.902 36.873 30.934 36.937 ;
			RECT	31.238 36.873 31.27 36.937 ;
			RECT	31.574 36.873 31.606 36.937 ;
			RECT	31.91 36.873 31.942 36.937 ;
			RECT	32.246 36.873 32.278 36.937 ;
			RECT	32.582 36.873 32.614 36.937 ;
			RECT	32.918 36.873 32.95 36.937 ;
			RECT	33.254 36.873 33.286 36.937 ;
			RECT	33.59 36.873 33.622 36.937 ;
			RECT	33.926 36.873 33.958 36.937 ;
			RECT	34.262 36.873 34.294 36.937 ;
			RECT	34.598 36.873 34.63 36.937 ;
			RECT	34.934 36.873 34.966 36.937 ;
			RECT	35.27 36.873 35.302 36.937 ;
			RECT	35.606 36.873 35.638 36.937 ;
			RECT	35.942 36.873 35.974 36.937 ;
			RECT	36.278 36.873 36.31 36.937 ;
			RECT	36.614 36.873 36.646 36.937 ;
			RECT	36.95 36.873 36.982 36.937 ;
			RECT	37.286 36.873 37.318 36.937 ;
			RECT	37.622 36.873 37.654 36.937 ;
			RECT	37.958 36.873 37.99 36.937 ;
			RECT	38.294 36.873 38.326 36.937 ;
			RECT	38.63 36.873 38.662 36.937 ;
			RECT	38.966 36.873 38.998 36.937 ;
			RECT	39.302 36.873 39.334 36.937 ;
			RECT	39.638 36.873 39.67 36.937 ;
			RECT	39.974 36.873 40.006 36.937 ;
			RECT	40.31 36.873 40.342 36.937 ;
			RECT	40.646 36.873 40.678 36.937 ;
			RECT	40.982 36.873 41.014 36.937 ;
			RECT	41.318 36.873 41.35 36.937 ;
			RECT	41.654 36.873 41.686 36.937 ;
			RECT	41.99 36.873 42.022 36.937 ;
			RECT	42.326 36.873 42.358 36.937 ;
			RECT	42.662 36.873 42.694 36.937 ;
			RECT	42.998 36.873 43.03 36.937 ;
			RECT	43.334 36.873 43.366 36.937 ;
			RECT	43.67 36.873 43.702 36.937 ;
			RECT	44.016 36.873 44.048 36.937 ;
			RECT	44.342 36.873 44.374 36.937 ;
			RECT	44.678 36.873 44.71 36.937 ;
			RECT	45.014 36.873 45.046 36.937 ;
			RECT	45.35 36.873 45.382 36.937 ;
			RECT	46.022 36.873 46.054 36.937 ;
			RECT	46.358 36.873 46.39 36.937 ;
			RECT	47.03 36.873 47.062 36.937 ;
			RECT	47.366 36.873 47.398 36.937 ;
			RECT	48.038 36.873 48.07 36.937 ;
			RECT	48.374 36.873 48.406 36.937 ;
			RECT	48.71 36.873 48.742 36.937 ;
			RECT	49.046 36.873 49.078 36.937 ;
			RECT	49.227 36.873 49.259 36.937 ;
			RECT	49.7 36.873 49.732 36.937 ;
			RECT	49.994 36.873 50.026 36.937 ;
			RECT	50.516 36.873 50.548 36.937 ;
			RECT	52.15 36.873 52.182 36.937 ;
			RECT	58.178 36.873 58.21 36.937 ;
			RECT	58.472 36.873 58.504 36.937 ;
			RECT	58.945 36.873 58.977 36.937 ;
			RECT	59.126 36.873 59.158 36.937 ;
			RECT	59.462 36.873 59.494 36.937 ;
			RECT	59.798 36.873 59.83 36.937 ;
			RECT	60.134 36.873 60.166 36.937 ;
			RECT	60.806 36.873 60.838 36.937 ;
			RECT	61.142 36.873 61.174 36.937 ;
			RECT	61.814 36.873 61.846 36.937 ;
			RECT	62.15 36.873 62.182 36.937 ;
			RECT	62.822 36.873 62.854 36.937 ;
			RECT	63.158 36.873 63.19 36.937 ;
			RECT	63.494 36.873 63.526 36.937 ;
			RECT	63.83 36.873 63.862 36.937 ;
			RECT	64.156 36.873 64.188 36.937 ;
			RECT	64.502 36.873 64.534 36.937 ;
			RECT	64.838 36.873 64.87 36.937 ;
			RECT	65.174 36.873 65.206 36.937 ;
			RECT	65.51 36.873 65.542 36.937 ;
			RECT	65.846 36.873 65.878 36.937 ;
			RECT	66.182 36.873 66.214 36.937 ;
			RECT	66.518 36.873 66.55 36.937 ;
			RECT	66.854 36.873 66.886 36.937 ;
			RECT	67.19 36.873 67.222 36.937 ;
			RECT	67.526 36.873 67.558 36.937 ;
			RECT	67.862 36.873 67.894 36.937 ;
			RECT	68.198 36.873 68.23 36.937 ;
			RECT	68.534 36.873 68.566 36.937 ;
			RECT	68.87 36.873 68.902 36.937 ;
			RECT	69.206 36.873 69.238 36.937 ;
			RECT	69.542 36.873 69.574 36.937 ;
			RECT	69.878 36.873 69.91 36.937 ;
			RECT	70.214 36.873 70.246 36.937 ;
			RECT	70.55 36.873 70.582 36.937 ;
			RECT	70.886 36.873 70.918 36.937 ;
			RECT	71.222 36.873 71.254 36.937 ;
			RECT	71.558 36.873 71.59 36.937 ;
			RECT	71.894 36.873 71.926 36.937 ;
			RECT	72.23 36.873 72.262 36.937 ;
			RECT	72.566 36.873 72.598 36.937 ;
			RECT	72.902 36.873 72.934 36.937 ;
			RECT	73.238 36.873 73.27 36.937 ;
			RECT	73.574 36.873 73.606 36.937 ;
			RECT	73.91 36.873 73.942 36.937 ;
			RECT	74.246 36.873 74.278 36.937 ;
			RECT	74.582 36.873 74.614 36.937 ;
			RECT	74.918 36.873 74.95 36.937 ;
			RECT	75.254 36.873 75.286 36.937 ;
			RECT	75.59 36.873 75.622 36.937 ;
			RECT	75.926 36.873 75.958 36.937 ;
			RECT	76.262 36.873 76.294 36.937 ;
			RECT	76.598 36.873 76.63 36.937 ;
			RECT	76.934 36.873 76.966 36.937 ;
			RECT	77.27 36.873 77.302 36.937 ;
			RECT	77.606 36.873 77.638 36.937 ;
			RECT	77.942 36.873 77.974 36.937 ;
			RECT	78.278 36.873 78.31 36.937 ;
			RECT	78.614 36.873 78.646 36.937 ;
			RECT	78.95 36.873 78.982 36.937 ;
			RECT	79.286 36.873 79.318 36.937 ;
			RECT	79.622 36.873 79.654 36.937 ;
			RECT	79.958 36.873 79.99 36.937 ;
			RECT	80.294 36.873 80.326 36.937 ;
			RECT	80.625 36.873 80.657 36.937 ;
			RECT	80.961 36.873 80.993 36.937 ;
			RECT	81.297 36.873 81.329 36.937 ;
			RECT	81.633 36.873 81.665 36.937 ;
			RECT	81.969 36.873 82.001 36.937 ;
			RECT	82.305 36.873 82.337 36.937 ;
			RECT	82.641 36.873 82.673 36.937 ;
			RECT	82.977 36.873 83.009 36.937 ;
			RECT	83.313 36.873 83.345 36.937 ;
			RECT	83.649 36.873 83.681 36.937 ;
			RECT	83.985 36.873 84.017 36.937 ;
			RECT	84.321 36.873 84.353 36.937 ;
			RECT	84.657 36.873 84.689 36.937 ;
			RECT	84.993 36.873 85.025 36.937 ;
			RECT	85.329 36.873 85.361 36.937 ;
			RECT	85.665 36.873 85.697 36.937 ;
			RECT	86.001 36.873 86.033 36.937 ;
			RECT	86.337 36.873 86.369 36.937 ;
			RECT	86.673 36.873 86.705 36.937 ;
			RECT	87.009 36.873 87.041 36.937 ;
			RECT	87.345 36.873 87.377 36.937 ;
			RECT	87.681 36.873 87.713 36.937 ;
			RECT	88.017 36.873 88.049 36.937 ;
			RECT	88.353 36.873 88.385 36.937 ;
			RECT	88.689 36.873 88.721 36.937 ;
			RECT	89.025 36.873 89.057 36.937 ;
			RECT	89.361 36.873 89.393 36.937 ;
			RECT	89.697 36.873 89.729 36.937 ;
			RECT	90.033 36.873 90.065 36.937 ;
			RECT	90.369 36.873 90.401 36.937 ;
			RECT	90.705 36.873 90.737 36.937 ;
			RECT	91.041 36.873 91.073 36.937 ;
			RECT	91.377 36.873 91.409 36.937 ;
			RECT	91.713 36.873 91.745 36.937 ;
			RECT	92.049 36.873 92.081 36.937 ;
			RECT	92.385 36.873 92.417 36.937 ;
			RECT	92.721 36.873 92.753 36.937 ;
			RECT	93.057 36.873 93.089 36.937 ;
			RECT	93.393 36.873 93.425 36.937 ;
			RECT	93.729 36.873 93.761 36.937 ;
			RECT	94.065 36.873 94.097 36.937 ;
			RECT	94.401 36.873 94.433 36.937 ;
			RECT	94.737 36.873 94.769 36.937 ;
			RECT	95.073 36.873 95.105 36.937 ;
			RECT	95.409 36.873 95.441 36.937 ;
			RECT	95.745 36.873 95.777 36.937 ;
			RECT	96.081 36.873 96.113 36.937 ;
			RECT	96.417 36.873 96.449 36.937 ;
			RECT	96.753 36.873 96.785 36.937 ;
			RECT	97.089 36.873 97.121 36.937 ;
			RECT	97.425 36.873 97.457 36.937 ;
			RECT	97.761 36.873 97.793 36.937 ;
			RECT	98.097 36.873 98.129 36.937 ;
			RECT	98.433 36.873 98.465 36.937 ;
			RECT	98.769 36.873 98.801 36.937 ;
			RECT	99.105 36.873 99.137 36.937 ;
			RECT	99.441 36.873 99.473 36.937 ;
			RECT	99.777 36.873 99.809 36.937 ;
			RECT	100.113 36.873 100.145 36.937 ;
			RECT	100.449 36.873 100.481 36.937 ;
			RECT	100.785 36.873 100.817 36.937 ;
			RECT	101.121 36.873 101.153 36.937 ;
			RECT	101.457 36.873 101.489 36.937 ;
			RECT	101.793 36.873 101.825 36.937 ;
			RECT	102.324 36.873 102.356 36.937 ;
			RECT	103.846 36.873 103.878 36.937 ;
			RECT	104.377 36.873 104.409 36.937 ;
			RECT	104.713 36.873 104.745 36.937 ;
			RECT	105.049 36.873 105.081 36.937 ;
			RECT	105.385 36.873 105.417 36.937 ;
			RECT	105.721 36.873 105.753 36.937 ;
			RECT	106.057 36.873 106.089 36.937 ;
			RECT	106.393 36.873 106.425 36.937 ;
			RECT	106.729 36.873 106.761 36.937 ;
			RECT	107.065 36.873 107.097 36.937 ;
			RECT	107.401 36.873 107.433 36.937 ;
			RECT	107.737 36.873 107.769 36.937 ;
			RECT	108.073 36.873 108.105 36.937 ;
			RECT	108.409 36.873 108.441 36.937 ;
			RECT	108.745 36.873 108.777 36.937 ;
			RECT	109.081 36.873 109.113 36.937 ;
			RECT	109.417 36.873 109.449 36.937 ;
			RECT	109.753 36.873 109.785 36.937 ;
			RECT	110.089 36.873 110.121 36.937 ;
			RECT	110.425 36.873 110.457 36.937 ;
			RECT	110.761 36.873 110.793 36.937 ;
			RECT	111.097 36.873 111.129 36.937 ;
			RECT	111.433 36.873 111.465 36.937 ;
			RECT	111.769 36.873 111.801 36.937 ;
			RECT	112.105 36.873 112.137 36.937 ;
			RECT	112.441 36.873 112.473 36.937 ;
			RECT	112.777 36.873 112.809 36.937 ;
			RECT	113.113 36.873 113.145 36.937 ;
			RECT	113.449 36.873 113.481 36.937 ;
			RECT	113.785 36.873 113.817 36.937 ;
			RECT	114.121 36.873 114.153 36.937 ;
			RECT	114.457 36.873 114.489 36.937 ;
			RECT	114.793 36.873 114.825 36.937 ;
			RECT	115.129 36.873 115.161 36.937 ;
			RECT	115.465 36.873 115.497 36.937 ;
			RECT	115.801 36.873 115.833 36.937 ;
			RECT	116.137 36.873 116.169 36.937 ;
			RECT	116.473 36.873 116.505 36.937 ;
			RECT	116.809 36.873 116.841 36.937 ;
			RECT	117.145 36.873 117.177 36.937 ;
			RECT	117.481 36.873 117.513 36.937 ;
			RECT	117.817 36.873 117.849 36.937 ;
			RECT	118.153 36.873 118.185 36.937 ;
			RECT	118.489 36.873 118.521 36.937 ;
			RECT	118.825 36.873 118.857 36.937 ;
			RECT	119.161 36.873 119.193 36.937 ;
			RECT	119.497 36.873 119.529 36.937 ;
			RECT	119.833 36.873 119.865 36.937 ;
			RECT	120.169 36.873 120.201 36.937 ;
			RECT	120.505 36.873 120.537 36.937 ;
			RECT	120.841 36.873 120.873 36.937 ;
			RECT	121.177 36.873 121.209 36.937 ;
			RECT	121.513 36.873 121.545 36.937 ;
			RECT	121.849 36.873 121.881 36.937 ;
			RECT	122.185 36.873 122.217 36.937 ;
			RECT	122.521 36.873 122.553 36.937 ;
			RECT	122.857 36.873 122.889 36.937 ;
			RECT	123.193 36.873 123.225 36.937 ;
			RECT	123.529 36.873 123.561 36.937 ;
			RECT	123.865 36.873 123.897 36.937 ;
			RECT	124.201 36.873 124.233 36.937 ;
			RECT	124.537 36.873 124.569 36.937 ;
			RECT	124.873 36.873 124.905 36.937 ;
			RECT	125.209 36.873 125.241 36.937 ;
			RECT	125.545 36.873 125.577 36.937 ;
			RECT	125.876 36.873 125.908 36.937 ;
			RECT	126.212 36.873 126.244 36.937 ;
			RECT	126.548 36.873 126.58 36.937 ;
			RECT	126.884 36.873 126.916 36.937 ;
			RECT	127.22 36.873 127.252 36.937 ;
			RECT	127.556 36.873 127.588 36.937 ;
			RECT	127.892 36.873 127.924 36.937 ;
			RECT	128.228 36.873 128.26 36.937 ;
			RECT	128.564 36.873 128.596 36.937 ;
			RECT	128.9 36.873 128.932 36.937 ;
			RECT	129.236 36.873 129.268 36.937 ;
			RECT	129.572 36.873 129.604 36.937 ;
			RECT	129.908 36.873 129.94 36.937 ;
			RECT	130.244 36.873 130.276 36.937 ;
			RECT	130.58 36.873 130.612 36.937 ;
			RECT	130.916 36.873 130.948 36.937 ;
			RECT	131.252 36.873 131.284 36.937 ;
			RECT	131.588 36.873 131.62 36.937 ;
			RECT	131.924 36.873 131.956 36.937 ;
			RECT	132.26 36.873 132.292 36.937 ;
			RECT	132.596 36.873 132.628 36.937 ;
			RECT	132.932 36.873 132.964 36.937 ;
			RECT	133.268 36.873 133.3 36.937 ;
			RECT	133.604 36.873 133.636 36.937 ;
			RECT	133.94 36.873 133.972 36.937 ;
			RECT	134.276 36.873 134.308 36.937 ;
			RECT	134.612 36.873 134.644 36.937 ;
			RECT	134.948 36.873 134.98 36.937 ;
			RECT	135.284 36.873 135.316 36.937 ;
			RECT	135.62 36.873 135.652 36.937 ;
			RECT	135.956 36.873 135.988 36.937 ;
			RECT	136.292 36.873 136.324 36.937 ;
			RECT	136.628 36.873 136.66 36.937 ;
			RECT	136.964 36.873 136.996 36.937 ;
			RECT	137.3 36.873 137.332 36.937 ;
			RECT	137.636 36.873 137.668 36.937 ;
			RECT	137.972 36.873 138.004 36.937 ;
			RECT	138.308 36.873 138.34 36.937 ;
			RECT	138.644 36.873 138.676 36.937 ;
			RECT	138.98 36.873 139.012 36.937 ;
			RECT	139.316 36.873 139.348 36.937 ;
			RECT	139.652 36.873 139.684 36.937 ;
			RECT	139.988 36.873 140.02 36.937 ;
			RECT	140.324 36.873 140.356 36.937 ;
			RECT	140.66 36.873 140.692 36.937 ;
			RECT	140.996 36.873 141.028 36.937 ;
			RECT	141.332 36.873 141.364 36.937 ;
			RECT	141.668 36.873 141.7 36.937 ;
			RECT	142.014 36.873 142.046 36.937 ;
			RECT	142.34 36.873 142.372 36.937 ;
			RECT	142.676 36.873 142.708 36.937 ;
			RECT	143.012 36.873 143.044 36.937 ;
			RECT	143.348 36.873 143.38 36.937 ;
			RECT	144.02 36.873 144.052 36.937 ;
			RECT	144.356 36.873 144.388 36.937 ;
			RECT	145.028 36.873 145.06 36.937 ;
			RECT	145.364 36.873 145.396 36.937 ;
			RECT	146.036 36.873 146.068 36.937 ;
			RECT	146.372 36.873 146.404 36.937 ;
			RECT	146.708 36.873 146.74 36.937 ;
			RECT	147.044 36.873 147.076 36.937 ;
			RECT	147.225 36.873 147.257 36.937 ;
			RECT	147.698 36.873 147.73 36.937 ;
			RECT	147.992 36.873 148.024 36.937 ;
			RECT	148.514 36.873 148.546 36.937 ;
			RECT	150.148 36.873 150.18 36.937 ;
			RECT	156.176 36.873 156.208 36.937 ;
			RECT	156.47 36.873 156.502 36.937 ;
			RECT	156.943 36.873 156.975 36.937 ;
			RECT	157.124 36.873 157.156 36.937 ;
			RECT	157.46 36.873 157.492 36.937 ;
			RECT	157.796 36.873 157.828 36.937 ;
			RECT	158.132 36.873 158.164 36.937 ;
			RECT	158.804 36.873 158.836 36.937 ;
			RECT	159.14 36.873 159.172 36.937 ;
			RECT	159.812 36.873 159.844 36.937 ;
			RECT	160.148 36.873 160.18 36.937 ;
			RECT	160.82 36.873 160.852 36.937 ;
			RECT	161.156 36.873 161.188 36.937 ;
			RECT	161.492 36.873 161.524 36.937 ;
			RECT	161.828 36.873 161.86 36.937 ;
			RECT	162.154 36.873 162.186 36.937 ;
			RECT	162.5 36.873 162.532 36.937 ;
			RECT	162.836 36.873 162.868 36.937 ;
			RECT	163.172 36.873 163.204 36.937 ;
			RECT	163.508 36.873 163.54 36.937 ;
			RECT	163.844 36.873 163.876 36.937 ;
			RECT	164.18 36.873 164.212 36.937 ;
			RECT	164.516 36.873 164.548 36.937 ;
			RECT	164.852 36.873 164.884 36.937 ;
			RECT	165.188 36.873 165.22 36.937 ;
			RECT	165.524 36.873 165.556 36.937 ;
			RECT	165.86 36.873 165.892 36.937 ;
			RECT	166.196 36.873 166.228 36.937 ;
			RECT	166.532 36.873 166.564 36.937 ;
			RECT	166.868 36.873 166.9 36.937 ;
			RECT	167.204 36.873 167.236 36.937 ;
			RECT	167.54 36.873 167.572 36.937 ;
			RECT	167.876 36.873 167.908 36.937 ;
			RECT	168.212 36.873 168.244 36.937 ;
			RECT	168.548 36.873 168.58 36.937 ;
			RECT	168.884 36.873 168.916 36.937 ;
			RECT	169.22 36.873 169.252 36.937 ;
			RECT	169.556 36.873 169.588 36.937 ;
			RECT	169.892 36.873 169.924 36.937 ;
			RECT	170.228 36.873 170.26 36.937 ;
			RECT	170.564 36.873 170.596 36.937 ;
			RECT	170.9 36.873 170.932 36.937 ;
			RECT	171.236 36.873 171.268 36.937 ;
			RECT	171.572 36.873 171.604 36.937 ;
			RECT	171.908 36.873 171.94 36.937 ;
			RECT	172.244 36.873 172.276 36.937 ;
			RECT	172.58 36.873 172.612 36.937 ;
			RECT	172.916 36.873 172.948 36.937 ;
			RECT	173.252 36.873 173.284 36.937 ;
			RECT	173.588 36.873 173.62 36.937 ;
			RECT	173.924 36.873 173.956 36.937 ;
			RECT	174.26 36.873 174.292 36.937 ;
			RECT	174.596 36.873 174.628 36.937 ;
			RECT	174.932 36.873 174.964 36.937 ;
			RECT	175.268 36.873 175.3 36.937 ;
			RECT	175.604 36.873 175.636 36.937 ;
			RECT	175.94 36.873 175.972 36.937 ;
			RECT	176.276 36.873 176.308 36.937 ;
			RECT	176.612 36.873 176.644 36.937 ;
			RECT	176.948 36.873 176.98 36.937 ;
			RECT	177.284 36.873 177.316 36.937 ;
			RECT	177.62 36.873 177.652 36.937 ;
			RECT	177.956 36.873 177.988 36.937 ;
			RECT	178.292 36.873 178.324 36.937 ;
			RECT	178.623 36.873 178.655 36.937 ;
			RECT	178.959 36.873 178.991 36.937 ;
			RECT	179.295 36.873 179.327 36.937 ;
			RECT	179.631 36.873 179.663 36.937 ;
			RECT	179.967 36.873 179.999 36.937 ;
			RECT	180.303 36.873 180.335 36.937 ;
			RECT	180.639 36.873 180.671 36.937 ;
			RECT	180.975 36.873 181.007 36.937 ;
			RECT	181.311 36.873 181.343 36.937 ;
			RECT	181.647 36.873 181.679 36.937 ;
			RECT	181.983 36.873 182.015 36.937 ;
			RECT	182.319 36.873 182.351 36.937 ;
			RECT	182.655 36.873 182.687 36.937 ;
			RECT	182.991 36.873 183.023 36.937 ;
			RECT	183.327 36.873 183.359 36.937 ;
			RECT	183.663 36.873 183.695 36.937 ;
			RECT	183.999 36.873 184.031 36.937 ;
			RECT	184.335 36.873 184.367 36.937 ;
			RECT	184.671 36.873 184.703 36.937 ;
			RECT	185.007 36.873 185.039 36.937 ;
			RECT	185.343 36.873 185.375 36.937 ;
			RECT	185.679 36.873 185.711 36.937 ;
			RECT	186.015 36.873 186.047 36.937 ;
			RECT	186.351 36.873 186.383 36.937 ;
			RECT	186.687 36.873 186.719 36.937 ;
			RECT	187.023 36.873 187.055 36.937 ;
			RECT	187.359 36.873 187.391 36.937 ;
			RECT	187.695 36.873 187.727 36.937 ;
			RECT	188.031 36.873 188.063 36.937 ;
			RECT	188.367 36.873 188.399 36.937 ;
			RECT	188.703 36.873 188.735 36.937 ;
			RECT	189.039 36.873 189.071 36.937 ;
			RECT	189.375 36.873 189.407 36.937 ;
			RECT	189.711 36.873 189.743 36.937 ;
			RECT	190.047 36.873 190.079 36.937 ;
			RECT	190.383 36.873 190.415 36.937 ;
			RECT	190.719 36.873 190.751 36.937 ;
			RECT	191.055 36.873 191.087 36.937 ;
			RECT	191.391 36.873 191.423 36.937 ;
			RECT	191.727 36.873 191.759 36.937 ;
			RECT	192.063 36.873 192.095 36.937 ;
			RECT	192.399 36.873 192.431 36.937 ;
			RECT	192.735 36.873 192.767 36.937 ;
			RECT	193.071 36.873 193.103 36.937 ;
			RECT	193.407 36.873 193.439 36.937 ;
			RECT	193.743 36.873 193.775 36.937 ;
			RECT	194.079 36.873 194.111 36.937 ;
			RECT	194.415 36.873 194.447 36.937 ;
			RECT	194.751 36.873 194.783 36.937 ;
			RECT	195.087 36.873 195.119 36.937 ;
			RECT	195.423 36.873 195.455 36.937 ;
			RECT	195.759 36.873 195.791 36.937 ;
			RECT	196.095 36.873 196.127 36.937 ;
			RECT	196.431 36.873 196.463 36.937 ;
			RECT	196.767 36.873 196.799 36.937 ;
			RECT	197.103 36.873 197.135 36.937 ;
			RECT	197.439 36.873 197.471 36.937 ;
			RECT	197.775 36.873 197.807 36.937 ;
			RECT	198.111 36.873 198.143 36.937 ;
			RECT	198.447 36.873 198.479 36.937 ;
			RECT	198.783 36.873 198.815 36.937 ;
			RECT	199.119 36.873 199.151 36.937 ;
			RECT	199.455 36.873 199.487 36.937 ;
			RECT	199.791 36.873 199.823 36.937 ;
			RECT	200.322 36.873 200.354 36.937 ;
			RECT	201.14 36.873 201.204 36.937 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 41.656 201.665 41.776 ;
			LAYER	J3 ;
			RECT	5.848 41.684 5.88 41.748 ;
			RECT	45.35 41.684 45.382 41.748 ;
			RECT	45.696 41.684 45.728 41.748 ;
			RECT	62.476 41.684 62.508 41.748 ;
			RECT	62.822 41.684 62.854 41.748 ;
			RECT	102.324 41.684 102.356 41.748 ;
			RECT	103.846 41.684 103.878 41.748 ;
			RECT	143.348 41.684 143.38 41.748 ;
			RECT	143.694 41.684 143.726 41.748 ;
			RECT	160.474 41.684 160.506 41.748 ;
			RECT	160.82 41.684 160.852 41.748 ;
			RECT	200.322 41.684 200.354 41.748 ;
			RECT	201.14 41.684 201.204 41.748 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 45.423 201.665 45.543 ;
			LAYER	J3 ;
			RECT	5.064 45.451 5.096 45.515 ;
			RECT	6.379 45.451 6.411 45.515 ;
			RECT	6.715 45.451 6.747 45.515 ;
			RECT	7.051 45.451 7.083 45.515 ;
			RECT	7.387 45.451 7.419 45.515 ;
			RECT	7.723 45.451 7.755 45.515 ;
			RECT	8.059 45.451 8.091 45.515 ;
			RECT	8.395 45.451 8.427 45.515 ;
			RECT	8.731 45.451 8.763 45.515 ;
			RECT	9.067 45.451 9.099 45.515 ;
			RECT	9.403 45.451 9.435 45.515 ;
			RECT	9.739 45.451 9.771 45.515 ;
			RECT	10.075 45.451 10.107 45.515 ;
			RECT	10.411 45.451 10.443 45.515 ;
			RECT	10.747 45.451 10.779 45.515 ;
			RECT	11.083 45.451 11.115 45.515 ;
			RECT	11.419 45.451 11.451 45.515 ;
			RECT	11.755 45.451 11.787 45.515 ;
			RECT	12.091 45.451 12.123 45.515 ;
			RECT	12.427 45.451 12.459 45.515 ;
			RECT	12.763 45.451 12.795 45.515 ;
			RECT	13.099 45.451 13.131 45.515 ;
			RECT	13.435 45.451 13.467 45.515 ;
			RECT	13.771 45.451 13.803 45.515 ;
			RECT	14.107 45.451 14.139 45.515 ;
			RECT	14.443 45.451 14.475 45.515 ;
			RECT	14.779 45.451 14.811 45.515 ;
			RECT	15.115 45.451 15.147 45.515 ;
			RECT	15.451 45.451 15.483 45.515 ;
			RECT	15.787 45.451 15.819 45.515 ;
			RECT	16.123 45.451 16.155 45.515 ;
			RECT	16.459 45.451 16.491 45.515 ;
			RECT	16.795 45.451 16.827 45.515 ;
			RECT	17.131 45.451 17.163 45.515 ;
			RECT	17.467 45.451 17.499 45.515 ;
			RECT	17.803 45.451 17.835 45.515 ;
			RECT	18.139 45.451 18.171 45.515 ;
			RECT	18.475 45.451 18.507 45.515 ;
			RECT	18.811 45.451 18.843 45.515 ;
			RECT	19.147 45.451 19.179 45.515 ;
			RECT	19.483 45.451 19.515 45.515 ;
			RECT	19.819 45.451 19.851 45.515 ;
			RECT	20.155 45.451 20.187 45.515 ;
			RECT	20.491 45.451 20.523 45.515 ;
			RECT	20.827 45.451 20.859 45.515 ;
			RECT	21.163 45.451 21.195 45.515 ;
			RECT	21.499 45.451 21.531 45.515 ;
			RECT	21.835 45.451 21.867 45.515 ;
			RECT	22.171 45.451 22.203 45.515 ;
			RECT	22.507 45.451 22.539 45.515 ;
			RECT	22.843 45.451 22.875 45.515 ;
			RECT	23.179 45.451 23.211 45.515 ;
			RECT	23.515 45.451 23.547 45.515 ;
			RECT	23.851 45.451 23.883 45.515 ;
			RECT	24.187 45.451 24.219 45.515 ;
			RECT	24.523 45.451 24.555 45.515 ;
			RECT	24.859 45.451 24.891 45.515 ;
			RECT	25.195 45.451 25.227 45.515 ;
			RECT	25.531 45.451 25.563 45.515 ;
			RECT	25.867 45.451 25.899 45.515 ;
			RECT	26.203 45.451 26.235 45.515 ;
			RECT	26.539 45.451 26.571 45.515 ;
			RECT	26.875 45.451 26.907 45.515 ;
			RECT	27.211 45.451 27.243 45.515 ;
			RECT	27.547 45.451 27.579 45.515 ;
			RECT	27.878 45.451 27.91 45.515 ;
			RECT	28.214 45.451 28.246 45.515 ;
			RECT	28.55 45.451 28.582 45.515 ;
			RECT	28.886 45.451 28.918 45.515 ;
			RECT	29.222 45.451 29.254 45.515 ;
			RECT	29.558 45.451 29.59 45.515 ;
			RECT	29.894 45.451 29.926 45.515 ;
			RECT	30.23 45.451 30.262 45.515 ;
			RECT	30.566 45.451 30.598 45.515 ;
			RECT	30.902 45.451 30.934 45.515 ;
			RECT	31.238 45.451 31.27 45.515 ;
			RECT	31.574 45.451 31.606 45.515 ;
			RECT	31.91 45.451 31.942 45.515 ;
			RECT	32.246 45.451 32.278 45.515 ;
			RECT	32.582 45.451 32.614 45.515 ;
			RECT	32.918 45.451 32.95 45.515 ;
			RECT	33.254 45.451 33.286 45.515 ;
			RECT	33.59 45.451 33.622 45.515 ;
			RECT	33.926 45.451 33.958 45.515 ;
			RECT	34.262 45.451 34.294 45.515 ;
			RECT	34.598 45.451 34.63 45.515 ;
			RECT	34.934 45.451 34.966 45.515 ;
			RECT	35.27 45.451 35.302 45.515 ;
			RECT	35.606 45.451 35.638 45.515 ;
			RECT	35.942 45.451 35.974 45.515 ;
			RECT	36.278 45.451 36.31 45.515 ;
			RECT	36.614 45.451 36.646 45.515 ;
			RECT	36.95 45.451 36.982 45.515 ;
			RECT	37.286 45.451 37.318 45.515 ;
			RECT	37.622 45.451 37.654 45.515 ;
			RECT	37.958 45.451 37.99 45.515 ;
			RECT	38.294 45.451 38.326 45.515 ;
			RECT	38.63 45.451 38.662 45.515 ;
			RECT	38.966 45.451 38.998 45.515 ;
			RECT	39.302 45.451 39.334 45.515 ;
			RECT	39.638 45.451 39.67 45.515 ;
			RECT	39.974 45.451 40.006 45.515 ;
			RECT	40.31 45.451 40.342 45.515 ;
			RECT	40.646 45.451 40.678 45.515 ;
			RECT	40.982 45.451 41.014 45.515 ;
			RECT	41.318 45.451 41.35 45.515 ;
			RECT	41.654 45.451 41.686 45.515 ;
			RECT	41.99 45.451 42.022 45.515 ;
			RECT	42.326 45.451 42.358 45.515 ;
			RECT	42.662 45.451 42.694 45.515 ;
			RECT	42.998 45.451 43.03 45.515 ;
			RECT	43.334 45.451 43.366 45.515 ;
			RECT	43.67 45.451 43.702 45.515 ;
			RECT	44.016 45.451 44.048 45.515 ;
			RECT	44.342 45.451 44.374 45.515 ;
			RECT	44.678 45.451 44.71 45.515 ;
			RECT	45.014 45.451 45.046 45.515 ;
			RECT	45.35 45.451 45.382 45.515 ;
			RECT	45.686 45.451 45.718 45.515 ;
			RECT	46.022 45.451 46.054 45.515 ;
			RECT	46.358 45.451 46.39 45.515 ;
			RECT	46.694 45.451 46.726 45.515 ;
			RECT	47.03 45.451 47.062 45.515 ;
			RECT	47.366 45.451 47.398 45.515 ;
			RECT	47.702 45.451 47.734 45.515 ;
			RECT	48.038 45.451 48.07 45.515 ;
			RECT	48.374 45.451 48.406 45.515 ;
			RECT	48.71 45.451 48.742 45.515 ;
			RECT	49.046 45.451 49.078 45.515 ;
			RECT	49.691 45.451 49.723 45.515 ;
			RECT	52.121 45.451 52.153 45.515 ;
			RECT	58.481 45.451 58.513 45.515 ;
			RECT	59.126 45.451 59.158 45.515 ;
			RECT	59.462 45.451 59.494 45.515 ;
			RECT	59.798 45.451 59.83 45.515 ;
			RECT	60.134 45.451 60.166 45.515 ;
			RECT	60.47 45.451 60.502 45.515 ;
			RECT	60.806 45.451 60.838 45.515 ;
			RECT	61.142 45.451 61.174 45.515 ;
			RECT	61.478 45.451 61.51 45.515 ;
			RECT	61.814 45.451 61.846 45.515 ;
			RECT	62.15 45.451 62.182 45.515 ;
			RECT	62.486 45.451 62.518 45.515 ;
			RECT	62.822 45.451 62.854 45.515 ;
			RECT	63.158 45.451 63.19 45.515 ;
			RECT	63.494 45.451 63.526 45.515 ;
			RECT	63.83 45.451 63.862 45.515 ;
			RECT	64.156 45.451 64.188 45.515 ;
			RECT	64.502 45.451 64.534 45.515 ;
			RECT	64.838 45.451 64.87 45.515 ;
			RECT	65.174 45.451 65.206 45.515 ;
			RECT	65.51 45.451 65.542 45.515 ;
			RECT	65.846 45.451 65.878 45.515 ;
			RECT	66.182 45.451 66.214 45.515 ;
			RECT	66.518 45.451 66.55 45.515 ;
			RECT	66.854 45.451 66.886 45.515 ;
			RECT	67.19 45.451 67.222 45.515 ;
			RECT	67.526 45.451 67.558 45.515 ;
			RECT	67.862 45.451 67.894 45.515 ;
			RECT	68.198 45.451 68.23 45.515 ;
			RECT	68.534 45.451 68.566 45.515 ;
			RECT	68.87 45.451 68.902 45.515 ;
			RECT	69.206 45.451 69.238 45.515 ;
			RECT	69.542 45.451 69.574 45.515 ;
			RECT	69.878 45.451 69.91 45.515 ;
			RECT	70.214 45.451 70.246 45.515 ;
			RECT	70.55 45.451 70.582 45.515 ;
			RECT	70.886 45.451 70.918 45.515 ;
			RECT	71.222 45.451 71.254 45.515 ;
			RECT	71.558 45.451 71.59 45.515 ;
			RECT	71.894 45.451 71.926 45.515 ;
			RECT	72.23 45.451 72.262 45.515 ;
			RECT	72.566 45.451 72.598 45.515 ;
			RECT	72.902 45.451 72.934 45.515 ;
			RECT	73.238 45.451 73.27 45.515 ;
			RECT	73.574 45.451 73.606 45.515 ;
			RECT	73.91 45.451 73.942 45.515 ;
			RECT	74.246 45.451 74.278 45.515 ;
			RECT	74.582 45.451 74.614 45.515 ;
			RECT	74.918 45.451 74.95 45.515 ;
			RECT	75.254 45.451 75.286 45.515 ;
			RECT	75.59 45.451 75.622 45.515 ;
			RECT	75.926 45.451 75.958 45.515 ;
			RECT	76.262 45.451 76.294 45.515 ;
			RECT	76.598 45.451 76.63 45.515 ;
			RECT	76.934 45.451 76.966 45.515 ;
			RECT	77.27 45.451 77.302 45.515 ;
			RECT	77.606 45.451 77.638 45.515 ;
			RECT	77.942 45.451 77.974 45.515 ;
			RECT	78.278 45.451 78.31 45.515 ;
			RECT	78.614 45.451 78.646 45.515 ;
			RECT	78.95 45.451 78.982 45.515 ;
			RECT	79.286 45.451 79.318 45.515 ;
			RECT	79.622 45.451 79.654 45.515 ;
			RECT	79.958 45.451 79.99 45.515 ;
			RECT	80.294 45.451 80.326 45.515 ;
			RECT	80.625 45.451 80.657 45.515 ;
			RECT	80.961 45.451 80.993 45.515 ;
			RECT	81.297 45.451 81.329 45.515 ;
			RECT	81.633 45.451 81.665 45.515 ;
			RECT	81.969 45.451 82.001 45.515 ;
			RECT	82.305 45.451 82.337 45.515 ;
			RECT	82.641 45.451 82.673 45.515 ;
			RECT	82.977 45.451 83.009 45.515 ;
			RECT	83.313 45.451 83.345 45.515 ;
			RECT	83.649 45.451 83.681 45.515 ;
			RECT	83.985 45.451 84.017 45.515 ;
			RECT	84.321 45.451 84.353 45.515 ;
			RECT	84.657 45.451 84.689 45.515 ;
			RECT	84.993 45.451 85.025 45.515 ;
			RECT	85.329 45.451 85.361 45.515 ;
			RECT	85.665 45.451 85.697 45.515 ;
			RECT	86.001 45.451 86.033 45.515 ;
			RECT	86.337 45.451 86.369 45.515 ;
			RECT	86.673 45.451 86.705 45.515 ;
			RECT	87.009 45.451 87.041 45.515 ;
			RECT	87.345 45.451 87.377 45.515 ;
			RECT	87.681 45.451 87.713 45.515 ;
			RECT	88.017 45.451 88.049 45.515 ;
			RECT	88.353 45.451 88.385 45.515 ;
			RECT	88.689 45.451 88.721 45.515 ;
			RECT	89.025 45.451 89.057 45.515 ;
			RECT	89.361 45.451 89.393 45.515 ;
			RECT	89.697 45.451 89.729 45.515 ;
			RECT	90.033 45.451 90.065 45.515 ;
			RECT	90.369 45.451 90.401 45.515 ;
			RECT	90.705 45.451 90.737 45.515 ;
			RECT	91.041 45.451 91.073 45.515 ;
			RECT	91.377 45.451 91.409 45.515 ;
			RECT	91.713 45.451 91.745 45.515 ;
			RECT	92.049 45.451 92.081 45.515 ;
			RECT	92.385 45.451 92.417 45.515 ;
			RECT	92.721 45.451 92.753 45.515 ;
			RECT	93.057 45.451 93.089 45.515 ;
			RECT	93.393 45.451 93.425 45.515 ;
			RECT	93.729 45.451 93.761 45.515 ;
			RECT	94.065 45.451 94.097 45.515 ;
			RECT	94.401 45.451 94.433 45.515 ;
			RECT	94.737 45.451 94.769 45.515 ;
			RECT	95.073 45.451 95.105 45.515 ;
			RECT	95.409 45.451 95.441 45.515 ;
			RECT	95.745 45.451 95.777 45.515 ;
			RECT	96.081 45.451 96.113 45.515 ;
			RECT	96.417 45.451 96.449 45.515 ;
			RECT	96.753 45.451 96.785 45.515 ;
			RECT	97.089 45.451 97.121 45.515 ;
			RECT	97.425 45.451 97.457 45.515 ;
			RECT	97.761 45.451 97.793 45.515 ;
			RECT	98.097 45.451 98.129 45.515 ;
			RECT	98.433 45.451 98.465 45.515 ;
			RECT	98.769 45.451 98.801 45.515 ;
			RECT	99.105 45.451 99.137 45.515 ;
			RECT	99.441 45.451 99.473 45.515 ;
			RECT	99.777 45.451 99.809 45.515 ;
			RECT	100.113 45.451 100.145 45.515 ;
			RECT	100.449 45.451 100.481 45.515 ;
			RECT	100.785 45.451 100.817 45.515 ;
			RECT	101.121 45.451 101.153 45.515 ;
			RECT	101.457 45.451 101.489 45.515 ;
			RECT	101.793 45.451 101.825 45.515 ;
			RECT	104.377 45.451 104.409 45.515 ;
			RECT	104.713 45.451 104.745 45.515 ;
			RECT	105.049 45.451 105.081 45.515 ;
			RECT	105.385 45.451 105.417 45.515 ;
			RECT	105.721 45.451 105.753 45.515 ;
			RECT	106.057 45.451 106.089 45.515 ;
			RECT	106.393 45.451 106.425 45.515 ;
			RECT	106.729 45.451 106.761 45.515 ;
			RECT	107.065 45.451 107.097 45.515 ;
			RECT	107.401 45.451 107.433 45.515 ;
			RECT	107.737 45.451 107.769 45.515 ;
			RECT	108.073 45.451 108.105 45.515 ;
			RECT	108.409 45.451 108.441 45.515 ;
			RECT	108.745 45.451 108.777 45.515 ;
			RECT	109.081 45.451 109.113 45.515 ;
			RECT	109.417 45.451 109.449 45.515 ;
			RECT	109.753 45.451 109.785 45.515 ;
			RECT	110.089 45.451 110.121 45.515 ;
			RECT	110.425 45.451 110.457 45.515 ;
			RECT	110.761 45.451 110.793 45.515 ;
			RECT	111.097 45.451 111.129 45.515 ;
			RECT	111.433 45.451 111.465 45.515 ;
			RECT	111.769 45.451 111.801 45.515 ;
			RECT	112.105 45.451 112.137 45.515 ;
			RECT	112.441 45.451 112.473 45.515 ;
			RECT	112.777 45.451 112.809 45.515 ;
			RECT	113.113 45.451 113.145 45.515 ;
			RECT	113.449 45.451 113.481 45.515 ;
			RECT	113.785 45.451 113.817 45.515 ;
			RECT	114.121 45.451 114.153 45.515 ;
			RECT	114.457 45.451 114.489 45.515 ;
			RECT	114.793 45.451 114.825 45.515 ;
			RECT	115.129 45.451 115.161 45.515 ;
			RECT	115.465 45.451 115.497 45.515 ;
			RECT	115.801 45.451 115.833 45.515 ;
			RECT	116.137 45.451 116.169 45.515 ;
			RECT	116.473 45.451 116.505 45.515 ;
			RECT	116.809 45.451 116.841 45.515 ;
			RECT	117.145 45.451 117.177 45.515 ;
			RECT	117.481 45.451 117.513 45.515 ;
			RECT	117.817 45.451 117.849 45.515 ;
			RECT	118.153 45.451 118.185 45.515 ;
			RECT	118.489 45.451 118.521 45.515 ;
			RECT	118.825 45.451 118.857 45.515 ;
			RECT	119.161 45.451 119.193 45.515 ;
			RECT	119.497 45.451 119.529 45.515 ;
			RECT	119.833 45.451 119.865 45.515 ;
			RECT	120.169 45.451 120.201 45.515 ;
			RECT	120.505 45.451 120.537 45.515 ;
			RECT	120.841 45.451 120.873 45.515 ;
			RECT	121.177 45.451 121.209 45.515 ;
			RECT	121.513 45.451 121.545 45.515 ;
			RECT	121.849 45.451 121.881 45.515 ;
			RECT	122.185 45.451 122.217 45.515 ;
			RECT	122.521 45.451 122.553 45.515 ;
			RECT	122.857 45.451 122.889 45.515 ;
			RECT	123.193 45.451 123.225 45.515 ;
			RECT	123.529 45.451 123.561 45.515 ;
			RECT	123.865 45.451 123.897 45.515 ;
			RECT	124.201 45.451 124.233 45.515 ;
			RECT	124.537 45.451 124.569 45.515 ;
			RECT	124.873 45.451 124.905 45.515 ;
			RECT	125.209 45.451 125.241 45.515 ;
			RECT	125.545 45.451 125.577 45.515 ;
			RECT	125.876 45.451 125.908 45.515 ;
			RECT	126.212 45.451 126.244 45.515 ;
			RECT	126.548 45.451 126.58 45.515 ;
			RECT	126.884 45.451 126.916 45.515 ;
			RECT	127.22 45.451 127.252 45.515 ;
			RECT	127.556 45.451 127.588 45.515 ;
			RECT	127.892 45.451 127.924 45.515 ;
			RECT	128.228 45.451 128.26 45.515 ;
			RECT	128.564 45.451 128.596 45.515 ;
			RECT	128.9 45.451 128.932 45.515 ;
			RECT	129.236 45.451 129.268 45.515 ;
			RECT	129.572 45.451 129.604 45.515 ;
			RECT	129.908 45.451 129.94 45.515 ;
			RECT	130.244 45.451 130.276 45.515 ;
			RECT	130.58 45.451 130.612 45.515 ;
			RECT	130.916 45.451 130.948 45.515 ;
			RECT	131.252 45.451 131.284 45.515 ;
			RECT	131.588 45.451 131.62 45.515 ;
			RECT	131.924 45.451 131.956 45.515 ;
			RECT	132.26 45.451 132.292 45.515 ;
			RECT	132.596 45.451 132.628 45.515 ;
			RECT	132.932 45.451 132.964 45.515 ;
			RECT	133.268 45.451 133.3 45.515 ;
			RECT	133.604 45.451 133.636 45.515 ;
			RECT	133.94 45.451 133.972 45.515 ;
			RECT	134.276 45.451 134.308 45.515 ;
			RECT	134.612 45.451 134.644 45.515 ;
			RECT	134.948 45.451 134.98 45.515 ;
			RECT	135.284 45.451 135.316 45.515 ;
			RECT	135.62 45.451 135.652 45.515 ;
			RECT	135.956 45.451 135.988 45.515 ;
			RECT	136.292 45.451 136.324 45.515 ;
			RECT	136.628 45.451 136.66 45.515 ;
			RECT	136.964 45.451 136.996 45.515 ;
			RECT	137.3 45.451 137.332 45.515 ;
			RECT	137.636 45.451 137.668 45.515 ;
			RECT	137.972 45.451 138.004 45.515 ;
			RECT	138.308 45.451 138.34 45.515 ;
			RECT	138.644 45.451 138.676 45.515 ;
			RECT	138.98 45.451 139.012 45.515 ;
			RECT	139.316 45.451 139.348 45.515 ;
			RECT	139.652 45.451 139.684 45.515 ;
			RECT	139.988 45.451 140.02 45.515 ;
			RECT	140.324 45.451 140.356 45.515 ;
			RECT	140.66 45.451 140.692 45.515 ;
			RECT	140.996 45.451 141.028 45.515 ;
			RECT	141.332 45.451 141.364 45.515 ;
			RECT	141.668 45.451 141.7 45.515 ;
			RECT	142.014 45.451 142.046 45.515 ;
			RECT	142.34 45.451 142.372 45.515 ;
			RECT	142.676 45.451 142.708 45.515 ;
			RECT	143.012 45.451 143.044 45.515 ;
			RECT	143.348 45.451 143.38 45.515 ;
			RECT	143.684 45.451 143.716 45.515 ;
			RECT	144.02 45.451 144.052 45.515 ;
			RECT	144.356 45.451 144.388 45.515 ;
			RECT	144.692 45.451 144.724 45.515 ;
			RECT	145.028 45.451 145.06 45.515 ;
			RECT	145.364 45.451 145.396 45.515 ;
			RECT	145.7 45.451 145.732 45.515 ;
			RECT	146.036 45.451 146.068 45.515 ;
			RECT	146.372 45.451 146.404 45.515 ;
			RECT	146.708 45.451 146.74 45.515 ;
			RECT	147.044 45.451 147.076 45.515 ;
			RECT	147.689 45.451 147.721 45.515 ;
			RECT	150.119 45.451 150.151 45.515 ;
			RECT	156.479 45.451 156.511 45.515 ;
			RECT	157.124 45.451 157.156 45.515 ;
			RECT	157.46 45.451 157.492 45.515 ;
			RECT	157.796 45.451 157.828 45.515 ;
			RECT	158.132 45.451 158.164 45.515 ;
			RECT	158.468 45.451 158.5 45.515 ;
			RECT	158.804 45.451 158.836 45.515 ;
			RECT	159.14 45.451 159.172 45.515 ;
			RECT	159.476 45.451 159.508 45.515 ;
			RECT	159.812 45.451 159.844 45.515 ;
			RECT	160.148 45.451 160.18 45.515 ;
			RECT	160.484 45.451 160.516 45.515 ;
			RECT	160.82 45.451 160.852 45.515 ;
			RECT	161.156 45.451 161.188 45.515 ;
			RECT	161.492 45.451 161.524 45.515 ;
			RECT	161.828 45.451 161.86 45.515 ;
			RECT	162.154 45.451 162.186 45.515 ;
			RECT	162.5 45.451 162.532 45.515 ;
			RECT	162.836 45.451 162.868 45.515 ;
			RECT	163.172 45.451 163.204 45.515 ;
			RECT	163.508 45.451 163.54 45.515 ;
			RECT	163.844 45.451 163.876 45.515 ;
			RECT	164.18 45.451 164.212 45.515 ;
			RECT	164.516 45.451 164.548 45.515 ;
			RECT	164.852 45.451 164.884 45.515 ;
			RECT	165.188 45.451 165.22 45.515 ;
			RECT	165.524 45.451 165.556 45.515 ;
			RECT	165.86 45.451 165.892 45.515 ;
			RECT	166.196 45.451 166.228 45.515 ;
			RECT	166.532 45.451 166.564 45.515 ;
			RECT	166.868 45.451 166.9 45.515 ;
			RECT	167.204 45.451 167.236 45.515 ;
			RECT	167.54 45.451 167.572 45.515 ;
			RECT	167.876 45.451 167.908 45.515 ;
			RECT	168.212 45.451 168.244 45.515 ;
			RECT	168.548 45.451 168.58 45.515 ;
			RECT	168.884 45.451 168.916 45.515 ;
			RECT	169.22 45.451 169.252 45.515 ;
			RECT	169.556 45.451 169.588 45.515 ;
			RECT	169.892 45.451 169.924 45.515 ;
			RECT	170.228 45.451 170.26 45.515 ;
			RECT	170.564 45.451 170.596 45.515 ;
			RECT	170.9 45.451 170.932 45.515 ;
			RECT	171.236 45.451 171.268 45.515 ;
			RECT	171.572 45.451 171.604 45.515 ;
			RECT	171.908 45.451 171.94 45.515 ;
			RECT	172.244 45.451 172.276 45.515 ;
			RECT	172.58 45.451 172.612 45.515 ;
			RECT	172.916 45.451 172.948 45.515 ;
			RECT	173.252 45.451 173.284 45.515 ;
			RECT	173.588 45.451 173.62 45.515 ;
			RECT	173.924 45.451 173.956 45.515 ;
			RECT	174.26 45.451 174.292 45.515 ;
			RECT	174.596 45.451 174.628 45.515 ;
			RECT	174.932 45.451 174.964 45.515 ;
			RECT	175.268 45.451 175.3 45.515 ;
			RECT	175.604 45.451 175.636 45.515 ;
			RECT	175.94 45.451 175.972 45.515 ;
			RECT	176.276 45.451 176.308 45.515 ;
			RECT	176.612 45.451 176.644 45.515 ;
			RECT	176.948 45.451 176.98 45.515 ;
			RECT	177.284 45.451 177.316 45.515 ;
			RECT	177.62 45.451 177.652 45.515 ;
			RECT	177.956 45.451 177.988 45.515 ;
			RECT	178.292 45.451 178.324 45.515 ;
			RECT	178.623 45.451 178.655 45.515 ;
			RECT	178.959 45.451 178.991 45.515 ;
			RECT	179.295 45.451 179.327 45.515 ;
			RECT	179.631 45.451 179.663 45.515 ;
			RECT	179.967 45.451 179.999 45.515 ;
			RECT	180.303 45.451 180.335 45.515 ;
			RECT	180.639 45.451 180.671 45.515 ;
			RECT	180.975 45.451 181.007 45.515 ;
			RECT	181.311 45.451 181.343 45.515 ;
			RECT	181.647 45.451 181.679 45.515 ;
			RECT	181.983 45.451 182.015 45.515 ;
			RECT	182.319 45.451 182.351 45.515 ;
			RECT	182.655 45.451 182.687 45.515 ;
			RECT	182.991 45.451 183.023 45.515 ;
			RECT	183.327 45.451 183.359 45.515 ;
			RECT	183.663 45.451 183.695 45.515 ;
			RECT	183.999 45.451 184.031 45.515 ;
			RECT	184.335 45.451 184.367 45.515 ;
			RECT	184.671 45.451 184.703 45.515 ;
			RECT	185.007 45.451 185.039 45.515 ;
			RECT	185.343 45.451 185.375 45.515 ;
			RECT	185.679 45.451 185.711 45.515 ;
			RECT	186.015 45.451 186.047 45.515 ;
			RECT	186.351 45.451 186.383 45.515 ;
			RECT	186.687 45.451 186.719 45.515 ;
			RECT	187.023 45.451 187.055 45.515 ;
			RECT	187.359 45.451 187.391 45.515 ;
			RECT	187.695 45.451 187.727 45.515 ;
			RECT	188.031 45.451 188.063 45.515 ;
			RECT	188.367 45.451 188.399 45.515 ;
			RECT	188.703 45.451 188.735 45.515 ;
			RECT	189.039 45.451 189.071 45.515 ;
			RECT	189.375 45.451 189.407 45.515 ;
			RECT	189.711 45.451 189.743 45.515 ;
			RECT	190.047 45.451 190.079 45.515 ;
			RECT	190.383 45.451 190.415 45.515 ;
			RECT	190.719 45.451 190.751 45.515 ;
			RECT	191.055 45.451 191.087 45.515 ;
			RECT	191.391 45.451 191.423 45.515 ;
			RECT	191.727 45.451 191.759 45.515 ;
			RECT	192.063 45.451 192.095 45.515 ;
			RECT	192.399 45.451 192.431 45.515 ;
			RECT	192.735 45.451 192.767 45.515 ;
			RECT	193.071 45.451 193.103 45.515 ;
			RECT	193.407 45.451 193.439 45.515 ;
			RECT	193.743 45.451 193.775 45.515 ;
			RECT	194.079 45.451 194.111 45.515 ;
			RECT	194.415 45.451 194.447 45.515 ;
			RECT	194.751 45.451 194.783 45.515 ;
			RECT	195.087 45.451 195.119 45.515 ;
			RECT	195.423 45.451 195.455 45.515 ;
			RECT	195.759 45.451 195.791 45.515 ;
			RECT	196.095 45.451 196.127 45.515 ;
			RECT	196.431 45.451 196.463 45.515 ;
			RECT	196.767 45.451 196.799 45.515 ;
			RECT	197.103 45.451 197.135 45.515 ;
			RECT	197.439 45.451 197.471 45.515 ;
			RECT	197.775 45.451 197.807 45.515 ;
			RECT	198.111 45.451 198.143 45.515 ;
			RECT	198.447 45.451 198.479 45.515 ;
			RECT	198.783 45.451 198.815 45.515 ;
			RECT	199.119 45.451 199.151 45.515 ;
			RECT	199.455 45.451 199.487 45.515 ;
			RECT	199.791 45.451 199.823 45.515 ;
			RECT	201.14 45.451 201.204 45.515 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 46.918 201.665 47.038 ;
			LAYER	J3 ;
			RECT	5.514 46.946 5.578 47.01 ;
			RECT	6.379 46.946 6.411 47.01 ;
			RECT	6.715 46.946 6.747 47.01 ;
			RECT	7.051 46.946 7.083 47.01 ;
			RECT	7.387 46.946 7.419 47.01 ;
			RECT	7.723 46.946 7.755 47.01 ;
			RECT	8.059 46.946 8.091 47.01 ;
			RECT	8.395 46.946 8.427 47.01 ;
			RECT	8.731 46.946 8.763 47.01 ;
			RECT	9.067 46.946 9.099 47.01 ;
			RECT	9.403 46.946 9.435 47.01 ;
			RECT	9.739 46.946 9.771 47.01 ;
			RECT	10.075 46.946 10.107 47.01 ;
			RECT	10.411 46.946 10.443 47.01 ;
			RECT	10.747 46.946 10.779 47.01 ;
			RECT	11.083 46.946 11.115 47.01 ;
			RECT	11.419 46.946 11.451 47.01 ;
			RECT	11.755 46.946 11.787 47.01 ;
			RECT	12.091 46.946 12.123 47.01 ;
			RECT	12.427 46.946 12.459 47.01 ;
			RECT	12.763 46.946 12.795 47.01 ;
			RECT	13.099 46.946 13.131 47.01 ;
			RECT	13.435 46.946 13.467 47.01 ;
			RECT	13.771 46.946 13.803 47.01 ;
			RECT	14.107 46.946 14.139 47.01 ;
			RECT	14.443 46.946 14.475 47.01 ;
			RECT	14.779 46.946 14.811 47.01 ;
			RECT	15.115 46.946 15.147 47.01 ;
			RECT	15.451 46.946 15.483 47.01 ;
			RECT	15.787 46.946 15.819 47.01 ;
			RECT	16.123 46.946 16.155 47.01 ;
			RECT	16.459 46.946 16.491 47.01 ;
			RECT	16.795 46.946 16.827 47.01 ;
			RECT	17.131 46.946 17.163 47.01 ;
			RECT	17.467 46.946 17.499 47.01 ;
			RECT	17.803 46.946 17.835 47.01 ;
			RECT	18.139 46.946 18.171 47.01 ;
			RECT	18.475 46.946 18.507 47.01 ;
			RECT	18.811 46.946 18.843 47.01 ;
			RECT	19.147 46.946 19.179 47.01 ;
			RECT	19.483 46.946 19.515 47.01 ;
			RECT	19.819 46.946 19.851 47.01 ;
			RECT	20.155 46.946 20.187 47.01 ;
			RECT	20.491 46.946 20.523 47.01 ;
			RECT	20.827 46.946 20.859 47.01 ;
			RECT	21.163 46.946 21.195 47.01 ;
			RECT	21.499 46.946 21.531 47.01 ;
			RECT	21.835 46.946 21.867 47.01 ;
			RECT	22.171 46.946 22.203 47.01 ;
			RECT	22.507 46.946 22.539 47.01 ;
			RECT	22.843 46.946 22.875 47.01 ;
			RECT	23.179 46.946 23.211 47.01 ;
			RECT	23.515 46.946 23.547 47.01 ;
			RECT	23.851 46.946 23.883 47.01 ;
			RECT	24.187 46.946 24.219 47.01 ;
			RECT	24.523 46.946 24.555 47.01 ;
			RECT	24.859 46.946 24.891 47.01 ;
			RECT	25.195 46.946 25.227 47.01 ;
			RECT	25.531 46.946 25.563 47.01 ;
			RECT	25.867 46.946 25.899 47.01 ;
			RECT	26.203 46.946 26.235 47.01 ;
			RECT	26.539 46.946 26.571 47.01 ;
			RECT	26.875 46.946 26.907 47.01 ;
			RECT	27.211 46.946 27.243 47.01 ;
			RECT	27.547 46.946 27.579 47.01 ;
			RECT	27.878 46.946 27.91 47.01 ;
			RECT	28.214 46.946 28.246 47.01 ;
			RECT	28.55 46.946 28.582 47.01 ;
			RECT	28.886 46.946 28.918 47.01 ;
			RECT	29.222 46.946 29.254 47.01 ;
			RECT	29.558 46.946 29.59 47.01 ;
			RECT	29.894 46.946 29.926 47.01 ;
			RECT	30.23 46.946 30.262 47.01 ;
			RECT	30.566 46.946 30.598 47.01 ;
			RECT	30.902 46.946 30.934 47.01 ;
			RECT	31.238 46.946 31.27 47.01 ;
			RECT	31.574 46.946 31.606 47.01 ;
			RECT	31.91 46.946 31.942 47.01 ;
			RECT	32.246 46.946 32.278 47.01 ;
			RECT	32.582 46.946 32.614 47.01 ;
			RECT	32.918 46.946 32.95 47.01 ;
			RECT	33.254 46.946 33.286 47.01 ;
			RECT	33.59 46.946 33.622 47.01 ;
			RECT	33.926 46.946 33.958 47.01 ;
			RECT	34.262 46.946 34.294 47.01 ;
			RECT	34.598 46.946 34.63 47.01 ;
			RECT	34.934 46.946 34.966 47.01 ;
			RECT	35.27 46.946 35.302 47.01 ;
			RECT	35.606 46.946 35.638 47.01 ;
			RECT	35.942 46.946 35.974 47.01 ;
			RECT	36.278 46.946 36.31 47.01 ;
			RECT	36.614 46.946 36.646 47.01 ;
			RECT	36.95 46.946 36.982 47.01 ;
			RECT	37.286 46.946 37.318 47.01 ;
			RECT	37.622 46.946 37.654 47.01 ;
			RECT	37.958 46.946 37.99 47.01 ;
			RECT	38.294 46.946 38.326 47.01 ;
			RECT	38.63 46.946 38.662 47.01 ;
			RECT	38.966 46.946 38.998 47.01 ;
			RECT	39.302 46.946 39.334 47.01 ;
			RECT	39.638 46.946 39.67 47.01 ;
			RECT	39.974 46.946 40.006 47.01 ;
			RECT	40.31 46.946 40.342 47.01 ;
			RECT	40.646 46.946 40.678 47.01 ;
			RECT	40.982 46.946 41.014 47.01 ;
			RECT	41.318 46.946 41.35 47.01 ;
			RECT	41.654 46.946 41.686 47.01 ;
			RECT	41.99 46.946 42.022 47.01 ;
			RECT	42.326 46.946 42.358 47.01 ;
			RECT	42.662 46.946 42.694 47.01 ;
			RECT	42.998 46.946 43.03 47.01 ;
			RECT	43.334 46.946 43.366 47.01 ;
			RECT	43.67 46.946 43.702 47.01 ;
			RECT	44.342 46.946 44.374 47.01 ;
			RECT	44.678 46.946 44.71 47.01 ;
			RECT	45.014 46.946 45.046 47.01 ;
			RECT	45.35 46.946 45.382 47.01 ;
			RECT	45.686 46.946 45.718 47.01 ;
			RECT	46.022 46.946 46.054 47.01 ;
			RECT	46.358 46.946 46.39 47.01 ;
			RECT	46.694 46.946 46.726 47.01 ;
			RECT	47.03 46.946 47.062 47.01 ;
			RECT	47.366 46.946 47.398 47.01 ;
			RECT	47.702 46.946 47.734 47.01 ;
			RECT	48.038 46.946 48.07 47.01 ;
			RECT	48.374 46.946 48.406 47.01 ;
			RECT	48.71 46.946 48.742 47.01 ;
			RECT	49.046 46.946 49.078 47.01 ;
			RECT	49.457 46.946 49.489 47.01 ;
			RECT	50.433 46.946 50.465 47.01 ;
			RECT	51.274 46.946 51.306 47.01 ;
			RECT	51.794 46.946 51.826 47.01 ;
			RECT	54.657 46.946 54.689 47.01 ;
			RECT	56.144 46.946 56.176 47.01 ;
			RECT	56.664 46.946 56.696 47.01 ;
			RECT	57.507 46.946 57.571 47.01 ;
			RECT	58.715 46.946 58.747 47.01 ;
			RECT	59.126 46.946 59.158 47.01 ;
			RECT	59.462 46.946 59.494 47.01 ;
			RECT	59.798 46.946 59.83 47.01 ;
			RECT	60.134 46.946 60.166 47.01 ;
			RECT	60.47 46.946 60.502 47.01 ;
			RECT	60.806 46.946 60.838 47.01 ;
			RECT	61.142 46.946 61.174 47.01 ;
			RECT	61.478 46.946 61.51 47.01 ;
			RECT	61.814 46.946 61.846 47.01 ;
			RECT	62.15 46.946 62.182 47.01 ;
			RECT	62.486 46.946 62.518 47.01 ;
			RECT	62.822 46.946 62.854 47.01 ;
			RECT	63.158 46.946 63.19 47.01 ;
			RECT	63.494 46.946 63.526 47.01 ;
			RECT	63.83 46.946 63.862 47.01 ;
			RECT	64.502 46.946 64.534 47.01 ;
			RECT	64.838 46.946 64.87 47.01 ;
			RECT	65.174 46.946 65.206 47.01 ;
			RECT	65.51 46.946 65.542 47.01 ;
			RECT	65.846 46.946 65.878 47.01 ;
			RECT	66.182 46.946 66.214 47.01 ;
			RECT	66.518 46.946 66.55 47.01 ;
			RECT	66.854 46.946 66.886 47.01 ;
			RECT	67.19 46.946 67.222 47.01 ;
			RECT	67.526 46.946 67.558 47.01 ;
			RECT	67.862 46.946 67.894 47.01 ;
			RECT	68.198 46.946 68.23 47.01 ;
			RECT	68.534 46.946 68.566 47.01 ;
			RECT	68.87 46.946 68.902 47.01 ;
			RECT	69.206 46.946 69.238 47.01 ;
			RECT	69.542 46.946 69.574 47.01 ;
			RECT	69.878 46.946 69.91 47.01 ;
			RECT	70.214 46.946 70.246 47.01 ;
			RECT	70.55 46.946 70.582 47.01 ;
			RECT	70.886 46.946 70.918 47.01 ;
			RECT	71.222 46.946 71.254 47.01 ;
			RECT	71.558 46.946 71.59 47.01 ;
			RECT	71.894 46.946 71.926 47.01 ;
			RECT	72.23 46.946 72.262 47.01 ;
			RECT	72.566 46.946 72.598 47.01 ;
			RECT	72.902 46.946 72.934 47.01 ;
			RECT	73.238 46.946 73.27 47.01 ;
			RECT	73.574 46.946 73.606 47.01 ;
			RECT	73.91 46.946 73.942 47.01 ;
			RECT	74.246 46.946 74.278 47.01 ;
			RECT	74.582 46.946 74.614 47.01 ;
			RECT	74.918 46.946 74.95 47.01 ;
			RECT	75.254 46.946 75.286 47.01 ;
			RECT	75.59 46.946 75.622 47.01 ;
			RECT	75.926 46.946 75.958 47.01 ;
			RECT	76.262 46.946 76.294 47.01 ;
			RECT	76.598 46.946 76.63 47.01 ;
			RECT	76.934 46.946 76.966 47.01 ;
			RECT	77.27 46.946 77.302 47.01 ;
			RECT	77.606 46.946 77.638 47.01 ;
			RECT	77.942 46.946 77.974 47.01 ;
			RECT	78.278 46.946 78.31 47.01 ;
			RECT	78.614 46.946 78.646 47.01 ;
			RECT	78.95 46.946 78.982 47.01 ;
			RECT	79.286 46.946 79.318 47.01 ;
			RECT	79.622 46.946 79.654 47.01 ;
			RECT	79.958 46.946 79.99 47.01 ;
			RECT	80.294 46.946 80.326 47.01 ;
			RECT	80.625 46.946 80.657 47.01 ;
			RECT	80.961 46.946 80.993 47.01 ;
			RECT	81.297 46.946 81.329 47.01 ;
			RECT	81.633 46.946 81.665 47.01 ;
			RECT	81.969 46.946 82.001 47.01 ;
			RECT	82.305 46.946 82.337 47.01 ;
			RECT	82.641 46.946 82.673 47.01 ;
			RECT	82.977 46.946 83.009 47.01 ;
			RECT	83.313 46.946 83.345 47.01 ;
			RECT	83.649 46.946 83.681 47.01 ;
			RECT	83.985 46.946 84.017 47.01 ;
			RECT	84.321 46.946 84.353 47.01 ;
			RECT	84.657 46.946 84.689 47.01 ;
			RECT	84.993 46.946 85.025 47.01 ;
			RECT	85.329 46.946 85.361 47.01 ;
			RECT	85.665 46.946 85.697 47.01 ;
			RECT	86.001 46.946 86.033 47.01 ;
			RECT	86.337 46.946 86.369 47.01 ;
			RECT	86.673 46.946 86.705 47.01 ;
			RECT	87.009 46.946 87.041 47.01 ;
			RECT	87.345 46.946 87.377 47.01 ;
			RECT	87.681 46.946 87.713 47.01 ;
			RECT	88.017 46.946 88.049 47.01 ;
			RECT	88.353 46.946 88.385 47.01 ;
			RECT	88.689 46.946 88.721 47.01 ;
			RECT	89.025 46.946 89.057 47.01 ;
			RECT	89.361 46.946 89.393 47.01 ;
			RECT	89.697 46.946 89.729 47.01 ;
			RECT	90.033 46.946 90.065 47.01 ;
			RECT	90.369 46.946 90.401 47.01 ;
			RECT	90.705 46.946 90.737 47.01 ;
			RECT	91.041 46.946 91.073 47.01 ;
			RECT	91.377 46.946 91.409 47.01 ;
			RECT	91.713 46.946 91.745 47.01 ;
			RECT	92.049 46.946 92.081 47.01 ;
			RECT	92.385 46.946 92.417 47.01 ;
			RECT	92.721 46.946 92.753 47.01 ;
			RECT	93.057 46.946 93.089 47.01 ;
			RECT	93.393 46.946 93.425 47.01 ;
			RECT	93.729 46.946 93.761 47.01 ;
			RECT	94.065 46.946 94.097 47.01 ;
			RECT	94.401 46.946 94.433 47.01 ;
			RECT	94.737 46.946 94.769 47.01 ;
			RECT	95.073 46.946 95.105 47.01 ;
			RECT	95.409 46.946 95.441 47.01 ;
			RECT	95.745 46.946 95.777 47.01 ;
			RECT	96.081 46.946 96.113 47.01 ;
			RECT	96.417 46.946 96.449 47.01 ;
			RECT	96.753 46.946 96.785 47.01 ;
			RECT	97.089 46.946 97.121 47.01 ;
			RECT	97.425 46.946 97.457 47.01 ;
			RECT	97.761 46.946 97.793 47.01 ;
			RECT	98.097 46.946 98.129 47.01 ;
			RECT	98.433 46.946 98.465 47.01 ;
			RECT	98.769 46.946 98.801 47.01 ;
			RECT	99.105 46.946 99.137 47.01 ;
			RECT	99.441 46.946 99.473 47.01 ;
			RECT	99.777 46.946 99.809 47.01 ;
			RECT	100.113 46.946 100.145 47.01 ;
			RECT	100.449 46.946 100.481 47.01 ;
			RECT	100.785 46.946 100.817 47.01 ;
			RECT	101.121 46.946 101.153 47.01 ;
			RECT	101.457 46.946 101.489 47.01 ;
			RECT	101.793 46.946 101.825 47.01 ;
			RECT	102.626 46.946 102.69 47.01 ;
			RECT	103.512 46.946 103.576 47.01 ;
			RECT	104.377 46.946 104.409 47.01 ;
			RECT	104.713 46.946 104.745 47.01 ;
			RECT	105.049 46.946 105.081 47.01 ;
			RECT	105.385 46.946 105.417 47.01 ;
			RECT	105.721 46.946 105.753 47.01 ;
			RECT	106.057 46.946 106.089 47.01 ;
			RECT	106.393 46.946 106.425 47.01 ;
			RECT	106.729 46.946 106.761 47.01 ;
			RECT	107.065 46.946 107.097 47.01 ;
			RECT	107.401 46.946 107.433 47.01 ;
			RECT	107.737 46.946 107.769 47.01 ;
			RECT	108.073 46.946 108.105 47.01 ;
			RECT	108.409 46.946 108.441 47.01 ;
			RECT	108.745 46.946 108.777 47.01 ;
			RECT	109.081 46.946 109.113 47.01 ;
			RECT	109.417 46.946 109.449 47.01 ;
			RECT	109.753 46.946 109.785 47.01 ;
			RECT	110.089 46.946 110.121 47.01 ;
			RECT	110.425 46.946 110.457 47.01 ;
			RECT	110.761 46.946 110.793 47.01 ;
			RECT	111.097 46.946 111.129 47.01 ;
			RECT	111.433 46.946 111.465 47.01 ;
			RECT	111.769 46.946 111.801 47.01 ;
			RECT	112.105 46.946 112.137 47.01 ;
			RECT	112.441 46.946 112.473 47.01 ;
			RECT	112.777 46.946 112.809 47.01 ;
			RECT	113.113 46.946 113.145 47.01 ;
			RECT	113.449 46.946 113.481 47.01 ;
			RECT	113.785 46.946 113.817 47.01 ;
			RECT	114.121 46.946 114.153 47.01 ;
			RECT	114.457 46.946 114.489 47.01 ;
			RECT	114.793 46.946 114.825 47.01 ;
			RECT	115.129 46.946 115.161 47.01 ;
			RECT	115.465 46.946 115.497 47.01 ;
			RECT	115.801 46.946 115.833 47.01 ;
			RECT	116.137 46.946 116.169 47.01 ;
			RECT	116.473 46.946 116.505 47.01 ;
			RECT	116.809 46.946 116.841 47.01 ;
			RECT	117.145 46.946 117.177 47.01 ;
			RECT	117.481 46.946 117.513 47.01 ;
			RECT	117.817 46.946 117.849 47.01 ;
			RECT	118.153 46.946 118.185 47.01 ;
			RECT	118.489 46.946 118.521 47.01 ;
			RECT	118.825 46.946 118.857 47.01 ;
			RECT	119.161 46.946 119.193 47.01 ;
			RECT	119.497 46.946 119.529 47.01 ;
			RECT	119.833 46.946 119.865 47.01 ;
			RECT	120.169 46.946 120.201 47.01 ;
			RECT	120.505 46.946 120.537 47.01 ;
			RECT	120.841 46.946 120.873 47.01 ;
			RECT	121.177 46.946 121.209 47.01 ;
			RECT	121.513 46.946 121.545 47.01 ;
			RECT	121.849 46.946 121.881 47.01 ;
			RECT	122.185 46.946 122.217 47.01 ;
			RECT	122.521 46.946 122.553 47.01 ;
			RECT	122.857 46.946 122.889 47.01 ;
			RECT	123.193 46.946 123.225 47.01 ;
			RECT	123.529 46.946 123.561 47.01 ;
			RECT	123.865 46.946 123.897 47.01 ;
			RECT	124.201 46.946 124.233 47.01 ;
			RECT	124.537 46.946 124.569 47.01 ;
			RECT	124.873 46.946 124.905 47.01 ;
			RECT	125.209 46.946 125.241 47.01 ;
			RECT	125.545 46.946 125.577 47.01 ;
			RECT	125.876 46.946 125.908 47.01 ;
			RECT	126.212 46.946 126.244 47.01 ;
			RECT	126.548 46.946 126.58 47.01 ;
			RECT	126.884 46.946 126.916 47.01 ;
			RECT	127.22 46.946 127.252 47.01 ;
			RECT	127.556 46.946 127.588 47.01 ;
			RECT	127.892 46.946 127.924 47.01 ;
			RECT	128.228 46.946 128.26 47.01 ;
			RECT	128.564 46.946 128.596 47.01 ;
			RECT	128.9 46.946 128.932 47.01 ;
			RECT	129.236 46.946 129.268 47.01 ;
			RECT	129.572 46.946 129.604 47.01 ;
			RECT	129.908 46.946 129.94 47.01 ;
			RECT	130.244 46.946 130.276 47.01 ;
			RECT	130.58 46.946 130.612 47.01 ;
			RECT	130.916 46.946 130.948 47.01 ;
			RECT	131.252 46.946 131.284 47.01 ;
			RECT	131.588 46.946 131.62 47.01 ;
			RECT	131.924 46.946 131.956 47.01 ;
			RECT	132.26 46.946 132.292 47.01 ;
			RECT	132.596 46.946 132.628 47.01 ;
			RECT	132.932 46.946 132.964 47.01 ;
			RECT	133.268 46.946 133.3 47.01 ;
			RECT	133.604 46.946 133.636 47.01 ;
			RECT	133.94 46.946 133.972 47.01 ;
			RECT	134.276 46.946 134.308 47.01 ;
			RECT	134.612 46.946 134.644 47.01 ;
			RECT	134.948 46.946 134.98 47.01 ;
			RECT	135.284 46.946 135.316 47.01 ;
			RECT	135.62 46.946 135.652 47.01 ;
			RECT	135.956 46.946 135.988 47.01 ;
			RECT	136.292 46.946 136.324 47.01 ;
			RECT	136.628 46.946 136.66 47.01 ;
			RECT	136.964 46.946 136.996 47.01 ;
			RECT	137.3 46.946 137.332 47.01 ;
			RECT	137.636 46.946 137.668 47.01 ;
			RECT	137.972 46.946 138.004 47.01 ;
			RECT	138.308 46.946 138.34 47.01 ;
			RECT	138.644 46.946 138.676 47.01 ;
			RECT	138.98 46.946 139.012 47.01 ;
			RECT	139.316 46.946 139.348 47.01 ;
			RECT	139.652 46.946 139.684 47.01 ;
			RECT	139.988 46.946 140.02 47.01 ;
			RECT	140.324 46.946 140.356 47.01 ;
			RECT	140.66 46.946 140.692 47.01 ;
			RECT	140.996 46.946 141.028 47.01 ;
			RECT	141.332 46.946 141.364 47.01 ;
			RECT	141.668 46.946 141.7 47.01 ;
			RECT	142.34 46.946 142.372 47.01 ;
			RECT	142.676 46.946 142.708 47.01 ;
			RECT	143.012 46.946 143.044 47.01 ;
			RECT	143.348 46.946 143.38 47.01 ;
			RECT	143.684 46.946 143.716 47.01 ;
			RECT	144.02 46.946 144.052 47.01 ;
			RECT	144.356 46.946 144.388 47.01 ;
			RECT	144.692 46.946 144.724 47.01 ;
			RECT	145.028 46.946 145.06 47.01 ;
			RECT	145.364 46.946 145.396 47.01 ;
			RECT	145.7 46.946 145.732 47.01 ;
			RECT	146.036 46.946 146.068 47.01 ;
			RECT	146.372 46.946 146.404 47.01 ;
			RECT	146.708 46.946 146.74 47.01 ;
			RECT	147.044 46.946 147.076 47.01 ;
			RECT	147.455 46.946 147.487 47.01 ;
			RECT	148.431 46.946 148.463 47.01 ;
			RECT	149.272 46.946 149.304 47.01 ;
			RECT	149.792 46.946 149.824 47.01 ;
			RECT	152.655 46.946 152.687 47.01 ;
			RECT	154.142 46.946 154.174 47.01 ;
			RECT	154.662 46.946 154.694 47.01 ;
			RECT	155.505 46.946 155.569 47.01 ;
			RECT	156.713 46.946 156.745 47.01 ;
			RECT	157.124 46.946 157.156 47.01 ;
			RECT	157.46 46.946 157.492 47.01 ;
			RECT	157.796 46.946 157.828 47.01 ;
			RECT	158.132 46.946 158.164 47.01 ;
			RECT	158.468 46.946 158.5 47.01 ;
			RECT	158.804 46.946 158.836 47.01 ;
			RECT	159.14 46.946 159.172 47.01 ;
			RECT	159.476 46.946 159.508 47.01 ;
			RECT	159.812 46.946 159.844 47.01 ;
			RECT	160.148 46.946 160.18 47.01 ;
			RECT	160.484 46.946 160.516 47.01 ;
			RECT	160.82 46.946 160.852 47.01 ;
			RECT	161.156 46.946 161.188 47.01 ;
			RECT	161.492 46.946 161.524 47.01 ;
			RECT	161.828 46.946 161.86 47.01 ;
			RECT	162.5 46.946 162.532 47.01 ;
			RECT	162.836 46.946 162.868 47.01 ;
			RECT	163.172 46.946 163.204 47.01 ;
			RECT	163.508 46.946 163.54 47.01 ;
			RECT	163.844 46.946 163.876 47.01 ;
			RECT	164.18 46.946 164.212 47.01 ;
			RECT	164.516 46.946 164.548 47.01 ;
			RECT	164.852 46.946 164.884 47.01 ;
			RECT	165.188 46.946 165.22 47.01 ;
			RECT	165.524 46.946 165.556 47.01 ;
			RECT	165.86 46.946 165.892 47.01 ;
			RECT	166.196 46.946 166.228 47.01 ;
			RECT	166.532 46.946 166.564 47.01 ;
			RECT	166.868 46.946 166.9 47.01 ;
			RECT	167.204 46.946 167.236 47.01 ;
			RECT	167.54 46.946 167.572 47.01 ;
			RECT	167.876 46.946 167.908 47.01 ;
			RECT	168.212 46.946 168.244 47.01 ;
			RECT	168.548 46.946 168.58 47.01 ;
			RECT	168.884 46.946 168.916 47.01 ;
			RECT	169.22 46.946 169.252 47.01 ;
			RECT	169.556 46.946 169.588 47.01 ;
			RECT	169.892 46.946 169.924 47.01 ;
			RECT	170.228 46.946 170.26 47.01 ;
			RECT	170.564 46.946 170.596 47.01 ;
			RECT	170.9 46.946 170.932 47.01 ;
			RECT	171.236 46.946 171.268 47.01 ;
			RECT	171.572 46.946 171.604 47.01 ;
			RECT	171.908 46.946 171.94 47.01 ;
			RECT	172.244 46.946 172.276 47.01 ;
			RECT	172.58 46.946 172.612 47.01 ;
			RECT	172.916 46.946 172.948 47.01 ;
			RECT	173.252 46.946 173.284 47.01 ;
			RECT	173.588 46.946 173.62 47.01 ;
			RECT	173.924 46.946 173.956 47.01 ;
			RECT	174.26 46.946 174.292 47.01 ;
			RECT	174.596 46.946 174.628 47.01 ;
			RECT	174.932 46.946 174.964 47.01 ;
			RECT	175.268 46.946 175.3 47.01 ;
			RECT	175.604 46.946 175.636 47.01 ;
			RECT	175.94 46.946 175.972 47.01 ;
			RECT	176.276 46.946 176.308 47.01 ;
			RECT	176.612 46.946 176.644 47.01 ;
			RECT	176.948 46.946 176.98 47.01 ;
			RECT	177.284 46.946 177.316 47.01 ;
			RECT	177.62 46.946 177.652 47.01 ;
			RECT	177.956 46.946 177.988 47.01 ;
			RECT	178.292 46.946 178.324 47.01 ;
			RECT	178.623 46.946 178.655 47.01 ;
			RECT	178.959 46.946 178.991 47.01 ;
			RECT	179.295 46.946 179.327 47.01 ;
			RECT	179.631 46.946 179.663 47.01 ;
			RECT	179.967 46.946 179.999 47.01 ;
			RECT	180.303 46.946 180.335 47.01 ;
			RECT	180.639 46.946 180.671 47.01 ;
			RECT	180.975 46.946 181.007 47.01 ;
			RECT	181.311 46.946 181.343 47.01 ;
			RECT	181.647 46.946 181.679 47.01 ;
			RECT	181.983 46.946 182.015 47.01 ;
			RECT	182.319 46.946 182.351 47.01 ;
			RECT	182.655 46.946 182.687 47.01 ;
			RECT	182.991 46.946 183.023 47.01 ;
			RECT	183.327 46.946 183.359 47.01 ;
			RECT	183.663 46.946 183.695 47.01 ;
			RECT	183.999 46.946 184.031 47.01 ;
			RECT	184.335 46.946 184.367 47.01 ;
			RECT	184.671 46.946 184.703 47.01 ;
			RECT	185.007 46.946 185.039 47.01 ;
			RECT	185.343 46.946 185.375 47.01 ;
			RECT	185.679 46.946 185.711 47.01 ;
			RECT	186.015 46.946 186.047 47.01 ;
			RECT	186.351 46.946 186.383 47.01 ;
			RECT	186.687 46.946 186.719 47.01 ;
			RECT	187.023 46.946 187.055 47.01 ;
			RECT	187.359 46.946 187.391 47.01 ;
			RECT	187.695 46.946 187.727 47.01 ;
			RECT	188.031 46.946 188.063 47.01 ;
			RECT	188.367 46.946 188.399 47.01 ;
			RECT	188.703 46.946 188.735 47.01 ;
			RECT	189.039 46.946 189.071 47.01 ;
			RECT	189.375 46.946 189.407 47.01 ;
			RECT	189.711 46.946 189.743 47.01 ;
			RECT	190.047 46.946 190.079 47.01 ;
			RECT	190.383 46.946 190.415 47.01 ;
			RECT	190.719 46.946 190.751 47.01 ;
			RECT	191.055 46.946 191.087 47.01 ;
			RECT	191.391 46.946 191.423 47.01 ;
			RECT	191.727 46.946 191.759 47.01 ;
			RECT	192.063 46.946 192.095 47.01 ;
			RECT	192.399 46.946 192.431 47.01 ;
			RECT	192.735 46.946 192.767 47.01 ;
			RECT	193.071 46.946 193.103 47.01 ;
			RECT	193.407 46.946 193.439 47.01 ;
			RECT	193.743 46.946 193.775 47.01 ;
			RECT	194.079 46.946 194.111 47.01 ;
			RECT	194.415 46.946 194.447 47.01 ;
			RECT	194.751 46.946 194.783 47.01 ;
			RECT	195.087 46.946 195.119 47.01 ;
			RECT	195.423 46.946 195.455 47.01 ;
			RECT	195.759 46.946 195.791 47.01 ;
			RECT	196.095 46.946 196.127 47.01 ;
			RECT	196.431 46.946 196.463 47.01 ;
			RECT	196.767 46.946 196.799 47.01 ;
			RECT	197.103 46.946 197.135 47.01 ;
			RECT	197.439 46.946 197.471 47.01 ;
			RECT	197.775 46.946 197.807 47.01 ;
			RECT	198.111 46.946 198.143 47.01 ;
			RECT	198.447 46.946 198.479 47.01 ;
			RECT	198.783 46.946 198.815 47.01 ;
			RECT	199.119 46.946 199.151 47.01 ;
			RECT	199.455 46.946 199.487 47.01 ;
			RECT	199.791 46.946 199.823 47.01 ;
			RECT	200.624 46.946 200.688 47.01 ;
			RECT	201.14 46.946 201.204 47.01 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 48.443 201.665 48.563 ;
			LAYER	J3 ;
			RECT	5.514 48.471 5.578 48.535 ;
			RECT	49.457 48.471 49.489 48.535 ;
			RECT	49.691 48.471 49.723 48.535 ;
			RECT	50.433 48.471 50.465 48.535 ;
			RECT	51.274 48.471 51.306 48.535 ;
			RECT	51.794 48.471 51.826 48.535 ;
			RECT	54.657 48.471 54.689 48.535 ;
			RECT	56.144 48.471 56.176 48.535 ;
			RECT	56.664 48.471 56.696 48.535 ;
			RECT	57.507 48.471 57.571 48.535 ;
			RECT	58.481 48.471 58.513 48.535 ;
			RECT	58.715 48.471 58.747 48.535 ;
			RECT	102.626 48.471 102.69 48.535 ;
			RECT	103.512 48.471 103.576 48.535 ;
			RECT	147.455 48.471 147.487 48.535 ;
			RECT	147.689 48.471 147.721 48.535 ;
			RECT	148.431 48.471 148.463 48.535 ;
			RECT	149.272 48.471 149.304 48.535 ;
			RECT	149.792 48.471 149.824 48.535 ;
			RECT	152.655 48.471 152.687 48.535 ;
			RECT	154.142 48.471 154.174 48.535 ;
			RECT	154.662 48.471 154.694 48.535 ;
			RECT	155.505 48.471 155.569 48.535 ;
			RECT	156.479 48.471 156.511 48.535 ;
			RECT	156.713 48.471 156.745 48.535 ;
			RECT	200.624 48.471 200.688 48.535 ;
			RECT	201.14 48.471 201.204 48.535 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 49.598 201.665 49.708 ;
			LAYER	J3 ;
			RECT	5.514 49.621 5.578 49.685 ;
			RECT	102.626 49.621 102.69 49.685 ;
			RECT	103.512 49.621 103.576 49.685 ;
			RECT	200.624 49.621 200.688 49.685 ;
			RECT	201.156 49.621 201.188 49.685 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 33.063 201.665 33.153 ;
			LAYER	J3 ;
			RECT	5.675 33.076 5.707 33.14 ;
			RECT	49.691 33.076 49.723 33.14 ;
			RECT	54.676 33.095 54.708 33.127 ;
			RECT	58.481 33.076 58.513 33.14 ;
			RECT	102.497 33.076 102.529 33.14 ;
			RECT	103.673 33.076 103.705 33.14 ;
			RECT	147.689 33.076 147.721 33.14 ;
			RECT	152.674 33.095 152.706 33.127 ;
			RECT	156.479 33.076 156.511 33.14 ;
			RECT	200.495 33.076 200.527 33.14 ;
			RECT	201.14 33.092 201.204 33.124 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 49.023 201.665 49.113 ;
			LAYER	J3 ;
			RECT	5.675 49.036 5.707 49.1 ;
			RECT	49.691 49.036 49.723 49.1 ;
			RECT	54.657 49.052 54.689 49.084 ;
			RECT	58.481 49.036 58.513 49.1 ;
			RECT	102.497 49.036 102.529 49.1 ;
			RECT	103.673 49.036 103.705 49.1 ;
			RECT	147.689 49.036 147.721 49.1 ;
			RECT	152.655 49.052 152.687 49.084 ;
			RECT	156.479 49.036 156.511 49.1 ;
			RECT	200.495 49.036 200.527 49.1 ;
			RECT	201.14 49.052 201.204 49.084 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 81.678 201.665 81.768 ;
			LAYER	J3 ;
			RECT	1.067 81.691 1.099 81.755 ;
			RECT	1.223 81.691 1.255 81.755 ;
			RECT	5.675 81.691 5.707 81.755 ;
			RECT	49.691 81.691 49.723 81.755 ;
			RECT	58.481 81.691 58.513 81.755 ;
			RECT	102.497 81.691 102.529 81.755 ;
			RECT	103.673 81.691 103.705 81.755 ;
			RECT	147.689 81.691 147.721 81.755 ;
			RECT	156.479 81.691 156.511 81.755 ;
			RECT	200.495 81.691 200.527 81.755 ;
			RECT	201.14 81.707 201.204 81.739 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 0.408 201.665 0.498 ;
			LAYER	J3 ;
			RECT	1.067 0.421 1.099 0.485 ;
			RECT	1.223 0.421 1.255 0.485 ;
			RECT	5.675 0.421 5.707 0.485 ;
			RECT	49.691 0.421 49.723 0.485 ;
			RECT	58.481 0.421 58.513 0.485 ;
			RECT	102.497 0.421 102.529 0.485 ;
			RECT	103.673 0.421 103.705 0.485 ;
			RECT	147.689 0.421 147.721 0.485 ;
			RECT	156.479 0.421 156.511 0.485 ;
			RECT	200.495 0.421 200.527 0.485 ;
			RECT	201.14 0.437 201.204 0.469 ;
		END

	END VDDCE

	PIN VDDPE
		USE POWER ;
		DIRECTION INOUT ;
		PORT
			LAYER	C4 ;
			RECT	0.294 81.251 201.665 81.361 ;
			LAYER	J3 ;
			RECT	1.822 81.29 1.886 81.322 ;
			RECT	5.164 81.274 5.196 81.338 ;
			RECT	50.379 81.29 50.443 81.322 ;
			RECT	51.274 81.274 51.306 81.338 ;
			RECT	51.794 81.29 51.826 81.322 ;
			RECT	53.707 81.29 53.739 81.322 ;
			RECT	54.676 81.274 54.708 81.338 ;
			RECT	55.232 81.29 55.264 81.322 ;
			RECT	56.136 81.274 56.168 81.338 ;
			RECT	56.668 81.274 56.7 81.338 ;
			RECT	57.531 81.29 57.595 81.322 ;
			RECT	148.377 81.29 148.441 81.322 ;
			RECT	149.272 81.274 149.304 81.338 ;
			RECT	149.792 81.29 149.824 81.322 ;
			RECT	151.705 81.29 151.737 81.322 ;
			RECT	152.674 81.274 152.706 81.338 ;
			RECT	153.23 81.29 153.262 81.322 ;
			RECT	154.134 81.274 154.166 81.338 ;
			RECT	154.666 81.274 154.698 81.338 ;
			RECT	155.529 81.29 155.593 81.322 ;
			RECT	201.004 81.274 201.036 81.338 ;
			RECT	201.306 81.274 201.338 81.338 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 77.411 201.665 77.521 ;
			LAYER	J3 ;
			RECT	1.822 77.45 1.886 77.482 ;
			RECT	5.164 77.434 5.196 77.498 ;
			RECT	50.379 77.45 50.443 77.482 ;
			RECT	51.274 77.434 51.306 77.498 ;
			RECT	51.794 77.45 51.826 77.482 ;
			RECT	53.707 77.45 53.739 77.482 ;
			RECT	54.676 77.434 54.708 77.498 ;
			RECT	55.232 77.45 55.264 77.482 ;
			RECT	56.136 77.434 56.168 77.498 ;
			RECT	56.668 77.434 56.7 77.498 ;
			RECT	57.531 77.45 57.595 77.482 ;
			RECT	148.377 77.45 148.441 77.482 ;
			RECT	149.272 77.434 149.304 77.498 ;
			RECT	149.792 77.45 149.824 77.482 ;
			RECT	151.705 77.45 151.737 77.482 ;
			RECT	152.674 77.434 152.706 77.498 ;
			RECT	153.23 77.45 153.262 77.482 ;
			RECT	154.134 77.434 154.166 77.498 ;
			RECT	154.666 77.434 154.698 77.498 ;
			RECT	155.529 77.45 155.593 77.482 ;
			RECT	201.004 77.434 201.036 77.498 ;
			RECT	201.306 77.434 201.338 77.498 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 29.615 201.665 29.725 ;
			LAYER	J3 ;
			RECT	1.822 29.654 1.886 29.686 ;
			RECT	5.164 29.638 5.196 29.702 ;
			RECT	50.379 29.654 50.443 29.686 ;
			RECT	51.274 29.638 51.306 29.702 ;
			RECT	51.794 29.654 51.826 29.686 ;
			RECT	53.707 29.654 53.739 29.686 ;
			RECT	54.676 29.638 54.708 29.702 ;
			RECT	55.232 29.654 55.264 29.686 ;
			RECT	56.136 29.638 56.168 29.702 ;
			RECT	56.668 29.638 56.7 29.702 ;
			RECT	57.531 29.654 57.595 29.686 ;
			RECT	148.377 29.654 148.441 29.686 ;
			RECT	149.272 29.638 149.304 29.702 ;
			RECT	149.792 29.654 149.824 29.686 ;
			RECT	151.705 29.654 151.737 29.686 ;
			RECT	152.674 29.638 152.706 29.702 ;
			RECT	153.23 29.654 153.262 29.686 ;
			RECT	154.134 29.638 154.166 29.702 ;
			RECT	154.666 29.638 154.698 29.702 ;
			RECT	155.529 29.654 155.593 29.686 ;
			RECT	201.004 29.638 201.036 29.702 ;
			RECT	201.306 29.638 201.338 29.702 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 27.695 201.665 27.805 ;
			LAYER	J3 ;
			RECT	1.822 27.734 1.886 27.766 ;
			RECT	5.164 27.718 5.196 27.782 ;
			RECT	50.379 27.734 50.443 27.766 ;
			RECT	51.274 27.718 51.306 27.782 ;
			RECT	51.794 27.734 51.826 27.766 ;
			RECT	53.707 27.734 53.739 27.766 ;
			RECT	54.676 27.718 54.708 27.782 ;
			RECT	55.232 27.734 55.264 27.766 ;
			RECT	56.136 27.718 56.168 27.782 ;
			RECT	56.668 27.718 56.7 27.782 ;
			RECT	57.531 27.734 57.595 27.766 ;
			RECT	148.377 27.734 148.441 27.766 ;
			RECT	149.272 27.718 149.304 27.782 ;
			RECT	149.792 27.734 149.824 27.766 ;
			RECT	151.705 27.734 151.737 27.766 ;
			RECT	152.674 27.718 152.706 27.782 ;
			RECT	153.23 27.734 153.262 27.766 ;
			RECT	154.134 27.718 154.166 27.782 ;
			RECT	154.666 27.718 154.698 27.782 ;
			RECT	155.529 27.734 155.593 27.766 ;
			RECT	201.004 27.718 201.036 27.782 ;
			RECT	201.306 27.718 201.338 27.782 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 25.775 201.665 25.885 ;
			LAYER	J3 ;
			RECT	1.822 25.814 1.886 25.846 ;
			RECT	5.164 25.798 5.196 25.862 ;
			RECT	50.379 25.814 50.443 25.846 ;
			RECT	51.274 25.798 51.306 25.862 ;
			RECT	51.794 25.814 51.826 25.846 ;
			RECT	53.707 25.814 53.739 25.846 ;
			RECT	54.676 25.798 54.708 25.862 ;
			RECT	55.232 25.814 55.264 25.846 ;
			RECT	56.136 25.798 56.168 25.862 ;
			RECT	56.668 25.798 56.7 25.862 ;
			RECT	57.531 25.814 57.595 25.846 ;
			RECT	148.377 25.814 148.441 25.846 ;
			RECT	149.272 25.798 149.304 25.862 ;
			RECT	149.792 25.814 149.824 25.846 ;
			RECT	151.705 25.814 151.737 25.846 ;
			RECT	152.674 25.798 152.706 25.862 ;
			RECT	153.23 25.814 153.262 25.846 ;
			RECT	154.134 25.798 154.166 25.862 ;
			RECT	154.666 25.798 154.698 25.862 ;
			RECT	155.529 25.814 155.593 25.846 ;
			RECT	201.004 25.798 201.036 25.862 ;
			RECT	201.306 25.798 201.338 25.862 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 23.855 201.665 23.965 ;
			LAYER	J3 ;
			RECT	1.822 23.894 1.886 23.926 ;
			RECT	5.164 23.878 5.196 23.942 ;
			RECT	50.379 23.894 50.443 23.926 ;
			RECT	51.274 23.878 51.306 23.942 ;
			RECT	51.794 23.894 51.826 23.926 ;
			RECT	53.707 23.894 53.739 23.926 ;
			RECT	54.676 23.878 54.708 23.942 ;
			RECT	55.232 23.894 55.264 23.926 ;
			RECT	56.136 23.878 56.168 23.942 ;
			RECT	56.668 23.878 56.7 23.942 ;
			RECT	57.531 23.894 57.595 23.926 ;
			RECT	148.377 23.894 148.441 23.926 ;
			RECT	149.272 23.878 149.304 23.942 ;
			RECT	149.792 23.894 149.824 23.926 ;
			RECT	151.705 23.894 151.737 23.926 ;
			RECT	152.674 23.878 152.706 23.942 ;
			RECT	153.23 23.894 153.262 23.926 ;
			RECT	154.134 23.878 154.166 23.942 ;
			RECT	154.666 23.878 154.698 23.942 ;
			RECT	155.529 23.894 155.593 23.926 ;
			RECT	201.004 23.878 201.036 23.942 ;
			RECT	201.306 23.878 201.338 23.942 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 21.935 201.665 22.045 ;
			LAYER	J3 ;
			RECT	1.822 21.974 1.886 22.006 ;
			RECT	5.164 21.958 5.196 22.022 ;
			RECT	50.379 21.974 50.443 22.006 ;
			RECT	51.274 21.958 51.306 22.022 ;
			RECT	51.794 21.974 51.826 22.006 ;
			RECT	53.707 21.974 53.739 22.006 ;
			RECT	54.676 21.958 54.708 22.022 ;
			RECT	55.232 21.974 55.264 22.006 ;
			RECT	56.136 21.958 56.168 22.022 ;
			RECT	56.668 21.958 56.7 22.022 ;
			RECT	57.531 21.974 57.595 22.006 ;
			RECT	148.377 21.974 148.441 22.006 ;
			RECT	149.272 21.958 149.304 22.022 ;
			RECT	149.792 21.974 149.824 22.006 ;
			RECT	151.705 21.974 151.737 22.006 ;
			RECT	152.674 21.958 152.706 22.022 ;
			RECT	153.23 21.974 153.262 22.006 ;
			RECT	154.134 21.958 154.166 22.022 ;
			RECT	154.666 21.958 154.698 22.022 ;
			RECT	155.529 21.974 155.593 22.006 ;
			RECT	201.004 21.958 201.036 22.022 ;
			RECT	201.306 21.958 201.338 22.022 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 20.015 201.665 20.125 ;
			LAYER	J3 ;
			RECT	1.822 20.054 1.886 20.086 ;
			RECT	5.164 20.038 5.196 20.102 ;
			RECT	50.379 20.054 50.443 20.086 ;
			RECT	51.274 20.038 51.306 20.102 ;
			RECT	51.794 20.054 51.826 20.086 ;
			RECT	53.707 20.054 53.739 20.086 ;
			RECT	54.676 20.038 54.708 20.102 ;
			RECT	55.232 20.054 55.264 20.086 ;
			RECT	56.136 20.038 56.168 20.102 ;
			RECT	56.668 20.038 56.7 20.102 ;
			RECT	57.531 20.054 57.595 20.086 ;
			RECT	148.377 20.054 148.441 20.086 ;
			RECT	149.272 20.038 149.304 20.102 ;
			RECT	149.792 20.054 149.824 20.086 ;
			RECT	151.705 20.054 151.737 20.086 ;
			RECT	152.674 20.038 152.706 20.102 ;
			RECT	153.23 20.054 153.262 20.086 ;
			RECT	154.134 20.038 154.166 20.102 ;
			RECT	154.666 20.038 154.698 20.102 ;
			RECT	155.529 20.054 155.593 20.086 ;
			RECT	201.004 20.038 201.036 20.102 ;
			RECT	201.306 20.038 201.338 20.102 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 18.095 201.665 18.205 ;
			LAYER	J3 ;
			RECT	1.822 18.134 1.886 18.166 ;
			RECT	5.164 18.118 5.196 18.182 ;
			RECT	50.379 18.134 50.443 18.166 ;
			RECT	51.274 18.118 51.306 18.182 ;
			RECT	51.794 18.134 51.826 18.166 ;
			RECT	53.707 18.134 53.739 18.166 ;
			RECT	54.676 18.118 54.708 18.182 ;
			RECT	55.232 18.134 55.264 18.166 ;
			RECT	56.136 18.118 56.168 18.182 ;
			RECT	56.668 18.118 56.7 18.182 ;
			RECT	57.531 18.134 57.595 18.166 ;
			RECT	148.377 18.134 148.441 18.166 ;
			RECT	149.272 18.118 149.304 18.182 ;
			RECT	149.792 18.134 149.824 18.166 ;
			RECT	151.705 18.134 151.737 18.166 ;
			RECT	152.674 18.118 152.706 18.182 ;
			RECT	153.23 18.134 153.262 18.166 ;
			RECT	154.134 18.118 154.166 18.182 ;
			RECT	154.666 18.118 154.698 18.182 ;
			RECT	155.529 18.134 155.593 18.166 ;
			RECT	201.004 18.118 201.036 18.182 ;
			RECT	201.306 18.118 201.338 18.182 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 75.491 201.665 75.601 ;
			LAYER	J3 ;
			RECT	1.822 75.53 1.886 75.562 ;
			RECT	5.164 75.514 5.196 75.578 ;
			RECT	50.379 75.53 50.443 75.562 ;
			RECT	51.274 75.514 51.306 75.578 ;
			RECT	51.794 75.53 51.826 75.562 ;
			RECT	53.707 75.53 53.739 75.562 ;
			RECT	54.676 75.514 54.708 75.578 ;
			RECT	55.232 75.53 55.264 75.562 ;
			RECT	56.136 75.514 56.168 75.578 ;
			RECT	56.668 75.514 56.7 75.578 ;
			RECT	57.531 75.53 57.595 75.562 ;
			RECT	148.377 75.53 148.441 75.562 ;
			RECT	149.272 75.514 149.304 75.578 ;
			RECT	149.792 75.53 149.824 75.562 ;
			RECT	151.705 75.53 151.737 75.562 ;
			RECT	152.674 75.514 152.706 75.578 ;
			RECT	153.23 75.53 153.262 75.562 ;
			RECT	154.134 75.514 154.166 75.578 ;
			RECT	154.666 75.514 154.698 75.578 ;
			RECT	155.529 75.53 155.593 75.562 ;
			RECT	201.004 75.514 201.036 75.578 ;
			RECT	201.306 75.514 201.338 75.578 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 16.175 201.665 16.285 ;
			LAYER	J3 ;
			RECT	1.822 16.214 1.886 16.246 ;
			RECT	5.164 16.198 5.196 16.262 ;
			RECT	50.379 16.214 50.443 16.246 ;
			RECT	51.274 16.198 51.306 16.262 ;
			RECT	51.794 16.214 51.826 16.246 ;
			RECT	53.707 16.214 53.739 16.246 ;
			RECT	54.676 16.198 54.708 16.262 ;
			RECT	55.232 16.214 55.264 16.246 ;
			RECT	56.136 16.198 56.168 16.262 ;
			RECT	56.668 16.198 56.7 16.262 ;
			RECT	57.531 16.214 57.595 16.246 ;
			RECT	148.377 16.214 148.441 16.246 ;
			RECT	149.272 16.198 149.304 16.262 ;
			RECT	149.792 16.214 149.824 16.246 ;
			RECT	151.705 16.214 151.737 16.246 ;
			RECT	152.674 16.198 152.706 16.262 ;
			RECT	153.23 16.214 153.262 16.246 ;
			RECT	154.134 16.198 154.166 16.262 ;
			RECT	154.666 16.198 154.698 16.262 ;
			RECT	155.529 16.214 155.593 16.246 ;
			RECT	201.004 16.198 201.036 16.262 ;
			RECT	201.306 16.198 201.338 16.262 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 14.255 201.665 14.365 ;
			LAYER	J3 ;
			RECT	1.822 14.294 1.886 14.326 ;
			RECT	5.164 14.278 5.196 14.342 ;
			RECT	50.379 14.294 50.443 14.326 ;
			RECT	51.274 14.278 51.306 14.342 ;
			RECT	51.794 14.294 51.826 14.326 ;
			RECT	53.707 14.294 53.739 14.326 ;
			RECT	54.676 14.278 54.708 14.342 ;
			RECT	55.232 14.294 55.264 14.326 ;
			RECT	56.136 14.278 56.168 14.342 ;
			RECT	56.668 14.278 56.7 14.342 ;
			RECT	57.531 14.294 57.595 14.326 ;
			RECT	148.377 14.294 148.441 14.326 ;
			RECT	149.272 14.278 149.304 14.342 ;
			RECT	149.792 14.294 149.824 14.326 ;
			RECT	151.705 14.294 151.737 14.326 ;
			RECT	152.674 14.278 152.706 14.342 ;
			RECT	153.23 14.294 153.262 14.326 ;
			RECT	154.134 14.278 154.166 14.342 ;
			RECT	154.666 14.278 154.698 14.342 ;
			RECT	155.529 14.294 155.593 14.326 ;
			RECT	201.004 14.278 201.036 14.342 ;
			RECT	201.306 14.278 201.338 14.342 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 12.335 201.665 12.445 ;
			LAYER	J3 ;
			RECT	1.822 12.374 1.886 12.406 ;
			RECT	5.164 12.358 5.196 12.422 ;
			RECT	50.379 12.374 50.443 12.406 ;
			RECT	51.274 12.358 51.306 12.422 ;
			RECT	51.794 12.374 51.826 12.406 ;
			RECT	53.707 12.374 53.739 12.406 ;
			RECT	54.676 12.358 54.708 12.422 ;
			RECT	55.232 12.374 55.264 12.406 ;
			RECT	56.136 12.358 56.168 12.422 ;
			RECT	56.668 12.358 56.7 12.422 ;
			RECT	57.531 12.374 57.595 12.406 ;
			RECT	148.377 12.374 148.441 12.406 ;
			RECT	149.272 12.358 149.304 12.422 ;
			RECT	149.792 12.374 149.824 12.406 ;
			RECT	151.705 12.374 151.737 12.406 ;
			RECT	152.674 12.358 152.706 12.422 ;
			RECT	153.23 12.374 153.262 12.406 ;
			RECT	154.134 12.358 154.166 12.422 ;
			RECT	154.666 12.358 154.698 12.422 ;
			RECT	155.529 12.374 155.593 12.406 ;
			RECT	201.004 12.358 201.036 12.422 ;
			RECT	201.306 12.358 201.338 12.422 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 10.415 201.665 10.525 ;
			LAYER	J3 ;
			RECT	1.822 10.454 1.886 10.486 ;
			RECT	5.164 10.438 5.196 10.502 ;
			RECT	50.379 10.454 50.443 10.486 ;
			RECT	51.274 10.438 51.306 10.502 ;
			RECT	51.794 10.454 51.826 10.486 ;
			RECT	53.707 10.454 53.739 10.486 ;
			RECT	54.676 10.438 54.708 10.502 ;
			RECT	55.232 10.454 55.264 10.486 ;
			RECT	56.136 10.438 56.168 10.502 ;
			RECT	56.668 10.438 56.7 10.502 ;
			RECT	57.531 10.454 57.595 10.486 ;
			RECT	148.377 10.454 148.441 10.486 ;
			RECT	149.272 10.438 149.304 10.502 ;
			RECT	149.792 10.454 149.824 10.486 ;
			RECT	151.705 10.454 151.737 10.486 ;
			RECT	152.674 10.438 152.706 10.502 ;
			RECT	153.23 10.454 153.262 10.486 ;
			RECT	154.134 10.438 154.166 10.502 ;
			RECT	154.666 10.438 154.698 10.502 ;
			RECT	155.529 10.454 155.593 10.486 ;
			RECT	201.004 10.438 201.036 10.502 ;
			RECT	201.306 10.438 201.338 10.502 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 8.495 201.665 8.605 ;
			LAYER	J3 ;
			RECT	1.822 8.534 1.886 8.566 ;
			RECT	5.164 8.518 5.196 8.582 ;
			RECT	50.379 8.534 50.443 8.566 ;
			RECT	51.274 8.518 51.306 8.582 ;
			RECT	51.794 8.534 51.826 8.566 ;
			RECT	53.707 8.534 53.739 8.566 ;
			RECT	54.676 8.518 54.708 8.582 ;
			RECT	55.232 8.534 55.264 8.566 ;
			RECT	56.136 8.518 56.168 8.582 ;
			RECT	56.668 8.518 56.7 8.582 ;
			RECT	57.531 8.534 57.595 8.566 ;
			RECT	148.377 8.534 148.441 8.566 ;
			RECT	149.272 8.518 149.304 8.582 ;
			RECT	149.792 8.534 149.824 8.566 ;
			RECT	151.705 8.534 151.737 8.566 ;
			RECT	152.674 8.518 152.706 8.582 ;
			RECT	153.23 8.534 153.262 8.566 ;
			RECT	154.134 8.518 154.166 8.582 ;
			RECT	154.666 8.518 154.698 8.582 ;
			RECT	155.529 8.534 155.593 8.566 ;
			RECT	201.004 8.518 201.036 8.582 ;
			RECT	201.306 8.518 201.338 8.582 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 6.575 201.665 6.685 ;
			LAYER	J3 ;
			RECT	1.822 6.614 1.886 6.646 ;
			RECT	5.164 6.598 5.196 6.662 ;
			RECT	50.379 6.614 50.443 6.646 ;
			RECT	51.274 6.598 51.306 6.662 ;
			RECT	51.794 6.614 51.826 6.646 ;
			RECT	53.707 6.614 53.739 6.646 ;
			RECT	54.676 6.598 54.708 6.662 ;
			RECT	55.232 6.614 55.264 6.646 ;
			RECT	56.136 6.598 56.168 6.662 ;
			RECT	56.668 6.598 56.7 6.662 ;
			RECT	57.531 6.614 57.595 6.646 ;
			RECT	148.377 6.614 148.441 6.646 ;
			RECT	149.272 6.598 149.304 6.662 ;
			RECT	149.792 6.614 149.824 6.646 ;
			RECT	151.705 6.614 151.737 6.646 ;
			RECT	152.674 6.598 152.706 6.662 ;
			RECT	153.23 6.614 153.262 6.646 ;
			RECT	154.134 6.598 154.166 6.662 ;
			RECT	154.666 6.598 154.698 6.662 ;
			RECT	155.529 6.614 155.593 6.646 ;
			RECT	201.004 6.598 201.036 6.662 ;
			RECT	201.306 6.598 201.338 6.662 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 4.655 201.665 4.765 ;
			LAYER	J3 ;
			RECT	1.822 4.694 1.886 4.726 ;
			RECT	5.164 4.678 5.196 4.742 ;
			RECT	50.379 4.694 50.443 4.726 ;
			RECT	51.274 4.678 51.306 4.742 ;
			RECT	51.794 4.694 51.826 4.726 ;
			RECT	53.707 4.694 53.739 4.726 ;
			RECT	54.676 4.678 54.708 4.742 ;
			RECT	55.232 4.694 55.264 4.726 ;
			RECT	56.136 4.678 56.168 4.742 ;
			RECT	56.668 4.678 56.7 4.742 ;
			RECT	57.531 4.694 57.595 4.726 ;
			RECT	148.377 4.694 148.441 4.726 ;
			RECT	149.272 4.678 149.304 4.742 ;
			RECT	149.792 4.694 149.824 4.726 ;
			RECT	151.705 4.694 151.737 4.726 ;
			RECT	152.674 4.678 152.706 4.742 ;
			RECT	153.23 4.694 153.262 4.726 ;
			RECT	154.134 4.678 154.166 4.742 ;
			RECT	154.666 4.678 154.698 4.742 ;
			RECT	155.529 4.694 155.593 4.726 ;
			RECT	201.004 4.678 201.036 4.742 ;
			RECT	201.306 4.678 201.338 4.742 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 2.735 201.665 2.845 ;
			LAYER	J3 ;
			RECT	1.822 2.774 1.886 2.806 ;
			RECT	5.164 2.758 5.196 2.822 ;
			RECT	50.379 2.774 50.443 2.806 ;
			RECT	51.274 2.758 51.306 2.822 ;
			RECT	51.794 2.774 51.826 2.806 ;
			RECT	53.707 2.774 53.739 2.806 ;
			RECT	54.676 2.758 54.708 2.822 ;
			RECT	55.232 2.774 55.264 2.806 ;
			RECT	56.136 2.758 56.168 2.822 ;
			RECT	56.668 2.758 56.7 2.822 ;
			RECT	57.531 2.774 57.595 2.806 ;
			RECT	148.377 2.774 148.441 2.806 ;
			RECT	149.272 2.758 149.304 2.822 ;
			RECT	149.792 2.774 149.824 2.806 ;
			RECT	151.705 2.774 151.737 2.806 ;
			RECT	152.674 2.758 152.706 2.822 ;
			RECT	153.23 2.774 153.262 2.806 ;
			RECT	154.134 2.758 154.166 2.822 ;
			RECT	154.666 2.758 154.698 2.822 ;
			RECT	155.529 2.774 155.593 2.806 ;
			RECT	201.004 2.758 201.036 2.822 ;
			RECT	201.306 2.758 201.338 2.822 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 0.815 201.665 0.925 ;
			LAYER	J3 ;
			RECT	1.822 0.854 1.886 0.886 ;
			RECT	5.164 0.838 5.196 0.902 ;
			RECT	50.379 0.854 50.443 0.886 ;
			RECT	51.274 0.838 51.306 0.902 ;
			RECT	51.794 0.854 51.826 0.886 ;
			RECT	53.707 0.854 53.739 0.886 ;
			RECT	54.676 0.838 54.708 0.902 ;
			RECT	55.232 0.854 55.264 0.886 ;
			RECT	56.136 0.838 56.168 0.902 ;
			RECT	56.668 0.838 56.7 0.902 ;
			RECT	57.531 0.854 57.595 0.886 ;
			RECT	148.377 0.854 148.441 0.886 ;
			RECT	149.272 0.838 149.304 0.902 ;
			RECT	149.792 0.854 149.824 0.886 ;
			RECT	151.705 0.854 151.737 0.886 ;
			RECT	152.674 0.838 152.706 0.902 ;
			RECT	153.23 0.854 153.262 0.886 ;
			RECT	154.134 0.838 154.166 0.902 ;
			RECT	154.666 0.838 154.698 0.902 ;
			RECT	155.529 0.854 155.593 0.886 ;
			RECT	201.004 0.838 201.036 0.902 ;
			RECT	201.306 0.838 201.338 0.902 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 73.571 201.665 73.681 ;
			LAYER	J3 ;
			RECT	1.822 73.61 1.886 73.642 ;
			RECT	5.164 73.594 5.196 73.658 ;
			RECT	50.379 73.61 50.443 73.642 ;
			RECT	51.274 73.594 51.306 73.658 ;
			RECT	51.794 73.61 51.826 73.642 ;
			RECT	53.707 73.61 53.739 73.642 ;
			RECT	54.676 73.594 54.708 73.658 ;
			RECT	55.232 73.61 55.264 73.642 ;
			RECT	56.136 73.594 56.168 73.658 ;
			RECT	56.668 73.594 56.7 73.658 ;
			RECT	57.531 73.61 57.595 73.642 ;
			RECT	148.377 73.61 148.441 73.642 ;
			RECT	149.272 73.594 149.304 73.658 ;
			RECT	149.792 73.61 149.824 73.642 ;
			RECT	151.705 73.61 151.737 73.642 ;
			RECT	152.674 73.594 152.706 73.658 ;
			RECT	153.23 73.61 153.262 73.642 ;
			RECT	154.134 73.594 154.166 73.658 ;
			RECT	154.666 73.594 154.698 73.658 ;
			RECT	155.529 73.61 155.593 73.642 ;
			RECT	201.004 73.594 201.036 73.658 ;
			RECT	201.306 73.594 201.338 73.658 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 71.651 201.665 71.761 ;
			LAYER	J3 ;
			RECT	1.822 71.69 1.886 71.722 ;
			RECT	5.164 71.674 5.196 71.738 ;
			RECT	50.379 71.69 50.443 71.722 ;
			RECT	51.274 71.674 51.306 71.738 ;
			RECT	51.794 71.69 51.826 71.722 ;
			RECT	53.707 71.69 53.739 71.722 ;
			RECT	54.676 71.674 54.708 71.738 ;
			RECT	55.232 71.69 55.264 71.722 ;
			RECT	56.136 71.674 56.168 71.738 ;
			RECT	56.668 71.674 56.7 71.738 ;
			RECT	57.531 71.69 57.595 71.722 ;
			RECT	148.377 71.69 148.441 71.722 ;
			RECT	149.272 71.674 149.304 71.738 ;
			RECT	149.792 71.69 149.824 71.722 ;
			RECT	151.705 71.69 151.737 71.722 ;
			RECT	152.674 71.674 152.706 71.738 ;
			RECT	153.23 71.69 153.262 71.722 ;
			RECT	154.134 71.674 154.166 71.738 ;
			RECT	154.666 71.674 154.698 71.738 ;
			RECT	155.529 71.69 155.593 71.722 ;
			RECT	201.004 71.674 201.036 71.738 ;
			RECT	201.306 71.674 201.338 71.738 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 69.731 201.665 69.841 ;
			LAYER	J3 ;
			RECT	1.822 69.77 1.886 69.802 ;
			RECT	5.164 69.754 5.196 69.818 ;
			RECT	50.379 69.77 50.443 69.802 ;
			RECT	51.274 69.754 51.306 69.818 ;
			RECT	51.794 69.77 51.826 69.802 ;
			RECT	53.707 69.77 53.739 69.802 ;
			RECT	54.676 69.754 54.708 69.818 ;
			RECT	55.232 69.77 55.264 69.802 ;
			RECT	56.136 69.754 56.168 69.818 ;
			RECT	56.668 69.754 56.7 69.818 ;
			RECT	57.531 69.77 57.595 69.802 ;
			RECT	148.377 69.77 148.441 69.802 ;
			RECT	149.272 69.754 149.304 69.818 ;
			RECT	149.792 69.77 149.824 69.802 ;
			RECT	151.705 69.77 151.737 69.802 ;
			RECT	152.674 69.754 152.706 69.818 ;
			RECT	153.23 69.77 153.262 69.802 ;
			RECT	154.134 69.754 154.166 69.818 ;
			RECT	154.666 69.754 154.698 69.818 ;
			RECT	155.529 69.77 155.593 69.802 ;
			RECT	201.004 69.754 201.036 69.818 ;
			RECT	201.306 69.754 201.338 69.818 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 67.811 201.665 67.921 ;
			LAYER	J3 ;
			RECT	1.822 67.85 1.886 67.882 ;
			RECT	5.164 67.834 5.196 67.898 ;
			RECT	50.379 67.85 50.443 67.882 ;
			RECT	51.274 67.834 51.306 67.898 ;
			RECT	51.794 67.85 51.826 67.882 ;
			RECT	53.707 67.85 53.739 67.882 ;
			RECT	54.676 67.834 54.708 67.898 ;
			RECT	55.232 67.85 55.264 67.882 ;
			RECT	56.136 67.834 56.168 67.898 ;
			RECT	56.668 67.834 56.7 67.898 ;
			RECT	57.531 67.85 57.595 67.882 ;
			RECT	148.377 67.85 148.441 67.882 ;
			RECT	149.272 67.834 149.304 67.898 ;
			RECT	149.792 67.85 149.824 67.882 ;
			RECT	151.705 67.85 151.737 67.882 ;
			RECT	152.674 67.834 152.706 67.898 ;
			RECT	153.23 67.85 153.262 67.882 ;
			RECT	154.134 67.834 154.166 67.898 ;
			RECT	154.666 67.834 154.698 67.898 ;
			RECT	155.529 67.85 155.593 67.882 ;
			RECT	201.004 67.834 201.036 67.898 ;
			RECT	201.306 67.834 201.338 67.898 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 65.891 201.665 66.001 ;
			LAYER	J3 ;
			RECT	1.822 65.93 1.886 65.962 ;
			RECT	5.164 65.914 5.196 65.978 ;
			RECT	50.379 65.93 50.443 65.962 ;
			RECT	51.274 65.914 51.306 65.978 ;
			RECT	51.794 65.93 51.826 65.962 ;
			RECT	53.707 65.93 53.739 65.962 ;
			RECT	54.676 65.914 54.708 65.978 ;
			RECT	55.232 65.93 55.264 65.962 ;
			RECT	56.136 65.914 56.168 65.978 ;
			RECT	56.668 65.914 56.7 65.978 ;
			RECT	57.531 65.93 57.595 65.962 ;
			RECT	148.377 65.93 148.441 65.962 ;
			RECT	149.272 65.914 149.304 65.978 ;
			RECT	149.792 65.93 149.824 65.962 ;
			RECT	151.705 65.93 151.737 65.962 ;
			RECT	152.674 65.914 152.706 65.978 ;
			RECT	153.23 65.93 153.262 65.962 ;
			RECT	154.134 65.914 154.166 65.978 ;
			RECT	154.666 65.914 154.698 65.978 ;
			RECT	155.529 65.93 155.593 65.962 ;
			RECT	201.004 65.914 201.036 65.978 ;
			RECT	201.306 65.914 201.338 65.978 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 63.971 201.665 64.081 ;
			LAYER	J3 ;
			RECT	1.822 64.01 1.886 64.042 ;
			RECT	5.164 63.994 5.196 64.058 ;
			RECT	50.379 64.01 50.443 64.042 ;
			RECT	51.274 63.994 51.306 64.058 ;
			RECT	51.794 64.01 51.826 64.042 ;
			RECT	53.707 64.01 53.739 64.042 ;
			RECT	54.676 63.994 54.708 64.058 ;
			RECT	55.232 64.01 55.264 64.042 ;
			RECT	56.136 63.994 56.168 64.058 ;
			RECT	56.668 63.994 56.7 64.058 ;
			RECT	57.531 64.01 57.595 64.042 ;
			RECT	148.377 64.01 148.441 64.042 ;
			RECT	149.272 63.994 149.304 64.058 ;
			RECT	149.792 64.01 149.824 64.042 ;
			RECT	151.705 64.01 151.737 64.042 ;
			RECT	152.674 63.994 152.706 64.058 ;
			RECT	153.23 64.01 153.262 64.042 ;
			RECT	154.134 63.994 154.166 64.058 ;
			RECT	154.666 63.994 154.698 64.058 ;
			RECT	155.529 64.01 155.593 64.042 ;
			RECT	201.004 63.994 201.036 64.058 ;
			RECT	201.306 63.994 201.338 64.058 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 62.051 201.665 62.161 ;
			LAYER	J3 ;
			RECT	1.822 62.09 1.886 62.122 ;
			RECT	5.164 62.074 5.196 62.138 ;
			RECT	50.379 62.09 50.443 62.122 ;
			RECT	51.274 62.074 51.306 62.138 ;
			RECT	51.794 62.09 51.826 62.122 ;
			RECT	53.707 62.09 53.739 62.122 ;
			RECT	54.676 62.074 54.708 62.138 ;
			RECT	55.232 62.09 55.264 62.122 ;
			RECT	56.136 62.074 56.168 62.138 ;
			RECT	56.668 62.074 56.7 62.138 ;
			RECT	57.531 62.09 57.595 62.122 ;
			RECT	148.377 62.09 148.441 62.122 ;
			RECT	149.272 62.074 149.304 62.138 ;
			RECT	149.792 62.09 149.824 62.122 ;
			RECT	151.705 62.09 151.737 62.122 ;
			RECT	152.674 62.074 152.706 62.138 ;
			RECT	153.23 62.09 153.262 62.122 ;
			RECT	154.134 62.074 154.166 62.138 ;
			RECT	154.666 62.074 154.698 62.138 ;
			RECT	155.529 62.09 155.593 62.122 ;
			RECT	201.004 62.074 201.036 62.138 ;
			RECT	201.306 62.074 201.338 62.138 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 60.131 201.665 60.241 ;
			LAYER	J3 ;
			RECT	1.822 60.17 1.886 60.202 ;
			RECT	5.164 60.154 5.196 60.218 ;
			RECT	50.379 60.17 50.443 60.202 ;
			RECT	51.274 60.154 51.306 60.218 ;
			RECT	51.794 60.17 51.826 60.202 ;
			RECT	53.707 60.17 53.739 60.202 ;
			RECT	54.676 60.154 54.708 60.218 ;
			RECT	55.232 60.17 55.264 60.202 ;
			RECT	56.136 60.154 56.168 60.218 ;
			RECT	56.668 60.154 56.7 60.218 ;
			RECT	57.531 60.17 57.595 60.202 ;
			RECT	148.377 60.17 148.441 60.202 ;
			RECT	149.272 60.154 149.304 60.218 ;
			RECT	149.792 60.17 149.824 60.202 ;
			RECT	151.705 60.17 151.737 60.202 ;
			RECT	152.674 60.154 152.706 60.218 ;
			RECT	153.23 60.17 153.262 60.202 ;
			RECT	154.134 60.154 154.166 60.218 ;
			RECT	154.666 60.154 154.698 60.218 ;
			RECT	155.529 60.17 155.593 60.202 ;
			RECT	201.004 60.154 201.036 60.218 ;
			RECT	201.306 60.154 201.338 60.218 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 58.211 201.665 58.321 ;
			LAYER	J3 ;
			RECT	1.822 58.25 1.886 58.282 ;
			RECT	5.164 58.234 5.196 58.298 ;
			RECT	50.379 58.25 50.443 58.282 ;
			RECT	51.274 58.234 51.306 58.298 ;
			RECT	51.794 58.25 51.826 58.282 ;
			RECT	53.707 58.25 53.739 58.282 ;
			RECT	54.676 58.234 54.708 58.298 ;
			RECT	55.232 58.25 55.264 58.282 ;
			RECT	56.136 58.234 56.168 58.298 ;
			RECT	56.668 58.234 56.7 58.298 ;
			RECT	57.531 58.25 57.595 58.282 ;
			RECT	148.377 58.25 148.441 58.282 ;
			RECT	149.272 58.234 149.304 58.298 ;
			RECT	149.792 58.25 149.824 58.282 ;
			RECT	151.705 58.25 151.737 58.282 ;
			RECT	152.674 58.234 152.706 58.298 ;
			RECT	153.23 58.25 153.262 58.282 ;
			RECT	154.134 58.234 154.166 58.298 ;
			RECT	154.666 58.234 154.698 58.298 ;
			RECT	155.529 58.25 155.593 58.282 ;
			RECT	201.004 58.234 201.036 58.298 ;
			RECT	201.306 58.234 201.338 58.298 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 56.291 201.665 56.401 ;
			LAYER	J3 ;
			RECT	1.822 56.33 1.886 56.362 ;
			RECT	5.164 56.314 5.196 56.378 ;
			RECT	50.379 56.33 50.443 56.362 ;
			RECT	51.274 56.314 51.306 56.378 ;
			RECT	51.794 56.33 51.826 56.362 ;
			RECT	53.707 56.33 53.739 56.362 ;
			RECT	54.676 56.314 54.708 56.378 ;
			RECT	55.232 56.33 55.264 56.362 ;
			RECT	56.136 56.314 56.168 56.378 ;
			RECT	56.668 56.314 56.7 56.378 ;
			RECT	57.531 56.33 57.595 56.362 ;
			RECT	148.377 56.33 148.441 56.362 ;
			RECT	149.272 56.314 149.304 56.378 ;
			RECT	149.792 56.33 149.824 56.362 ;
			RECT	151.705 56.33 151.737 56.362 ;
			RECT	152.674 56.314 152.706 56.378 ;
			RECT	153.23 56.33 153.262 56.362 ;
			RECT	154.134 56.314 154.166 56.378 ;
			RECT	154.666 56.314 154.698 56.378 ;
			RECT	155.529 56.33 155.593 56.362 ;
			RECT	201.004 56.314 201.036 56.378 ;
			RECT	201.306 56.314 201.338 56.378 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 54.371 201.665 54.481 ;
			LAYER	J3 ;
			RECT	1.822 54.41 1.886 54.442 ;
			RECT	5.164 54.394 5.196 54.458 ;
			RECT	50.379 54.41 50.443 54.442 ;
			RECT	51.274 54.394 51.306 54.458 ;
			RECT	51.794 54.41 51.826 54.442 ;
			RECT	53.707 54.41 53.739 54.442 ;
			RECT	54.676 54.394 54.708 54.458 ;
			RECT	55.232 54.41 55.264 54.442 ;
			RECT	56.136 54.394 56.168 54.458 ;
			RECT	56.668 54.394 56.7 54.458 ;
			RECT	57.531 54.41 57.595 54.442 ;
			RECT	148.377 54.41 148.441 54.442 ;
			RECT	149.272 54.394 149.304 54.458 ;
			RECT	149.792 54.41 149.824 54.442 ;
			RECT	151.705 54.41 151.737 54.442 ;
			RECT	152.674 54.394 152.706 54.458 ;
			RECT	153.23 54.41 153.262 54.442 ;
			RECT	154.134 54.394 154.166 54.458 ;
			RECT	154.666 54.394 154.698 54.458 ;
			RECT	155.529 54.41 155.593 54.442 ;
			RECT	201.004 54.394 201.036 54.458 ;
			RECT	201.306 54.394 201.338 54.458 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 52.451 201.665 52.561 ;
			LAYER	J3 ;
			RECT	1.822 52.49 1.886 52.522 ;
			RECT	5.164 52.474 5.196 52.538 ;
			RECT	50.379 52.49 50.443 52.522 ;
			RECT	51.274 52.474 51.306 52.538 ;
			RECT	51.794 52.49 51.826 52.522 ;
			RECT	53.707 52.49 53.739 52.522 ;
			RECT	54.676 52.474 54.708 52.538 ;
			RECT	55.232 52.49 55.264 52.522 ;
			RECT	56.136 52.474 56.168 52.538 ;
			RECT	56.668 52.474 56.7 52.538 ;
			RECT	57.531 52.49 57.595 52.522 ;
			RECT	148.377 52.49 148.441 52.522 ;
			RECT	149.272 52.474 149.304 52.538 ;
			RECT	149.792 52.49 149.824 52.522 ;
			RECT	151.705 52.49 151.737 52.522 ;
			RECT	152.674 52.474 152.706 52.538 ;
			RECT	153.23 52.49 153.262 52.522 ;
			RECT	154.134 52.474 154.166 52.538 ;
			RECT	154.666 52.474 154.698 52.538 ;
			RECT	155.529 52.49 155.593 52.522 ;
			RECT	201.004 52.474 201.036 52.538 ;
			RECT	201.306 52.474 201.338 52.538 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 79.331 201.665 79.441 ;
			LAYER	J3 ;
			RECT	1.822 79.37 1.886 79.402 ;
			RECT	5.164 79.354 5.196 79.418 ;
			RECT	50.379 79.37 50.443 79.402 ;
			RECT	51.274 79.354 51.306 79.418 ;
			RECT	51.794 79.37 51.826 79.402 ;
			RECT	53.707 79.37 53.739 79.402 ;
			RECT	54.676 79.354 54.708 79.418 ;
			RECT	55.232 79.37 55.264 79.402 ;
			RECT	56.136 79.354 56.168 79.418 ;
			RECT	56.668 79.354 56.7 79.418 ;
			RECT	57.531 79.37 57.595 79.402 ;
			RECT	148.377 79.37 148.441 79.402 ;
			RECT	149.272 79.354 149.304 79.418 ;
			RECT	149.792 79.37 149.824 79.402 ;
			RECT	151.705 79.37 151.737 79.402 ;
			RECT	152.674 79.354 152.706 79.418 ;
			RECT	153.23 79.37 153.262 79.402 ;
			RECT	154.134 79.354 154.166 79.418 ;
			RECT	154.666 79.354 154.698 79.418 ;
			RECT	155.529 79.37 155.593 79.402 ;
			RECT	201.004 79.354 201.036 79.418 ;
			RECT	201.306 79.354 201.338 79.418 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 32.468 201.665 32.578 ;
			LAYER	J3 ;
			RECT	1.822 32.491 1.886 32.555 ;
			RECT	2.501 32.491 2.565 32.555 ;
			RECT	3.922 32.491 3.954 32.555 ;
			RECT	4.113 32.491 4.145 32.555 ;
			RECT	4.674 32.491 4.706 32.555 ;
			RECT	5.164 32.491 5.196 32.555 ;
			RECT	50.412 32.491 50.444 32.555 ;
			RECT	51.274 32.491 51.306 32.555 ;
			RECT	51.794 32.491 51.826 32.555 ;
			RECT	55.216 32.491 55.248 32.555 ;
			RECT	56.144 32.491 56.176 32.555 ;
			RECT	56.664 32.491 56.696 32.555 ;
			RECT	57.254 32.491 57.286 32.555 ;
			RECT	57.531 32.491 57.595 32.555 ;
			RECT	148.41 32.491 148.442 32.555 ;
			RECT	149.272 32.491 149.304 32.555 ;
			RECT	149.792 32.491 149.824 32.555 ;
			RECT	153.214 32.491 153.246 32.555 ;
			RECT	154.142 32.491 154.174 32.555 ;
			RECT	154.662 32.491 154.694 32.555 ;
			RECT	155.252 32.491 155.284 32.555 ;
			RECT	155.529 32.491 155.593 32.555 ;
			RECT	201.307 32.491 201.339 32.555 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 34.227 201.665 34.347 ;
			LAYER	J3 ;
			RECT	0.812 34.255 0.844 34.319 ;
			RECT	1.024 34.255 1.056 34.319 ;
			RECT	1.822 34.255 1.886 34.319 ;
			RECT	2.501 34.255 2.565 34.319 ;
			RECT	3.922 34.255 3.954 34.319 ;
			RECT	4.113 34.255 4.145 34.319 ;
			RECT	4.674 34.255 4.706 34.319 ;
			RECT	5.164 34.255 5.196 34.319 ;
			RECT	50.412 34.255 50.444 34.319 ;
			RECT	51.274 34.255 51.306 34.319 ;
			RECT	51.794 34.255 51.826 34.319 ;
			RECT	53.403 34.255 53.435 34.319 ;
			RECT	55.208 34.255 55.272 34.319 ;
			RECT	56.144 34.255 56.176 34.319 ;
			RECT	56.664 34.255 56.696 34.319 ;
			RECT	57.495 34.255 57.527 34.319 ;
			RECT	148.41 34.255 148.442 34.319 ;
			RECT	149.272 34.255 149.304 34.319 ;
			RECT	149.792 34.255 149.824 34.319 ;
			RECT	151.401 34.255 151.433 34.319 ;
			RECT	153.206 34.255 153.27 34.319 ;
			RECT	154.142 34.255 154.174 34.319 ;
			RECT	154.662 34.255 154.694 34.319 ;
			RECT	155.493 34.255 155.525 34.319 ;
			RECT	201.307 34.255 201.339 34.319 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 35.022 201.665 35.142 ;
			LAYER	J3 ;
			RECT	1.024 35.05 1.056 35.114 ;
			RECT	1.822 35.05 1.886 35.114 ;
			RECT	1.981 35.05 2.013 35.114 ;
			RECT	2.501 35.05 2.565 35.114 ;
			RECT	3.285 35.05 3.317 35.114 ;
			RECT	3.695 35.05 3.727 35.114 ;
			RECT	3.922 35.05 3.954 35.114 ;
			RECT	5.164 35.05 5.196 35.114 ;
			RECT	48.844 35.05 48.876 35.114 ;
			RECT	50.412 35.05 50.444 35.114 ;
			RECT	51.274 35.05 51.306 35.114 ;
			RECT	51.794 35.05 51.826 35.114 ;
			RECT	52.597 35.05 52.629 35.114 ;
			RECT	53.403 35.05 53.435 35.114 ;
			RECT	55.208 35.05 55.272 35.114 ;
			RECT	56.144 35.05 56.176 35.114 ;
			RECT	56.664 35.05 56.696 35.114 ;
			RECT	57.495 35.05 57.527 35.114 ;
			RECT	59.328 35.05 59.36 35.114 ;
			RECT	146.842 35.05 146.874 35.114 ;
			RECT	148.41 35.05 148.442 35.114 ;
			RECT	149.272 35.05 149.304 35.114 ;
			RECT	149.792 35.05 149.824 35.114 ;
			RECT	150.595 35.05 150.627 35.114 ;
			RECT	151.401 35.05 151.433 35.114 ;
			RECT	153.206 35.05 153.27 35.114 ;
			RECT	154.142 35.05 154.174 35.114 ;
			RECT	154.662 35.05 154.694 35.114 ;
			RECT	155.493 35.05 155.525 35.114 ;
			RECT	157.326 35.05 157.358 35.114 ;
			RECT	201.004 35.05 201.036 35.114 ;
			RECT	201.307 35.05 201.339 35.114 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 36.064 201.665 36.154 ;
			LAYER	J3 ;
			RECT	1.024 36.077 1.056 36.141 ;
			RECT	1.838 36.077 1.87 36.141 ;
			RECT	1.981 36.077 2.013 36.141 ;
			RECT	2.501 36.093 2.565 36.125 ;
			RECT	3.285 36.077 3.317 36.141 ;
			RECT	3.695 36.093 3.727 36.125 ;
			RECT	3.922 36.077 3.954 36.141 ;
			RECT	5.164 36.077 5.196 36.141 ;
			RECT	48.844 36.077 48.876 36.141 ;
			RECT	50.412 36.077 50.444 36.141 ;
			RECT	51.274 36.077 51.306 36.141 ;
			RECT	51.794 36.077 51.826 36.141 ;
			RECT	52.597 36.077 52.629 36.141 ;
			RECT	53.403 36.077 53.435 36.141 ;
			RECT	55.224 36.077 55.256 36.141 ;
			RECT	56.144 36.077 56.176 36.141 ;
			RECT	56.664 36.077 56.696 36.141 ;
			RECT	57.495 36.077 57.527 36.141 ;
			RECT	59.328 36.077 59.36 36.141 ;
			RECT	146.842 36.077 146.874 36.141 ;
			RECT	148.41 36.077 148.442 36.141 ;
			RECT	149.272 36.077 149.304 36.141 ;
			RECT	149.792 36.077 149.824 36.141 ;
			RECT	150.595 36.077 150.627 36.141 ;
			RECT	151.401 36.077 151.433 36.141 ;
			RECT	153.222 36.077 153.254 36.141 ;
			RECT	154.142 36.077 154.174 36.141 ;
			RECT	154.662 36.077 154.694 36.141 ;
			RECT	155.493 36.077 155.525 36.141 ;
			RECT	157.326 36.077 157.358 36.141 ;
			RECT	201.004 36.077 201.036 36.141 ;
			RECT	201.307 36.077 201.339 36.141 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 37.05 201.665 37.17 ;
			LAYER	J3 ;
			RECT	1.024 37.078 1.056 37.142 ;
			RECT	1.822 37.078 1.886 37.142 ;
			RECT	1.981 37.078 2.013 37.142 ;
			RECT	2.501 37.078 2.565 37.142 ;
			RECT	2.956 37.078 2.988 37.142 ;
			RECT	3.285 37.078 3.317 37.142 ;
			RECT	3.695 37.078 3.727 37.142 ;
			RECT	3.922 37.078 3.954 37.142 ;
			RECT	4.277 37.078 4.309 37.142 ;
			RECT	5.164 37.078 5.196 37.142 ;
			RECT	5.567 37.078 5.599 37.142 ;
			RECT	48.844 37.078 48.876 37.142 ;
			RECT	50.412 37.078 50.444 37.142 ;
			RECT	51.274 37.078 51.306 37.142 ;
			RECT	51.794 37.078 51.826 37.142 ;
			RECT	52.597 37.078 52.629 37.142 ;
			RECT	53.403 37.078 53.435 37.142 ;
			RECT	54.066 37.094 54.098 37.126 ;
			RECT	54.363 37.078 54.427 37.142 ;
			RECT	55.208 37.078 55.272 37.142 ;
			RECT	56.144 37.078 56.176 37.142 ;
			RECT	56.664 37.078 56.696 37.142 ;
			RECT	57.495 37.078 57.527 37.142 ;
			RECT	59.328 37.078 59.36 37.142 ;
			RECT	102.605 37.078 102.637 37.142 ;
			RECT	103.565 37.078 103.597 37.142 ;
			RECT	146.842 37.078 146.874 37.142 ;
			RECT	148.41 37.078 148.442 37.142 ;
			RECT	149.272 37.078 149.304 37.142 ;
			RECT	149.792 37.078 149.824 37.142 ;
			RECT	150.595 37.078 150.627 37.142 ;
			RECT	151.401 37.078 151.433 37.142 ;
			RECT	152.064 37.094 152.096 37.126 ;
			RECT	152.361 37.078 152.425 37.142 ;
			RECT	153.206 37.078 153.27 37.142 ;
			RECT	154.142 37.078 154.174 37.142 ;
			RECT	154.662 37.078 154.694 37.142 ;
			RECT	155.493 37.078 155.525 37.142 ;
			RECT	157.326 37.078 157.358 37.142 ;
			RECT	200.603 37.078 200.635 37.142 ;
			RECT	201.307 37.078 201.339 37.142 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 37.815 201.665 37.905 ;
			LAYER	J3 ;
			RECT	1.024 37.828 1.056 37.892 ;
			RECT	1.838 37.828 1.87 37.892 ;
			RECT	1.981 37.828 2.013 37.892 ;
			RECT	2.517 37.828 2.549 37.892 ;
			RECT	2.957 37.828 2.989 37.892 ;
			RECT	3.285 37.828 3.317 37.892 ;
			RECT	3.922 37.828 3.954 37.892 ;
			RECT	4.277 37.828 4.309 37.892 ;
			RECT	5.567 37.828 5.599 37.892 ;
			RECT	35.952 37.844 35.984 37.876 ;
			RECT	36.624 37.844 36.656 37.876 ;
			RECT	37.296 37.844 37.328 37.876 ;
			RECT	39.312 37.844 39.344 37.876 ;
			RECT	40.656 37.844 40.688 37.876 ;
			RECT	41.328 37.844 41.36 37.876 ;
			RECT	48.844 37.828 48.876 37.892 ;
			RECT	50.434 37.828 50.466 37.892 ;
			RECT	51.274 37.828 51.306 37.892 ;
			RECT	51.794 37.828 51.826 37.892 ;
			RECT	52.597 37.828 52.629 37.892 ;
			RECT	53.403 37.828 53.435 37.892 ;
			RECT	54.379 37.828 54.411 37.892 ;
			RECT	55.224 37.828 55.256 37.892 ;
			RECT	56.144 37.827 56.176 37.891 ;
			RECT	56.664 37.828 56.696 37.892 ;
			RECT	57.495 37.828 57.527 37.892 ;
			RECT	57.766 37.828 57.798 37.892 ;
			RECT	59.328 37.828 59.36 37.892 ;
			RECT	66.844 37.844 66.876 37.876 ;
			RECT	67.516 37.844 67.548 37.876 ;
			RECT	68.86 37.844 68.892 37.876 ;
			RECT	70.876 37.844 70.908 37.876 ;
			RECT	71.548 37.844 71.58 37.876 ;
			RECT	72.22 37.844 72.252 37.876 ;
			RECT	102.605 37.828 102.637 37.892 ;
			RECT	103.565 37.828 103.597 37.892 ;
			RECT	133.95 37.844 133.982 37.876 ;
			RECT	134.622 37.844 134.654 37.876 ;
			RECT	135.294 37.844 135.326 37.876 ;
			RECT	137.31 37.844 137.342 37.876 ;
			RECT	138.654 37.844 138.686 37.876 ;
			RECT	139.326 37.844 139.358 37.876 ;
			RECT	146.842 37.828 146.874 37.892 ;
			RECT	148.432 37.828 148.464 37.892 ;
			RECT	149.272 37.828 149.304 37.892 ;
			RECT	149.792 37.828 149.824 37.892 ;
			RECT	150.595 37.828 150.627 37.892 ;
			RECT	151.401 37.828 151.433 37.892 ;
			RECT	152.377 37.828 152.409 37.892 ;
			RECT	153.222 37.828 153.254 37.892 ;
			RECT	154.142 37.827 154.174 37.891 ;
			RECT	154.662 37.828 154.694 37.892 ;
			RECT	155.493 37.828 155.525 37.892 ;
			RECT	155.764 37.828 155.796 37.892 ;
			RECT	157.326 37.828 157.358 37.892 ;
			RECT	164.842 37.844 164.874 37.876 ;
			RECT	165.514 37.844 165.546 37.876 ;
			RECT	166.858 37.844 166.89 37.876 ;
			RECT	168.874 37.844 168.906 37.876 ;
			RECT	169.546 37.844 169.578 37.876 ;
			RECT	170.218 37.844 170.25 37.876 ;
			RECT	200.603 37.828 200.635 37.892 ;
			RECT	201.307 37.828 201.339 37.892 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 38.187 201.665 38.277 ;
			LAYER	J3 ;
			RECT	1.024 38.204 1.056 38.236 ;
			RECT	1.838 38.2 1.87 38.264 ;
			RECT	1.981 38.2 2.013 38.264 ;
			RECT	2.501 38.216 2.565 38.248 ;
			RECT	2.957 38.2 2.989 38.264 ;
			RECT	3.285 38.2 3.317 38.264 ;
			RECT	3.922 38.2 3.954 38.264 ;
			RECT	4.277 38.2 4.309 38.264 ;
			RECT	4.982 38.216 5.014 38.248 ;
			RECT	5.164 38.2 5.196 38.264 ;
			RECT	27.888 38.2 27.92 38.264 ;
			RECT	28.56 38.2 28.592 38.264 ;
			RECT	29.232 38.2 29.264 38.264 ;
			RECT	29.904 38.2 29.936 38.264 ;
			RECT	30.912 38.2 30.944 38.264 ;
			RECT	31.584 38.2 31.616 38.264 ;
			RECT	34.608 38.2 34.64 38.264 ;
			RECT	34.944 38.2 34.976 38.264 ;
			RECT	35.952 38.2 35.984 38.264 ;
			RECT	36.624 38.2 36.656 38.264 ;
			RECT	37.296 38.2 37.328 38.264 ;
			RECT	37.968 38.2 38 38.264 ;
			RECT	38.304 38.2 38.336 38.264 ;
			RECT	38.976 38.2 39.008 38.264 ;
			RECT	39.312 38.2 39.344 38.264 ;
			RECT	40.656 38.2 40.688 38.264 ;
			RECT	41.328 38.2 41.36 38.264 ;
			RECT	41.664 38.2 41.696 38.264 ;
			RECT	43.344 38.2 43.376 38.264 ;
			RECT	46.032 38.2 46.064 38.264 ;
			RECT	47.376 38.2 47.408 38.264 ;
			RECT	48.844 38.2 48.876 38.264 ;
			RECT	50.434 38.2 50.466 38.264 ;
			RECT	51.274 38.2 51.306 38.264 ;
			RECT	51.794 38.2 51.826 38.264 ;
			RECT	52.597 38.2 52.629 38.264 ;
			RECT	53.403 38.2 53.435 38.264 ;
			RECT	53.996 38.2 54.028 38.264 ;
			RECT	54.379 38.2 54.411 38.264 ;
			RECT	55.224 38.2 55.256 38.264 ;
			RECT	56.144 38.2 56.176 38.264 ;
			RECT	56.664 38.201 56.696 38.265 ;
			RECT	57.509 38.216 57.573 38.248 ;
			RECT	59.328 38.2 59.36 38.264 ;
			RECT	60.796 38.2 60.828 38.264 ;
			RECT	62.14 38.2 62.172 38.264 ;
			RECT	64.828 38.2 64.86 38.264 ;
			RECT	66.508 38.2 66.54 38.264 ;
			RECT	66.844 38.2 66.876 38.264 ;
			RECT	67.516 38.2 67.548 38.264 ;
			RECT	68.86 38.2 68.892 38.264 ;
			RECT	69.196 38.2 69.228 38.264 ;
			RECT	69.868 38.2 69.9 38.264 ;
			RECT	70.204 38.2 70.236 38.264 ;
			RECT	70.876 38.2 70.908 38.264 ;
			RECT	71.548 38.2 71.58 38.264 ;
			RECT	72.22 38.2 72.252 38.264 ;
			RECT	73.228 38.2 73.26 38.264 ;
			RECT	73.564 38.2 73.596 38.264 ;
			RECT	76.588 38.2 76.62 38.264 ;
			RECT	77.26 38.2 77.292 38.264 ;
			RECT	78.268 38.2 78.3 38.264 ;
			RECT	78.94 38.2 78.972 38.264 ;
			RECT	79.612 38.2 79.644 38.264 ;
			RECT	80.284 38.2 80.316 38.264 ;
			RECT	125.886 38.2 125.918 38.264 ;
			RECT	126.558 38.2 126.59 38.264 ;
			RECT	127.23 38.2 127.262 38.264 ;
			RECT	127.902 38.2 127.934 38.264 ;
			RECT	128.91 38.2 128.942 38.264 ;
			RECT	129.582 38.2 129.614 38.264 ;
			RECT	132.606 38.2 132.638 38.264 ;
			RECT	132.942 38.2 132.974 38.264 ;
			RECT	133.95 38.2 133.982 38.264 ;
			RECT	134.622 38.2 134.654 38.264 ;
			RECT	135.294 38.2 135.326 38.264 ;
			RECT	135.966 38.2 135.998 38.264 ;
			RECT	136.302 38.2 136.334 38.264 ;
			RECT	136.974 38.2 137.006 38.264 ;
			RECT	137.31 38.2 137.342 38.264 ;
			RECT	138.654 38.2 138.686 38.264 ;
			RECT	139.326 38.2 139.358 38.264 ;
			RECT	139.662 38.2 139.694 38.264 ;
			RECT	141.342 38.2 141.374 38.264 ;
			RECT	144.03 38.2 144.062 38.264 ;
			RECT	145.374 38.2 145.406 38.264 ;
			RECT	146.842 38.2 146.874 38.264 ;
			RECT	148.432 38.2 148.464 38.264 ;
			RECT	149.272 38.2 149.304 38.264 ;
			RECT	149.792 38.2 149.824 38.264 ;
			RECT	150.595 38.2 150.627 38.264 ;
			RECT	151.401 38.2 151.433 38.264 ;
			RECT	151.994 38.2 152.026 38.264 ;
			RECT	152.377 38.2 152.409 38.264 ;
			RECT	153.222 38.2 153.254 38.264 ;
			RECT	154.142 38.2 154.174 38.264 ;
			RECT	154.662 38.201 154.694 38.265 ;
			RECT	155.507 38.216 155.571 38.248 ;
			RECT	157.326 38.2 157.358 38.264 ;
			RECT	158.794 38.2 158.826 38.264 ;
			RECT	160.138 38.2 160.17 38.264 ;
			RECT	162.826 38.2 162.858 38.264 ;
			RECT	164.506 38.2 164.538 38.264 ;
			RECT	164.842 38.2 164.874 38.264 ;
			RECT	165.514 38.2 165.546 38.264 ;
			RECT	166.858 38.2 166.89 38.264 ;
			RECT	167.194 38.2 167.226 38.264 ;
			RECT	167.866 38.2 167.898 38.264 ;
			RECT	168.202 38.2 168.234 38.264 ;
			RECT	168.874 38.2 168.906 38.264 ;
			RECT	169.546 38.2 169.578 38.264 ;
			RECT	170.218 38.2 170.25 38.264 ;
			RECT	171.226 38.2 171.258 38.264 ;
			RECT	171.562 38.2 171.594 38.264 ;
			RECT	174.586 38.2 174.618 38.264 ;
			RECT	175.258 38.2 175.29 38.264 ;
			RECT	176.266 38.2 176.298 38.264 ;
			RECT	176.938 38.2 176.97 38.264 ;
			RECT	177.61 38.2 177.642 38.264 ;
			RECT	178.282 38.2 178.314 38.264 ;
			RECT	201.307 38.2 201.339 38.264 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 38.777 201.665 38.897 ;
			LAYER	J3 ;
			RECT	1.024 38.805 1.056 38.869 ;
			RECT	1.822 38.805 1.886 38.869 ;
			RECT	1.981 38.805 2.013 38.869 ;
			RECT	2.501 38.805 2.565 38.869 ;
			RECT	2.952 38.805 2.984 38.869 ;
			RECT	3.922 38.805 3.954 38.869 ;
			RECT	4.277 38.805 4.309 38.869 ;
			RECT	4.982 38.805 5.014 38.869 ;
			RECT	5.164 38.805 5.196 38.869 ;
			RECT	6.389 38.805 6.421 38.869 ;
			RECT	6.725 38.805 6.757 38.869 ;
			RECT	7.061 38.805 7.093 38.869 ;
			RECT	7.397 38.805 7.429 38.869 ;
			RECT	7.733 38.805 7.765 38.869 ;
			RECT	8.069 38.805 8.101 38.869 ;
			RECT	8.405 38.805 8.437 38.869 ;
			RECT	8.741 38.805 8.773 38.869 ;
			RECT	9.077 38.805 9.109 38.869 ;
			RECT	9.413 38.805 9.445 38.869 ;
			RECT	9.749 38.805 9.781 38.869 ;
			RECT	10.085 38.805 10.117 38.869 ;
			RECT	10.421 38.805 10.453 38.869 ;
			RECT	10.757 38.805 10.789 38.869 ;
			RECT	11.093 38.805 11.125 38.869 ;
			RECT	11.429 38.805 11.461 38.869 ;
			RECT	11.765 38.805 11.797 38.869 ;
			RECT	12.101 38.805 12.133 38.869 ;
			RECT	12.437 38.805 12.469 38.869 ;
			RECT	12.773 38.805 12.805 38.869 ;
			RECT	13.109 38.805 13.141 38.869 ;
			RECT	13.445 38.805 13.477 38.869 ;
			RECT	13.781 38.805 13.813 38.869 ;
			RECT	14.117 38.805 14.149 38.869 ;
			RECT	14.453 38.805 14.485 38.869 ;
			RECT	14.789 38.805 14.821 38.869 ;
			RECT	15.125 38.805 15.157 38.869 ;
			RECT	15.461 38.805 15.493 38.869 ;
			RECT	15.797 38.805 15.829 38.869 ;
			RECT	16.133 38.805 16.165 38.869 ;
			RECT	16.469 38.805 16.501 38.869 ;
			RECT	16.805 38.805 16.837 38.869 ;
			RECT	17.141 38.805 17.173 38.869 ;
			RECT	17.477 38.805 17.509 38.869 ;
			RECT	17.813 38.805 17.845 38.869 ;
			RECT	18.149 38.805 18.181 38.869 ;
			RECT	18.485 38.805 18.517 38.869 ;
			RECT	18.821 38.805 18.853 38.869 ;
			RECT	19.157 38.805 19.189 38.869 ;
			RECT	19.493 38.805 19.525 38.869 ;
			RECT	19.829 38.805 19.861 38.869 ;
			RECT	20.165 38.805 20.197 38.869 ;
			RECT	20.501 38.805 20.533 38.869 ;
			RECT	20.837 38.805 20.869 38.869 ;
			RECT	21.173 38.805 21.205 38.869 ;
			RECT	21.509 38.805 21.541 38.869 ;
			RECT	21.845 38.805 21.877 38.869 ;
			RECT	22.181 38.805 22.213 38.869 ;
			RECT	22.517 38.805 22.549 38.869 ;
			RECT	22.853 38.805 22.885 38.869 ;
			RECT	23.189 38.805 23.221 38.869 ;
			RECT	23.525 38.805 23.557 38.869 ;
			RECT	23.861 38.805 23.893 38.869 ;
			RECT	24.197 38.805 24.229 38.869 ;
			RECT	24.533 38.805 24.565 38.869 ;
			RECT	24.869 38.805 24.901 38.869 ;
			RECT	25.205 38.805 25.237 38.869 ;
			RECT	25.541 38.805 25.573 38.869 ;
			RECT	25.877 38.805 25.909 38.869 ;
			RECT	26.213 38.805 26.245 38.869 ;
			RECT	26.549 38.805 26.581 38.869 ;
			RECT	26.885 38.805 26.917 38.869 ;
			RECT	27.221 38.805 27.253 38.869 ;
			RECT	27.557 38.805 27.589 38.869 ;
			RECT	27.888 38.805 27.92 38.869 ;
			RECT	28.224 38.805 28.256 38.869 ;
			RECT	28.56 38.805 28.592 38.869 ;
			RECT	29.232 38.805 29.264 38.869 ;
			RECT	29.568 38.805 29.6 38.869 ;
			RECT	29.904 38.805 29.936 38.869 ;
			RECT	30.912 38.805 30.944 38.869 ;
			RECT	31.584 38.805 31.616 38.869 ;
			RECT	32.256 38.805 32.288 38.869 ;
			RECT	32.928 38.805 32.96 38.869 ;
			RECT	33.6 38.805 33.632 38.869 ;
			RECT	34.608 38.805 34.64 38.869 ;
			RECT	34.944 38.805 34.976 38.869 ;
			RECT	37.296 38.805 37.328 38.869 ;
			RECT	37.968 38.805 38 38.869 ;
			RECT	38.304 38.805 38.336 38.869 ;
			RECT	38.976 38.805 39.008 38.869 ;
			RECT	39.312 38.805 39.344 38.869 ;
			RECT	41.664 38.805 41.696 38.869 ;
			RECT	42 38.805 42.032 38.869 ;
			RECT	43.008 38.805 43.04 38.869 ;
			RECT	43.344 38.805 43.376 38.869 ;
			RECT	44.016 38.805 44.048 38.869 ;
			RECT	44.352 38.805 44.384 38.869 ;
			RECT	44.688 38.805 44.72 38.869 ;
			RECT	45.024 38.805 45.056 38.869 ;
			RECT	45.696 38.805 45.728 38.869 ;
			RECT	46.032 38.805 46.064 38.869 ;
			RECT	47.376 38.805 47.408 38.869 ;
			RECT	48.844 38.805 48.876 38.869 ;
			RECT	50.418 38.805 50.482 38.869 ;
			RECT	51.274 38.805 51.306 38.869 ;
			RECT	51.794 38.805 51.826 38.869 ;
			RECT	52.597 38.805 52.629 38.869 ;
			RECT	53.403 38.821 53.435 38.853 ;
			RECT	53.996 38.821 54.028 38.853 ;
			RECT	56.664 38.805 56.696 38.869 ;
			RECT	57.509 38.805 57.573 38.869 ;
			RECT	57.766 38.805 57.798 38.869 ;
			RECT	59.328 38.805 59.36 38.869 ;
			RECT	60.796 38.805 60.828 38.869 ;
			RECT	62.14 38.805 62.172 38.869 ;
			RECT	62.476 38.805 62.508 38.869 ;
			RECT	63.148 38.805 63.18 38.869 ;
			RECT	63.484 38.805 63.516 38.869 ;
			RECT	63.82 38.805 63.852 38.869 ;
			RECT	64.156 38.805 64.188 38.869 ;
			RECT	64.828 38.805 64.86 38.869 ;
			RECT	65.164 38.805 65.196 38.869 ;
			RECT	66.172 38.805 66.204 38.869 ;
			RECT	66.508 38.805 66.54 38.869 ;
			RECT	68.86 38.805 68.892 38.869 ;
			RECT	69.196 38.805 69.228 38.869 ;
			RECT	69.868 38.805 69.9 38.869 ;
			RECT	70.204 38.805 70.236 38.869 ;
			RECT	70.876 38.805 70.908 38.869 ;
			RECT	73.228 38.805 73.26 38.869 ;
			RECT	73.564 38.805 73.596 38.869 ;
			RECT	74.572 38.805 74.604 38.869 ;
			RECT	75.244 38.805 75.276 38.869 ;
			RECT	75.916 38.805 75.948 38.869 ;
			RECT	76.588 38.805 76.62 38.869 ;
			RECT	77.26 38.805 77.292 38.869 ;
			RECT	78.268 38.805 78.3 38.869 ;
			RECT	78.604 38.805 78.636 38.869 ;
			RECT	78.94 38.805 78.972 38.869 ;
			RECT	79.612 38.805 79.644 38.869 ;
			RECT	79.948 38.805 79.98 38.869 ;
			RECT	80.284 38.805 80.316 38.869 ;
			RECT	80.615 38.805 80.647 38.869 ;
			RECT	80.951 38.805 80.983 38.869 ;
			RECT	81.287 38.805 81.319 38.869 ;
			RECT	81.623 38.805 81.655 38.869 ;
			RECT	81.959 38.805 81.991 38.869 ;
			RECT	82.295 38.805 82.327 38.869 ;
			RECT	82.631 38.805 82.663 38.869 ;
			RECT	82.967 38.805 82.999 38.869 ;
			RECT	83.303 38.805 83.335 38.869 ;
			RECT	83.639 38.805 83.671 38.869 ;
			RECT	83.975 38.805 84.007 38.869 ;
			RECT	84.311 38.805 84.343 38.869 ;
			RECT	84.647 38.805 84.679 38.869 ;
			RECT	84.983 38.805 85.015 38.869 ;
			RECT	85.319 38.805 85.351 38.869 ;
			RECT	85.655 38.805 85.687 38.869 ;
			RECT	85.991 38.805 86.023 38.869 ;
			RECT	86.327 38.805 86.359 38.869 ;
			RECT	86.663 38.805 86.695 38.869 ;
			RECT	86.999 38.805 87.031 38.869 ;
			RECT	87.335 38.805 87.367 38.869 ;
			RECT	87.671 38.805 87.703 38.869 ;
			RECT	88.007 38.805 88.039 38.869 ;
			RECT	88.343 38.805 88.375 38.869 ;
			RECT	88.679 38.805 88.711 38.869 ;
			RECT	89.015 38.805 89.047 38.869 ;
			RECT	89.351 38.805 89.383 38.869 ;
			RECT	89.687 38.805 89.719 38.869 ;
			RECT	90.023 38.805 90.055 38.869 ;
			RECT	90.359 38.805 90.391 38.869 ;
			RECT	90.695 38.805 90.727 38.869 ;
			RECT	91.031 38.805 91.063 38.869 ;
			RECT	91.367 38.805 91.399 38.869 ;
			RECT	91.703 38.805 91.735 38.869 ;
			RECT	92.039 38.805 92.071 38.869 ;
			RECT	92.375 38.805 92.407 38.869 ;
			RECT	92.711 38.805 92.743 38.869 ;
			RECT	93.047 38.805 93.079 38.869 ;
			RECT	93.383 38.805 93.415 38.869 ;
			RECT	93.719 38.805 93.751 38.869 ;
			RECT	94.055 38.805 94.087 38.869 ;
			RECT	94.391 38.805 94.423 38.869 ;
			RECT	94.727 38.805 94.759 38.869 ;
			RECT	95.063 38.805 95.095 38.869 ;
			RECT	95.399 38.805 95.431 38.869 ;
			RECT	95.735 38.805 95.767 38.869 ;
			RECT	96.071 38.805 96.103 38.869 ;
			RECT	96.407 38.805 96.439 38.869 ;
			RECT	96.743 38.805 96.775 38.869 ;
			RECT	97.079 38.805 97.111 38.869 ;
			RECT	97.415 38.805 97.447 38.869 ;
			RECT	97.751 38.805 97.783 38.869 ;
			RECT	98.087 38.805 98.119 38.869 ;
			RECT	98.423 38.805 98.455 38.869 ;
			RECT	98.759 38.805 98.791 38.869 ;
			RECT	99.095 38.805 99.127 38.869 ;
			RECT	99.431 38.805 99.463 38.869 ;
			RECT	99.767 38.805 99.799 38.869 ;
			RECT	100.103 38.805 100.135 38.869 ;
			RECT	100.439 38.805 100.471 38.869 ;
			RECT	100.775 38.805 100.807 38.869 ;
			RECT	101.111 38.805 101.143 38.869 ;
			RECT	101.447 38.805 101.479 38.869 ;
			RECT	101.783 38.805 101.815 38.869 ;
			RECT	104.387 38.805 104.419 38.869 ;
			RECT	104.723 38.805 104.755 38.869 ;
			RECT	105.059 38.805 105.091 38.869 ;
			RECT	105.395 38.805 105.427 38.869 ;
			RECT	105.731 38.805 105.763 38.869 ;
			RECT	106.067 38.805 106.099 38.869 ;
			RECT	106.403 38.805 106.435 38.869 ;
			RECT	106.739 38.805 106.771 38.869 ;
			RECT	107.075 38.805 107.107 38.869 ;
			RECT	107.411 38.805 107.443 38.869 ;
			RECT	107.747 38.805 107.779 38.869 ;
			RECT	108.083 38.805 108.115 38.869 ;
			RECT	108.419 38.805 108.451 38.869 ;
			RECT	108.755 38.805 108.787 38.869 ;
			RECT	109.091 38.805 109.123 38.869 ;
			RECT	109.427 38.805 109.459 38.869 ;
			RECT	109.763 38.805 109.795 38.869 ;
			RECT	110.099 38.805 110.131 38.869 ;
			RECT	110.435 38.805 110.467 38.869 ;
			RECT	110.771 38.805 110.803 38.869 ;
			RECT	111.107 38.805 111.139 38.869 ;
			RECT	111.443 38.805 111.475 38.869 ;
			RECT	111.779 38.805 111.811 38.869 ;
			RECT	112.115 38.805 112.147 38.869 ;
			RECT	112.451 38.805 112.483 38.869 ;
			RECT	112.787 38.805 112.819 38.869 ;
			RECT	113.123 38.805 113.155 38.869 ;
			RECT	113.459 38.805 113.491 38.869 ;
			RECT	113.795 38.805 113.827 38.869 ;
			RECT	114.131 38.805 114.163 38.869 ;
			RECT	114.467 38.805 114.499 38.869 ;
			RECT	114.803 38.805 114.835 38.869 ;
			RECT	115.139 38.805 115.171 38.869 ;
			RECT	115.475 38.805 115.507 38.869 ;
			RECT	115.811 38.805 115.843 38.869 ;
			RECT	116.147 38.805 116.179 38.869 ;
			RECT	116.483 38.805 116.515 38.869 ;
			RECT	116.819 38.805 116.851 38.869 ;
			RECT	117.155 38.805 117.187 38.869 ;
			RECT	117.491 38.805 117.523 38.869 ;
			RECT	117.827 38.805 117.859 38.869 ;
			RECT	118.163 38.805 118.195 38.869 ;
			RECT	118.499 38.805 118.531 38.869 ;
			RECT	118.835 38.805 118.867 38.869 ;
			RECT	119.171 38.805 119.203 38.869 ;
			RECT	119.507 38.805 119.539 38.869 ;
			RECT	119.843 38.805 119.875 38.869 ;
			RECT	120.179 38.805 120.211 38.869 ;
			RECT	120.515 38.805 120.547 38.869 ;
			RECT	120.851 38.805 120.883 38.869 ;
			RECT	121.187 38.805 121.219 38.869 ;
			RECT	121.523 38.805 121.555 38.869 ;
			RECT	121.859 38.805 121.891 38.869 ;
			RECT	122.195 38.805 122.227 38.869 ;
			RECT	122.531 38.805 122.563 38.869 ;
			RECT	122.867 38.805 122.899 38.869 ;
			RECT	123.203 38.805 123.235 38.869 ;
			RECT	123.539 38.805 123.571 38.869 ;
			RECT	123.875 38.805 123.907 38.869 ;
			RECT	124.211 38.805 124.243 38.869 ;
			RECT	124.547 38.805 124.579 38.869 ;
			RECT	124.883 38.805 124.915 38.869 ;
			RECT	125.219 38.805 125.251 38.869 ;
			RECT	125.555 38.805 125.587 38.869 ;
			RECT	125.886 38.805 125.918 38.869 ;
			RECT	126.222 38.805 126.254 38.869 ;
			RECT	126.558 38.805 126.59 38.869 ;
			RECT	127.23 38.805 127.262 38.869 ;
			RECT	127.566 38.805 127.598 38.869 ;
			RECT	127.902 38.805 127.934 38.869 ;
			RECT	128.91 38.805 128.942 38.869 ;
			RECT	129.582 38.805 129.614 38.869 ;
			RECT	130.254 38.805 130.286 38.869 ;
			RECT	130.926 38.805 130.958 38.869 ;
			RECT	131.598 38.805 131.63 38.869 ;
			RECT	132.606 38.805 132.638 38.869 ;
			RECT	132.942 38.805 132.974 38.869 ;
			RECT	135.294 38.805 135.326 38.869 ;
			RECT	135.966 38.805 135.998 38.869 ;
			RECT	136.302 38.805 136.334 38.869 ;
			RECT	136.974 38.805 137.006 38.869 ;
			RECT	137.31 38.805 137.342 38.869 ;
			RECT	139.662 38.805 139.694 38.869 ;
			RECT	139.998 38.805 140.03 38.869 ;
			RECT	141.006 38.805 141.038 38.869 ;
			RECT	141.342 38.805 141.374 38.869 ;
			RECT	142.014 38.805 142.046 38.869 ;
			RECT	142.35 38.805 142.382 38.869 ;
			RECT	142.686 38.805 142.718 38.869 ;
			RECT	143.022 38.805 143.054 38.869 ;
			RECT	143.694 38.805 143.726 38.869 ;
			RECT	144.03 38.805 144.062 38.869 ;
			RECT	145.374 38.805 145.406 38.869 ;
			RECT	146.842 38.805 146.874 38.869 ;
			RECT	148.416 38.805 148.48 38.869 ;
			RECT	149.272 38.805 149.304 38.869 ;
			RECT	149.792 38.805 149.824 38.869 ;
			RECT	150.595 38.805 150.627 38.869 ;
			RECT	151.401 38.821 151.433 38.853 ;
			RECT	151.994 38.821 152.026 38.853 ;
			RECT	154.662 38.805 154.694 38.869 ;
			RECT	155.507 38.805 155.571 38.869 ;
			RECT	155.764 38.805 155.796 38.869 ;
			RECT	157.326 38.805 157.358 38.869 ;
			RECT	158.794 38.805 158.826 38.869 ;
			RECT	160.138 38.805 160.17 38.869 ;
			RECT	160.474 38.805 160.506 38.869 ;
			RECT	161.146 38.805 161.178 38.869 ;
			RECT	161.482 38.805 161.514 38.869 ;
			RECT	161.818 38.805 161.85 38.869 ;
			RECT	162.154 38.805 162.186 38.869 ;
			RECT	162.826 38.805 162.858 38.869 ;
			RECT	163.162 38.805 163.194 38.869 ;
			RECT	164.17 38.805 164.202 38.869 ;
			RECT	164.506 38.805 164.538 38.869 ;
			RECT	166.858 38.805 166.89 38.869 ;
			RECT	167.194 38.805 167.226 38.869 ;
			RECT	167.866 38.805 167.898 38.869 ;
			RECT	168.202 38.805 168.234 38.869 ;
			RECT	168.874 38.805 168.906 38.869 ;
			RECT	171.226 38.805 171.258 38.869 ;
			RECT	171.562 38.805 171.594 38.869 ;
			RECT	172.57 38.805 172.602 38.869 ;
			RECT	173.242 38.805 173.274 38.869 ;
			RECT	173.914 38.805 173.946 38.869 ;
			RECT	174.586 38.805 174.618 38.869 ;
			RECT	175.258 38.805 175.29 38.869 ;
			RECT	176.266 38.805 176.298 38.869 ;
			RECT	176.602 38.805 176.634 38.869 ;
			RECT	176.938 38.805 176.97 38.869 ;
			RECT	177.61 38.805 177.642 38.869 ;
			RECT	177.946 38.805 177.978 38.869 ;
			RECT	178.282 38.805 178.314 38.869 ;
			RECT	178.613 38.805 178.645 38.869 ;
			RECT	178.949 38.805 178.981 38.869 ;
			RECT	179.285 38.805 179.317 38.869 ;
			RECT	179.621 38.805 179.653 38.869 ;
			RECT	179.957 38.805 179.989 38.869 ;
			RECT	180.293 38.805 180.325 38.869 ;
			RECT	180.629 38.805 180.661 38.869 ;
			RECT	180.965 38.805 180.997 38.869 ;
			RECT	181.301 38.805 181.333 38.869 ;
			RECT	181.637 38.805 181.669 38.869 ;
			RECT	181.973 38.805 182.005 38.869 ;
			RECT	182.309 38.805 182.341 38.869 ;
			RECT	182.645 38.805 182.677 38.869 ;
			RECT	182.981 38.805 183.013 38.869 ;
			RECT	183.317 38.805 183.349 38.869 ;
			RECT	183.653 38.805 183.685 38.869 ;
			RECT	183.989 38.805 184.021 38.869 ;
			RECT	184.325 38.805 184.357 38.869 ;
			RECT	184.661 38.805 184.693 38.869 ;
			RECT	184.997 38.805 185.029 38.869 ;
			RECT	185.333 38.805 185.365 38.869 ;
			RECT	185.669 38.805 185.701 38.869 ;
			RECT	186.005 38.805 186.037 38.869 ;
			RECT	186.341 38.805 186.373 38.869 ;
			RECT	186.677 38.805 186.709 38.869 ;
			RECT	187.013 38.805 187.045 38.869 ;
			RECT	187.349 38.805 187.381 38.869 ;
			RECT	187.685 38.805 187.717 38.869 ;
			RECT	188.021 38.805 188.053 38.869 ;
			RECT	188.357 38.805 188.389 38.869 ;
			RECT	188.693 38.805 188.725 38.869 ;
			RECT	189.029 38.805 189.061 38.869 ;
			RECT	189.365 38.805 189.397 38.869 ;
			RECT	189.701 38.805 189.733 38.869 ;
			RECT	190.037 38.805 190.069 38.869 ;
			RECT	190.373 38.805 190.405 38.869 ;
			RECT	190.709 38.805 190.741 38.869 ;
			RECT	191.045 38.805 191.077 38.869 ;
			RECT	191.381 38.805 191.413 38.869 ;
			RECT	191.717 38.805 191.749 38.869 ;
			RECT	192.053 38.805 192.085 38.869 ;
			RECT	192.389 38.805 192.421 38.869 ;
			RECT	192.725 38.805 192.757 38.869 ;
			RECT	193.061 38.805 193.093 38.869 ;
			RECT	193.397 38.805 193.429 38.869 ;
			RECT	193.733 38.805 193.765 38.869 ;
			RECT	194.069 38.805 194.101 38.869 ;
			RECT	194.405 38.805 194.437 38.869 ;
			RECT	194.741 38.805 194.773 38.869 ;
			RECT	195.077 38.805 195.109 38.869 ;
			RECT	195.413 38.805 195.445 38.869 ;
			RECT	195.749 38.805 195.781 38.869 ;
			RECT	196.085 38.805 196.117 38.869 ;
			RECT	196.421 38.805 196.453 38.869 ;
			RECT	196.757 38.805 196.789 38.869 ;
			RECT	197.093 38.805 197.125 38.869 ;
			RECT	197.429 38.805 197.461 38.869 ;
			RECT	197.765 38.805 197.797 38.869 ;
			RECT	198.101 38.805 198.133 38.869 ;
			RECT	198.437 38.805 198.469 38.869 ;
			RECT	198.773 38.805 198.805 38.869 ;
			RECT	199.109 38.805 199.141 38.869 ;
			RECT	199.445 38.805 199.477 38.869 ;
			RECT	199.781 38.805 199.813 38.869 ;
			RECT	201.307 38.805 201.339 38.869 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 39.974 201.665 40.064 ;
			LAYER	J3 ;
			RECT	1.024 39.987 1.056 40.051 ;
			RECT	1.838 39.987 1.87 40.051 ;
			RECT	1.981 39.987 2.013 40.051 ;
			RECT	2.517 39.987 2.549 40.051 ;
			RECT	2.953 39.987 2.985 40.051 ;
			RECT	3.922 39.987 3.954 40.051 ;
			RECT	4.982 39.987 5.014 40.051 ;
			RECT	5.164 39.987 5.196 40.051 ;
			RECT	38.304 39.987 38.336 40.051 ;
			RECT	48.844 39.987 48.876 40.051 ;
			RECT	51.794 39.987 51.826 40.051 ;
			RECT	52.597 39.987 52.629 40.051 ;
			RECT	53.403 39.987 53.435 40.051 ;
			RECT	55.22 39.987 55.252 40.051 ;
			RECT	57.766 39.987 57.798 40.051 ;
			RECT	59.328 39.987 59.36 40.051 ;
			RECT	69.868 39.987 69.9 40.051 ;
			RECT	136.302 39.987 136.334 40.051 ;
			RECT	146.842 39.987 146.874 40.051 ;
			RECT	149.792 39.987 149.824 40.051 ;
			RECT	150.595 39.987 150.627 40.051 ;
			RECT	151.401 39.987 151.433 40.051 ;
			RECT	153.218 39.987 153.25 40.051 ;
			RECT	155.764 39.987 155.796 40.051 ;
			RECT	157.326 39.987 157.358 40.051 ;
			RECT	167.866 39.987 167.898 40.051 ;
			RECT	201.307 39.985 201.339 40.049 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 41.13 201.665 41.25 ;
			LAYER	J3 ;
			RECT	1.024 41.158 1.056 41.222 ;
			RECT	1.822 41.158 1.886 41.222 ;
			RECT	1.981 41.158 2.013 41.222 ;
			RECT	2.501 41.158 2.565 41.222 ;
			RECT	2.988 41.158 3.02 41.222 ;
			RECT	3.313 41.158 3.345 41.222 ;
			RECT	3.922 41.158 3.954 41.222 ;
			RECT	4.056 41.158 4.088 41.222 ;
			RECT	4.196 41.158 4.228 41.222 ;
			RECT	4.48 41.158 4.544 41.222 ;
			RECT	4.982 41.158 5.014 41.222 ;
			RECT	5.164 41.158 5.196 41.222 ;
			RECT	6.389 41.158 6.421 41.222 ;
			RECT	6.725 41.158 6.757 41.222 ;
			RECT	7.061 41.158 7.093 41.222 ;
			RECT	7.397 41.158 7.429 41.222 ;
			RECT	7.733 41.158 7.765 41.222 ;
			RECT	8.069 41.158 8.101 41.222 ;
			RECT	8.405 41.158 8.437 41.222 ;
			RECT	8.741 41.158 8.773 41.222 ;
			RECT	9.077 41.158 9.109 41.222 ;
			RECT	9.413 41.158 9.445 41.222 ;
			RECT	9.749 41.158 9.781 41.222 ;
			RECT	10.085 41.158 10.117 41.222 ;
			RECT	10.421 41.158 10.453 41.222 ;
			RECT	10.757 41.158 10.789 41.222 ;
			RECT	11.093 41.158 11.125 41.222 ;
			RECT	11.429 41.158 11.461 41.222 ;
			RECT	11.765 41.158 11.797 41.222 ;
			RECT	12.101 41.158 12.133 41.222 ;
			RECT	12.437 41.158 12.469 41.222 ;
			RECT	12.773 41.158 12.805 41.222 ;
			RECT	13.109 41.158 13.141 41.222 ;
			RECT	13.445 41.158 13.477 41.222 ;
			RECT	13.781 41.158 13.813 41.222 ;
			RECT	14.117 41.158 14.149 41.222 ;
			RECT	14.453 41.158 14.485 41.222 ;
			RECT	14.789 41.158 14.821 41.222 ;
			RECT	15.125 41.158 15.157 41.222 ;
			RECT	15.461 41.158 15.493 41.222 ;
			RECT	15.797 41.158 15.829 41.222 ;
			RECT	16.133 41.158 16.165 41.222 ;
			RECT	16.469 41.158 16.501 41.222 ;
			RECT	16.805 41.158 16.837 41.222 ;
			RECT	17.141 41.158 17.173 41.222 ;
			RECT	17.477 41.158 17.509 41.222 ;
			RECT	17.813 41.158 17.845 41.222 ;
			RECT	18.149 41.158 18.181 41.222 ;
			RECT	18.485 41.158 18.517 41.222 ;
			RECT	18.821 41.158 18.853 41.222 ;
			RECT	19.157 41.158 19.189 41.222 ;
			RECT	19.493 41.158 19.525 41.222 ;
			RECT	19.829 41.158 19.861 41.222 ;
			RECT	20.165 41.158 20.197 41.222 ;
			RECT	20.501 41.158 20.533 41.222 ;
			RECT	20.837 41.158 20.869 41.222 ;
			RECT	21.173 41.158 21.205 41.222 ;
			RECT	21.509 41.158 21.541 41.222 ;
			RECT	21.845 41.158 21.877 41.222 ;
			RECT	22.181 41.158 22.213 41.222 ;
			RECT	22.517 41.158 22.549 41.222 ;
			RECT	22.853 41.158 22.885 41.222 ;
			RECT	23.189 41.158 23.221 41.222 ;
			RECT	23.525 41.158 23.557 41.222 ;
			RECT	23.861 41.158 23.893 41.222 ;
			RECT	24.197 41.158 24.229 41.222 ;
			RECT	24.533 41.158 24.565 41.222 ;
			RECT	24.869 41.158 24.901 41.222 ;
			RECT	25.205 41.158 25.237 41.222 ;
			RECT	25.541 41.158 25.573 41.222 ;
			RECT	25.877 41.158 25.909 41.222 ;
			RECT	26.213 41.158 26.245 41.222 ;
			RECT	26.549 41.158 26.581 41.222 ;
			RECT	26.885 41.158 26.917 41.222 ;
			RECT	27.221 41.158 27.253 41.222 ;
			RECT	27.557 41.158 27.589 41.222 ;
			RECT	28.224 41.158 28.256 41.222 ;
			RECT	28.896 41.158 28.928 41.222 ;
			RECT	29.568 41.158 29.6 41.222 ;
			RECT	30.24 41.158 30.272 41.222 ;
			RECT	30.912 41.158 30.944 41.222 ;
			RECT	31.248 41.158 31.28 41.222 ;
			RECT	31.584 41.158 31.616 41.222 ;
			RECT	32.256 41.158 32.288 41.222 ;
			RECT	32.592 41.158 32.624 41.222 ;
			RECT	32.928 41.158 32.96 41.222 ;
			RECT	33.6 41.158 33.632 41.222 ;
			RECT	33.936 41.158 33.968 41.222 ;
			RECT	34.944 41.158 34.976 41.222 ;
			RECT	35.28 41.158 35.312 41.222 ;
			RECT	36.288 41.158 36.32 41.222 ;
			RECT	36.624 41.158 36.656 41.222 ;
			RECT	37.632 41.158 37.664 41.222 ;
			RECT	37.968 41.158 38 41.222 ;
			RECT	38.304 41.158 38.336 41.222 ;
			RECT	38.976 41.158 39.008 41.222 ;
			RECT	39.312 41.158 39.344 41.222 ;
			RECT	39.648 41.158 39.68 41.222 ;
			RECT	39.984 41.158 40.016 41.222 ;
			RECT	40.656 41.158 40.688 41.222 ;
			RECT	40.992 41.158 41.024 41.222 ;
			RECT	41.664 41.158 41.696 41.222 ;
			RECT	42 41.158 42.032 41.222 ;
			RECT	42.336 41.158 42.368 41.222 ;
			RECT	43.008 41.158 43.04 41.222 ;
			RECT	43.344 41.158 43.376 41.222 ;
			RECT	44.352 41.158 44.384 41.222 ;
			RECT	45.024 41.158 45.056 41.222 ;
			RECT	45.696 41.158 45.728 41.222 ;
			RECT	46.368 41.158 46.4 41.222 ;
			RECT	47.04 41.158 47.072 41.222 ;
			RECT	47.376 41.158 47.408 41.222 ;
			RECT	48.384 41.158 48.416 41.222 ;
			RECT	48.844 41.158 48.876 41.222 ;
			RECT	49.638 41.158 49.67 41.222 ;
			RECT	50.417 41.158 50.481 41.222 ;
			RECT	51.274 41.158 51.306 41.222 ;
			RECT	51.794 41.158 51.826 41.222 ;
			RECT	52.597 41.158 52.629 41.222 ;
			RECT	53.403 41.158 53.435 41.222 ;
			RECT	55.204 41.158 55.268 41.222 ;
			RECT	56.144 41.158 56.176 41.222 ;
			RECT	56.664 41.158 56.696 41.222 ;
			RECT	57.507 41.158 57.571 41.222 ;
			RECT	57.75 41.158 57.814 41.222 ;
			RECT	58.534 41.158 58.566 41.222 ;
			RECT	59.328 41.158 59.36 41.222 ;
			RECT	59.788 41.158 59.82 41.222 ;
			RECT	60.796 41.158 60.828 41.222 ;
			RECT	61.132 41.158 61.164 41.222 ;
			RECT	61.804 41.158 61.836 41.222 ;
			RECT	62.476 41.158 62.508 41.222 ;
			RECT	63.148 41.158 63.18 41.222 ;
			RECT	63.82 41.158 63.852 41.222 ;
			RECT	64.828 41.158 64.86 41.222 ;
			RECT	65.164 41.158 65.196 41.222 ;
			RECT	65.836 41.158 65.868 41.222 ;
			RECT	66.172 41.158 66.204 41.222 ;
			RECT	66.508 41.158 66.54 41.222 ;
			RECT	67.18 41.158 67.212 41.222 ;
			RECT	67.516 41.158 67.548 41.222 ;
			RECT	68.188 41.158 68.22 41.222 ;
			RECT	68.524 41.158 68.556 41.222 ;
			RECT	68.86 41.158 68.892 41.222 ;
			RECT	69.196 41.158 69.228 41.222 ;
			RECT	69.868 41.158 69.9 41.222 ;
			RECT	70.204 41.158 70.236 41.222 ;
			RECT	70.54 41.158 70.572 41.222 ;
			RECT	71.548 41.158 71.58 41.222 ;
			RECT	71.884 41.158 71.916 41.222 ;
			RECT	72.892 41.158 72.924 41.222 ;
			RECT	73.228 41.158 73.26 41.222 ;
			RECT	74.236 41.158 74.268 41.222 ;
			RECT	74.572 41.158 74.604 41.222 ;
			RECT	75.244 41.158 75.276 41.222 ;
			RECT	75.58 41.158 75.612 41.222 ;
			RECT	75.916 41.158 75.948 41.222 ;
			RECT	76.588 41.158 76.62 41.222 ;
			RECT	76.924 41.158 76.956 41.222 ;
			RECT	77.26 41.158 77.292 41.222 ;
			RECT	77.932 41.158 77.964 41.222 ;
			RECT	78.604 41.158 78.636 41.222 ;
			RECT	79.276 41.158 79.308 41.222 ;
			RECT	79.948 41.158 79.98 41.222 ;
			RECT	80.615 41.158 80.647 41.222 ;
			RECT	80.951 41.158 80.983 41.222 ;
			RECT	81.287 41.158 81.319 41.222 ;
			RECT	81.623 41.158 81.655 41.222 ;
			RECT	81.959 41.158 81.991 41.222 ;
			RECT	82.295 41.158 82.327 41.222 ;
			RECT	82.631 41.158 82.663 41.222 ;
			RECT	82.967 41.158 82.999 41.222 ;
			RECT	83.303 41.158 83.335 41.222 ;
			RECT	83.639 41.158 83.671 41.222 ;
			RECT	83.975 41.158 84.007 41.222 ;
			RECT	84.311 41.158 84.343 41.222 ;
			RECT	84.647 41.158 84.679 41.222 ;
			RECT	84.983 41.158 85.015 41.222 ;
			RECT	85.319 41.158 85.351 41.222 ;
			RECT	85.655 41.158 85.687 41.222 ;
			RECT	85.991 41.158 86.023 41.222 ;
			RECT	86.327 41.158 86.359 41.222 ;
			RECT	86.663 41.158 86.695 41.222 ;
			RECT	86.999 41.158 87.031 41.222 ;
			RECT	87.335 41.158 87.367 41.222 ;
			RECT	87.671 41.158 87.703 41.222 ;
			RECT	88.007 41.158 88.039 41.222 ;
			RECT	88.343 41.158 88.375 41.222 ;
			RECT	88.679 41.158 88.711 41.222 ;
			RECT	89.015 41.158 89.047 41.222 ;
			RECT	89.351 41.158 89.383 41.222 ;
			RECT	89.687 41.158 89.719 41.222 ;
			RECT	90.023 41.158 90.055 41.222 ;
			RECT	90.359 41.158 90.391 41.222 ;
			RECT	90.695 41.158 90.727 41.222 ;
			RECT	91.031 41.158 91.063 41.222 ;
			RECT	91.367 41.158 91.399 41.222 ;
			RECT	91.703 41.158 91.735 41.222 ;
			RECT	92.039 41.158 92.071 41.222 ;
			RECT	92.375 41.158 92.407 41.222 ;
			RECT	92.711 41.158 92.743 41.222 ;
			RECT	93.047 41.158 93.079 41.222 ;
			RECT	93.383 41.158 93.415 41.222 ;
			RECT	93.719 41.158 93.751 41.222 ;
			RECT	94.055 41.158 94.087 41.222 ;
			RECT	94.391 41.158 94.423 41.222 ;
			RECT	94.727 41.158 94.759 41.222 ;
			RECT	95.063 41.158 95.095 41.222 ;
			RECT	95.399 41.158 95.431 41.222 ;
			RECT	95.735 41.158 95.767 41.222 ;
			RECT	96.071 41.158 96.103 41.222 ;
			RECT	96.407 41.158 96.439 41.222 ;
			RECT	96.743 41.158 96.775 41.222 ;
			RECT	97.079 41.158 97.111 41.222 ;
			RECT	97.415 41.158 97.447 41.222 ;
			RECT	97.751 41.158 97.783 41.222 ;
			RECT	98.087 41.158 98.119 41.222 ;
			RECT	98.423 41.158 98.455 41.222 ;
			RECT	98.759 41.158 98.791 41.222 ;
			RECT	99.095 41.158 99.127 41.222 ;
			RECT	99.431 41.158 99.463 41.222 ;
			RECT	99.767 41.158 99.799 41.222 ;
			RECT	100.103 41.158 100.135 41.222 ;
			RECT	100.439 41.158 100.471 41.222 ;
			RECT	100.775 41.158 100.807 41.222 ;
			RECT	101.111 41.158 101.143 41.222 ;
			RECT	101.447 41.158 101.479 41.222 ;
			RECT	101.783 41.158 101.815 41.222 ;
			RECT	104.387 41.158 104.419 41.222 ;
			RECT	104.723 41.158 104.755 41.222 ;
			RECT	105.059 41.158 105.091 41.222 ;
			RECT	105.395 41.158 105.427 41.222 ;
			RECT	105.731 41.158 105.763 41.222 ;
			RECT	106.067 41.158 106.099 41.222 ;
			RECT	106.403 41.158 106.435 41.222 ;
			RECT	106.739 41.158 106.771 41.222 ;
			RECT	107.075 41.158 107.107 41.222 ;
			RECT	107.411 41.158 107.443 41.222 ;
			RECT	107.747 41.158 107.779 41.222 ;
			RECT	108.083 41.158 108.115 41.222 ;
			RECT	108.419 41.158 108.451 41.222 ;
			RECT	108.755 41.158 108.787 41.222 ;
			RECT	109.091 41.158 109.123 41.222 ;
			RECT	109.427 41.158 109.459 41.222 ;
			RECT	109.763 41.158 109.795 41.222 ;
			RECT	110.099 41.158 110.131 41.222 ;
			RECT	110.435 41.158 110.467 41.222 ;
			RECT	110.771 41.158 110.803 41.222 ;
			RECT	111.107 41.158 111.139 41.222 ;
			RECT	111.443 41.158 111.475 41.222 ;
			RECT	111.779 41.158 111.811 41.222 ;
			RECT	112.115 41.158 112.147 41.222 ;
			RECT	112.451 41.158 112.483 41.222 ;
			RECT	112.787 41.158 112.819 41.222 ;
			RECT	113.123 41.158 113.155 41.222 ;
			RECT	113.459 41.158 113.491 41.222 ;
			RECT	113.795 41.158 113.827 41.222 ;
			RECT	114.131 41.158 114.163 41.222 ;
			RECT	114.467 41.158 114.499 41.222 ;
			RECT	114.803 41.158 114.835 41.222 ;
			RECT	115.139 41.158 115.171 41.222 ;
			RECT	115.475 41.158 115.507 41.222 ;
			RECT	115.811 41.158 115.843 41.222 ;
			RECT	116.147 41.158 116.179 41.222 ;
			RECT	116.483 41.158 116.515 41.222 ;
			RECT	116.819 41.158 116.851 41.222 ;
			RECT	117.155 41.158 117.187 41.222 ;
			RECT	117.491 41.158 117.523 41.222 ;
			RECT	117.827 41.158 117.859 41.222 ;
			RECT	118.163 41.158 118.195 41.222 ;
			RECT	118.499 41.158 118.531 41.222 ;
			RECT	118.835 41.158 118.867 41.222 ;
			RECT	119.171 41.158 119.203 41.222 ;
			RECT	119.507 41.158 119.539 41.222 ;
			RECT	119.843 41.158 119.875 41.222 ;
			RECT	120.179 41.158 120.211 41.222 ;
			RECT	120.515 41.158 120.547 41.222 ;
			RECT	120.851 41.158 120.883 41.222 ;
			RECT	121.187 41.158 121.219 41.222 ;
			RECT	121.523 41.158 121.555 41.222 ;
			RECT	121.859 41.158 121.891 41.222 ;
			RECT	122.195 41.158 122.227 41.222 ;
			RECT	122.531 41.158 122.563 41.222 ;
			RECT	122.867 41.158 122.899 41.222 ;
			RECT	123.203 41.158 123.235 41.222 ;
			RECT	123.539 41.158 123.571 41.222 ;
			RECT	123.875 41.158 123.907 41.222 ;
			RECT	124.211 41.158 124.243 41.222 ;
			RECT	124.547 41.158 124.579 41.222 ;
			RECT	124.883 41.158 124.915 41.222 ;
			RECT	125.219 41.158 125.251 41.222 ;
			RECT	125.555 41.158 125.587 41.222 ;
			RECT	126.222 41.158 126.254 41.222 ;
			RECT	126.894 41.158 126.926 41.222 ;
			RECT	127.566 41.158 127.598 41.222 ;
			RECT	128.238 41.158 128.27 41.222 ;
			RECT	128.91 41.158 128.942 41.222 ;
			RECT	129.246 41.158 129.278 41.222 ;
			RECT	129.582 41.158 129.614 41.222 ;
			RECT	130.254 41.158 130.286 41.222 ;
			RECT	130.59 41.158 130.622 41.222 ;
			RECT	130.926 41.158 130.958 41.222 ;
			RECT	131.598 41.158 131.63 41.222 ;
			RECT	131.934 41.158 131.966 41.222 ;
			RECT	132.942 41.158 132.974 41.222 ;
			RECT	133.278 41.158 133.31 41.222 ;
			RECT	134.286 41.158 134.318 41.222 ;
			RECT	134.622 41.158 134.654 41.222 ;
			RECT	135.63 41.158 135.662 41.222 ;
			RECT	135.966 41.158 135.998 41.222 ;
			RECT	136.302 41.158 136.334 41.222 ;
			RECT	136.974 41.158 137.006 41.222 ;
			RECT	137.31 41.158 137.342 41.222 ;
			RECT	137.646 41.158 137.678 41.222 ;
			RECT	137.982 41.158 138.014 41.222 ;
			RECT	138.654 41.158 138.686 41.222 ;
			RECT	138.99 41.158 139.022 41.222 ;
			RECT	139.662 41.158 139.694 41.222 ;
			RECT	139.998 41.158 140.03 41.222 ;
			RECT	140.334 41.158 140.366 41.222 ;
			RECT	141.006 41.158 141.038 41.222 ;
			RECT	141.342 41.158 141.374 41.222 ;
			RECT	142.35 41.158 142.382 41.222 ;
			RECT	143.022 41.158 143.054 41.222 ;
			RECT	143.694 41.158 143.726 41.222 ;
			RECT	144.366 41.158 144.398 41.222 ;
			RECT	145.038 41.158 145.07 41.222 ;
			RECT	145.374 41.158 145.406 41.222 ;
			RECT	146.382 41.158 146.414 41.222 ;
			RECT	146.842 41.158 146.874 41.222 ;
			RECT	147.636 41.158 147.668 41.222 ;
			RECT	148.415 41.158 148.479 41.222 ;
			RECT	149.272 41.158 149.304 41.222 ;
			RECT	149.792 41.158 149.824 41.222 ;
			RECT	150.595 41.158 150.627 41.222 ;
			RECT	151.401 41.158 151.433 41.222 ;
			RECT	153.202 41.158 153.266 41.222 ;
			RECT	154.142 41.158 154.174 41.222 ;
			RECT	154.662 41.158 154.694 41.222 ;
			RECT	155.505 41.158 155.569 41.222 ;
			RECT	155.748 41.158 155.812 41.222 ;
			RECT	156.532 41.158 156.564 41.222 ;
			RECT	157.326 41.158 157.358 41.222 ;
			RECT	157.786 41.158 157.818 41.222 ;
			RECT	158.794 41.158 158.826 41.222 ;
			RECT	159.13 41.158 159.162 41.222 ;
			RECT	159.802 41.158 159.834 41.222 ;
			RECT	160.474 41.158 160.506 41.222 ;
			RECT	161.146 41.158 161.178 41.222 ;
			RECT	161.818 41.158 161.85 41.222 ;
			RECT	162.826 41.158 162.858 41.222 ;
			RECT	163.162 41.158 163.194 41.222 ;
			RECT	163.834 41.158 163.866 41.222 ;
			RECT	164.17 41.158 164.202 41.222 ;
			RECT	164.506 41.158 164.538 41.222 ;
			RECT	165.178 41.158 165.21 41.222 ;
			RECT	165.514 41.158 165.546 41.222 ;
			RECT	166.186 41.158 166.218 41.222 ;
			RECT	166.522 41.158 166.554 41.222 ;
			RECT	166.858 41.158 166.89 41.222 ;
			RECT	167.194 41.158 167.226 41.222 ;
			RECT	167.866 41.158 167.898 41.222 ;
			RECT	168.202 41.158 168.234 41.222 ;
			RECT	168.538 41.158 168.57 41.222 ;
			RECT	169.546 41.158 169.578 41.222 ;
			RECT	169.882 41.158 169.914 41.222 ;
			RECT	170.89 41.158 170.922 41.222 ;
			RECT	171.226 41.158 171.258 41.222 ;
			RECT	172.234 41.158 172.266 41.222 ;
			RECT	172.57 41.158 172.602 41.222 ;
			RECT	173.242 41.158 173.274 41.222 ;
			RECT	173.578 41.158 173.61 41.222 ;
			RECT	173.914 41.158 173.946 41.222 ;
			RECT	174.586 41.158 174.618 41.222 ;
			RECT	174.922 41.158 174.954 41.222 ;
			RECT	175.258 41.158 175.29 41.222 ;
			RECT	175.93 41.158 175.962 41.222 ;
			RECT	176.602 41.158 176.634 41.222 ;
			RECT	177.274 41.158 177.306 41.222 ;
			RECT	177.946 41.158 177.978 41.222 ;
			RECT	178.613 41.158 178.645 41.222 ;
			RECT	178.949 41.158 178.981 41.222 ;
			RECT	179.285 41.158 179.317 41.222 ;
			RECT	179.621 41.158 179.653 41.222 ;
			RECT	179.957 41.158 179.989 41.222 ;
			RECT	180.293 41.158 180.325 41.222 ;
			RECT	180.629 41.158 180.661 41.222 ;
			RECT	180.965 41.158 180.997 41.222 ;
			RECT	181.301 41.158 181.333 41.222 ;
			RECT	181.637 41.158 181.669 41.222 ;
			RECT	181.973 41.158 182.005 41.222 ;
			RECT	182.309 41.158 182.341 41.222 ;
			RECT	182.645 41.158 182.677 41.222 ;
			RECT	182.981 41.158 183.013 41.222 ;
			RECT	183.317 41.158 183.349 41.222 ;
			RECT	183.653 41.158 183.685 41.222 ;
			RECT	183.989 41.158 184.021 41.222 ;
			RECT	184.325 41.158 184.357 41.222 ;
			RECT	184.661 41.158 184.693 41.222 ;
			RECT	184.997 41.158 185.029 41.222 ;
			RECT	185.333 41.158 185.365 41.222 ;
			RECT	185.669 41.158 185.701 41.222 ;
			RECT	186.005 41.158 186.037 41.222 ;
			RECT	186.341 41.158 186.373 41.222 ;
			RECT	186.677 41.158 186.709 41.222 ;
			RECT	187.013 41.158 187.045 41.222 ;
			RECT	187.349 41.158 187.381 41.222 ;
			RECT	187.685 41.158 187.717 41.222 ;
			RECT	188.021 41.158 188.053 41.222 ;
			RECT	188.357 41.158 188.389 41.222 ;
			RECT	188.693 41.158 188.725 41.222 ;
			RECT	189.029 41.158 189.061 41.222 ;
			RECT	189.365 41.158 189.397 41.222 ;
			RECT	189.701 41.158 189.733 41.222 ;
			RECT	190.037 41.158 190.069 41.222 ;
			RECT	190.373 41.158 190.405 41.222 ;
			RECT	190.709 41.158 190.741 41.222 ;
			RECT	191.045 41.158 191.077 41.222 ;
			RECT	191.381 41.158 191.413 41.222 ;
			RECT	191.717 41.158 191.749 41.222 ;
			RECT	192.053 41.158 192.085 41.222 ;
			RECT	192.389 41.158 192.421 41.222 ;
			RECT	192.725 41.158 192.757 41.222 ;
			RECT	193.061 41.158 193.093 41.222 ;
			RECT	193.397 41.158 193.429 41.222 ;
			RECT	193.733 41.158 193.765 41.222 ;
			RECT	194.069 41.158 194.101 41.222 ;
			RECT	194.405 41.158 194.437 41.222 ;
			RECT	194.741 41.158 194.773 41.222 ;
			RECT	195.077 41.158 195.109 41.222 ;
			RECT	195.413 41.158 195.445 41.222 ;
			RECT	195.749 41.158 195.781 41.222 ;
			RECT	196.085 41.158 196.117 41.222 ;
			RECT	196.421 41.158 196.453 41.222 ;
			RECT	196.757 41.158 196.789 41.222 ;
			RECT	197.093 41.158 197.125 41.222 ;
			RECT	197.429 41.158 197.461 41.222 ;
			RECT	197.765 41.158 197.797 41.222 ;
			RECT	198.101 41.158 198.133 41.222 ;
			RECT	198.437 41.158 198.469 41.222 ;
			RECT	198.773 41.158 198.805 41.222 ;
			RECT	199.109 41.158 199.141 41.222 ;
			RECT	199.445 41.158 199.477 41.222 ;
			RECT	199.781 41.158 199.813 41.222 ;
			RECT	201.307 41.158 201.339 41.222 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 43.241 201.665 43.331 ;
			LAYER	J3 ;
			RECT	0.781 43.254 0.813 43.318 ;
			RECT	1.024 43.254 1.056 43.318 ;
			RECT	1.838 43.254 1.87 43.318 ;
			RECT	2.517 43.254 2.549 43.318 ;
			RECT	3.922 43.254 3.954 43.318 ;
			RECT	4.136 43.254 4.168 43.318 ;
			RECT	4.258 43.254 4.29 43.318 ;
			RECT	4.51 43.254 4.542 43.318 ;
			RECT	5.164 43.254 5.196 43.318 ;
			RECT	28.224 43.254 28.256 43.318 ;
			RECT	28.896 43.254 28.928 43.318 ;
			RECT	31.248 43.254 31.28 43.318 ;
			RECT	32.256 43.254 32.288 43.318 ;
			RECT	32.928 43.254 32.96 43.318 ;
			RECT	33.6 43.254 33.632 43.318 ;
			RECT	33.936 43.254 33.968 43.318 ;
			RECT	34.944 43.254 34.976 43.318 ;
			RECT	36.624 43.254 36.656 43.318 ;
			RECT	38.976 43.254 39.008 43.318 ;
			RECT	39.648 43.254 39.68 43.318 ;
			RECT	40.992 43.254 41.024 43.318 ;
			RECT	42 43.254 42.032 43.318 ;
			RECT	42.336 43.254 42.368 43.318 ;
			RECT	43.008 43.254 43.04 43.318 ;
			RECT	43.344 43.254 43.376 43.318 ;
			RECT	44.352 43.254 44.384 43.318 ;
			RECT	45.024 43.254 45.056 43.318 ;
			RECT	46.368 43.254 46.4 43.318 ;
			RECT	48.844 43.254 48.876 43.318 ;
			RECT	50.433 43.254 50.465 43.318 ;
			RECT	51.275 43.254 51.307 43.318 ;
			RECT	51.794 43.254 51.826 43.318 ;
			RECT	52.597 43.254 52.629 43.318 ;
			RECT	53.403 43.254 53.435 43.318 ;
			RECT	54.117 43.254 54.149 43.318 ;
			RECT	55.22 43.254 55.252 43.318 ;
			RECT	56.144 43.256 56.176 43.32 ;
			RECT	56.664 43.257 56.696 43.321 ;
			RECT	57.507 43.27 57.571 43.302 ;
			RECT	57.766 43.254 57.798 43.318 ;
			RECT	59.328 43.254 59.36 43.318 ;
			RECT	61.804 43.254 61.836 43.318 ;
			RECT	63.148 43.254 63.18 43.318 ;
			RECT	63.82 43.254 63.852 43.318 ;
			RECT	64.828 43.254 64.86 43.318 ;
			RECT	65.164 43.254 65.196 43.318 ;
			RECT	65.836 43.254 65.868 43.318 ;
			RECT	66.172 43.254 66.204 43.318 ;
			RECT	67.18 43.254 67.212 43.318 ;
			RECT	68.524 43.254 68.556 43.318 ;
			RECT	69.196 43.254 69.228 43.318 ;
			RECT	71.548 43.254 71.58 43.318 ;
			RECT	73.228 43.254 73.26 43.318 ;
			RECT	74.236 43.254 74.268 43.318 ;
			RECT	74.572 43.254 74.604 43.318 ;
			RECT	75.244 43.254 75.276 43.318 ;
			RECT	75.916 43.254 75.948 43.318 ;
			RECT	76.924 43.254 76.956 43.318 ;
			RECT	79.276 43.254 79.308 43.318 ;
			RECT	79.948 43.254 79.98 43.318 ;
			RECT	126.222 43.254 126.254 43.318 ;
			RECT	126.894 43.254 126.926 43.318 ;
			RECT	129.246 43.254 129.278 43.318 ;
			RECT	130.254 43.254 130.286 43.318 ;
			RECT	130.926 43.254 130.958 43.318 ;
			RECT	131.598 43.254 131.63 43.318 ;
			RECT	131.934 43.254 131.966 43.318 ;
			RECT	132.942 43.254 132.974 43.318 ;
			RECT	134.622 43.254 134.654 43.318 ;
			RECT	136.974 43.254 137.006 43.318 ;
			RECT	137.646 43.254 137.678 43.318 ;
			RECT	138.99 43.254 139.022 43.318 ;
			RECT	139.998 43.254 140.03 43.318 ;
			RECT	140.334 43.254 140.366 43.318 ;
			RECT	141.006 43.254 141.038 43.318 ;
			RECT	141.342 43.254 141.374 43.318 ;
			RECT	142.35 43.254 142.382 43.318 ;
			RECT	143.022 43.254 143.054 43.318 ;
			RECT	144.366 43.254 144.398 43.318 ;
			RECT	146.842 43.254 146.874 43.318 ;
			RECT	148.431 43.254 148.463 43.318 ;
			RECT	149.273 43.254 149.305 43.318 ;
			RECT	149.792 43.254 149.824 43.318 ;
			RECT	150.595 43.254 150.627 43.318 ;
			RECT	151.401 43.254 151.433 43.318 ;
			RECT	152.115 43.254 152.147 43.318 ;
			RECT	153.218 43.254 153.25 43.318 ;
			RECT	154.142 43.256 154.174 43.32 ;
			RECT	154.662 43.257 154.694 43.321 ;
			RECT	155.505 43.27 155.569 43.302 ;
			RECT	155.764 43.254 155.796 43.318 ;
			RECT	157.326 43.254 157.358 43.318 ;
			RECT	159.802 43.254 159.834 43.318 ;
			RECT	161.146 43.254 161.178 43.318 ;
			RECT	161.818 43.254 161.85 43.318 ;
			RECT	162.826 43.254 162.858 43.318 ;
			RECT	163.162 43.254 163.194 43.318 ;
			RECT	163.834 43.254 163.866 43.318 ;
			RECT	164.17 43.254 164.202 43.318 ;
			RECT	165.178 43.254 165.21 43.318 ;
			RECT	166.522 43.254 166.554 43.318 ;
			RECT	167.194 43.254 167.226 43.318 ;
			RECT	169.546 43.254 169.578 43.318 ;
			RECT	171.226 43.254 171.258 43.318 ;
			RECT	172.234 43.254 172.266 43.318 ;
			RECT	172.57 43.254 172.602 43.318 ;
			RECT	173.242 43.254 173.274 43.318 ;
			RECT	173.914 43.254 173.946 43.318 ;
			RECT	174.922 43.254 174.954 43.318 ;
			RECT	177.274 43.254 177.306 43.318 ;
			RECT	177.946 43.254 177.978 43.318 ;
			RECT	201.307 43.254 201.339 43.318 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 44.585 201.665 44.675 ;
			LAYER	J3 ;
			RECT	1.024 44.598 1.056 44.662 ;
			RECT	1.838 44.598 1.87 44.662 ;
			RECT	2.517 44.598 2.549 44.662 ;
			RECT	3.313 44.598 3.345 44.662 ;
			RECT	3.719 44.598 3.751 44.662 ;
			RECT	3.922 44.598 3.954 44.662 ;
			RECT	4.138 44.598 4.17 44.662 ;
			RECT	4.419 44.598 4.451 44.662 ;
			RECT	5.164 44.598 5.196 44.662 ;
			RECT	28.224 44.598 28.256 44.662 ;
			RECT	28.896 44.598 28.928 44.662 ;
			RECT	31.248 44.598 31.28 44.662 ;
			RECT	32.256 44.598 32.288 44.662 ;
			RECT	34.944 44.598 34.976 44.662 ;
			RECT	36.284 44.598 36.316 44.662 ;
			RECT	36.624 44.598 36.656 44.662 ;
			RECT	38.976 44.598 39.008 44.662 ;
			RECT	40.992 44.598 41.024 44.662 ;
			RECT	42 44.598 42.032 44.662 ;
			RECT	42.336 44.598 42.368 44.662 ;
			RECT	43.008 44.598 43.04 44.662 ;
			RECT	43.344 44.598 43.376 44.662 ;
			RECT	44.352 44.598 44.384 44.662 ;
			RECT	46.368 44.598 46.4 44.662 ;
			RECT	48.844 44.598 48.876 44.662 ;
			RECT	50.433 44.598 50.465 44.662 ;
			RECT	51.275 44.598 51.307 44.662 ;
			RECT	51.794 44.598 51.826 44.662 ;
			RECT	52.597 44.598 52.629 44.662 ;
			RECT	53.403 44.598 53.435 44.662 ;
			RECT	56.144 44.596 56.176 44.66 ;
			RECT	56.664 44.597 56.696 44.661 ;
			RECT	57.507 44.614 57.571 44.646 ;
			RECT	59.328 44.598 59.36 44.662 ;
			RECT	61.804 44.598 61.836 44.662 ;
			RECT	63.82 44.598 63.852 44.662 ;
			RECT	64.828 44.598 64.86 44.662 ;
			RECT	65.164 44.598 65.196 44.662 ;
			RECT	65.836 44.598 65.868 44.662 ;
			RECT	66.172 44.598 66.204 44.662 ;
			RECT	67.18 44.598 67.212 44.662 ;
			RECT	69.196 44.598 69.228 44.662 ;
			RECT	71.548 44.598 71.58 44.662 ;
			RECT	71.888 44.598 71.92 44.662 ;
			RECT	73.228 44.598 73.26 44.662 ;
			RECT	75.916 44.598 75.948 44.662 ;
			RECT	76.924 44.598 76.956 44.662 ;
			RECT	79.276 44.598 79.308 44.662 ;
			RECT	79.948 44.598 79.98 44.662 ;
			RECT	126.222 44.598 126.254 44.662 ;
			RECT	126.894 44.598 126.926 44.662 ;
			RECT	129.246 44.598 129.278 44.662 ;
			RECT	130.254 44.598 130.286 44.662 ;
			RECT	132.942 44.598 132.974 44.662 ;
			RECT	134.282 44.598 134.314 44.662 ;
			RECT	134.622 44.598 134.654 44.662 ;
			RECT	136.974 44.598 137.006 44.662 ;
			RECT	138.99 44.598 139.022 44.662 ;
			RECT	139.998 44.598 140.03 44.662 ;
			RECT	140.334 44.598 140.366 44.662 ;
			RECT	141.006 44.598 141.038 44.662 ;
			RECT	141.342 44.598 141.374 44.662 ;
			RECT	142.35 44.598 142.382 44.662 ;
			RECT	144.366 44.598 144.398 44.662 ;
			RECT	146.842 44.598 146.874 44.662 ;
			RECT	148.431 44.598 148.463 44.662 ;
			RECT	149.273 44.598 149.305 44.662 ;
			RECT	149.792 44.598 149.824 44.662 ;
			RECT	150.595 44.598 150.627 44.662 ;
			RECT	151.401 44.598 151.433 44.662 ;
			RECT	154.142 44.596 154.174 44.66 ;
			RECT	154.662 44.597 154.694 44.661 ;
			RECT	155.505 44.614 155.569 44.646 ;
			RECT	157.326 44.598 157.358 44.662 ;
			RECT	159.802 44.598 159.834 44.662 ;
			RECT	161.818 44.598 161.85 44.662 ;
			RECT	162.826 44.598 162.858 44.662 ;
			RECT	163.162 44.598 163.194 44.662 ;
			RECT	163.834 44.598 163.866 44.662 ;
			RECT	164.17 44.598 164.202 44.662 ;
			RECT	165.178 44.598 165.21 44.662 ;
			RECT	167.194 44.598 167.226 44.662 ;
			RECT	169.546 44.598 169.578 44.662 ;
			RECT	169.886 44.598 169.918 44.662 ;
			RECT	171.226 44.598 171.258 44.662 ;
			RECT	173.914 44.598 173.946 44.662 ;
			RECT	174.922 44.598 174.954 44.662 ;
			RECT	177.274 44.598 177.306 44.662 ;
			RECT	177.946 44.598 177.978 44.662 ;
			RECT	201.307 44.593 201.339 44.657 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 45.628 201.665 45.748 ;
			LAYER	J3 ;
			RECT	1.024 45.656 1.056 45.72 ;
			RECT	1.822 45.656 1.886 45.72 ;
			RECT	2.501 45.656 2.565 45.72 ;
			RECT	3.719 45.656 3.751 45.72 ;
			RECT	3.922 45.656 3.954 45.72 ;
			RECT	4.138 45.656 4.17 45.72 ;
			RECT	4.419 45.656 4.451 45.72 ;
			RECT	5.164 45.656 5.196 45.72 ;
			RECT	50.417 45.656 50.481 45.72 ;
			RECT	51.275 45.656 51.307 45.72 ;
			RECT	51.794 45.656 51.826 45.72 ;
			RECT	52.597 45.656 52.629 45.72 ;
			RECT	54.657 45.656 54.689 45.72 ;
			RECT	55.21 45.656 55.274 45.72 ;
			RECT	56.144 45.656 56.176 45.72 ;
			RECT	56.664 45.656 56.696 45.72 ;
			RECT	57.278 45.656 57.31 45.72 ;
			RECT	57.507 45.656 57.571 45.72 ;
			RECT	148.415 45.656 148.479 45.72 ;
			RECT	149.273 45.656 149.305 45.72 ;
			RECT	149.792 45.656 149.824 45.72 ;
			RECT	150.595 45.656 150.627 45.72 ;
			RECT	152.655 45.656 152.687 45.72 ;
			RECT	153.208 45.656 153.272 45.72 ;
			RECT	154.142 45.656 154.174 45.72 ;
			RECT	154.662 45.656 154.694 45.72 ;
			RECT	155.276 45.656 155.308 45.72 ;
			RECT	155.505 45.656 155.569 45.72 ;
			RECT	201.307 45.656 201.339 45.72 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 46.363 201.665 46.453 ;
			LAYER	J3 ;
			RECT	1.024 46.376 1.056 46.44 ;
			RECT	1.822 46.392 1.886 46.424 ;
			RECT	2.517 46.376 2.549 46.44 ;
			RECT	3.719 46.376 3.751 46.44 ;
			RECT	3.922 46.376 3.954 46.44 ;
			RECT	4.138 46.376 4.17 46.44 ;
			RECT	4.281 46.376 4.313 46.44 ;
			RECT	4.422 46.376 4.454 46.44 ;
			RECT	48.845 46.376 48.877 46.44 ;
			RECT	50.433 46.376 50.465 46.44 ;
			RECT	51.274 46.376 51.306 46.44 ;
			RECT	51.791 46.375 51.823 46.439 ;
			RECT	52.597 46.376 52.629 46.44 ;
			RECT	53.403 46.376 53.435 46.44 ;
			RECT	54.657 46.376 54.689 46.44 ;
			RECT	55.24 46.376 55.272 46.44 ;
			RECT	56.144 46.375 56.176 46.439 ;
			RECT	56.664 46.376 56.696 46.44 ;
			RECT	57.278 46.376 57.31 46.44 ;
			RECT	57.507 46.392 57.571 46.424 ;
			RECT	59.327 46.376 59.359 46.44 ;
			RECT	146.843 46.376 146.875 46.44 ;
			RECT	148.431 46.376 148.463 46.44 ;
			RECT	149.272 46.376 149.304 46.44 ;
			RECT	149.789 46.375 149.821 46.439 ;
			RECT	150.595 46.376 150.627 46.44 ;
			RECT	151.401 46.376 151.433 46.44 ;
			RECT	152.655 46.376 152.687 46.44 ;
			RECT	153.238 46.376 153.27 46.44 ;
			RECT	154.142 46.375 154.174 46.439 ;
			RECT	154.662 46.376 154.694 46.44 ;
			RECT	155.276 46.376 155.308 46.44 ;
			RECT	155.505 46.392 155.569 46.424 ;
			RECT	157.325 46.376 157.357 46.44 ;
			RECT	201.307 46.376 201.339 46.44 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 47.153 201.665 47.273 ;
			LAYER	J3 ;
			RECT	1.024 47.181 1.056 47.245 ;
			RECT	1.822 47.181 1.886 47.245 ;
			RECT	2.501 47.181 2.565 47.245 ;
			RECT	3.318 47.181 3.35 47.245 ;
			RECT	3.719 47.181 3.751 47.245 ;
			RECT	3.922 47.181 3.954 47.245 ;
			RECT	4.138 47.181 4.17 47.245 ;
			RECT	4.281 47.181 4.313 47.245 ;
			RECT	5.164 47.181 5.196 47.245 ;
			RECT	48.845 47.181 48.877 47.245 ;
			RECT	52.597 47.181 52.629 47.245 ;
			RECT	53.403 47.181 53.435 47.245 ;
			RECT	55.21 47.181 55.274 47.245 ;
			RECT	57.278 47.181 57.31 47.245 ;
			RECT	59.327 47.181 59.359 47.245 ;
			RECT	146.843 47.181 146.875 47.245 ;
			RECT	150.595 47.181 150.627 47.245 ;
			RECT	151.401 47.181 151.433 47.245 ;
			RECT	153.208 47.181 153.272 47.245 ;
			RECT	155.276 47.181 155.308 47.245 ;
			RECT	157.325 47.181 157.357 47.245 ;
			RECT	201.004 47.181 201.036 47.245 ;
			RECT	201.307 47.181 201.339 47.245 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 47.798 201.665 47.918 ;
			LAYER	J3 ;
			RECT	1.024 47.826 1.056 47.89 ;
			RECT	1.822 47.826 1.886 47.89 ;
			RECT	2.501 47.826 2.565 47.89 ;
			RECT	3.719 47.826 3.751 47.89 ;
			RECT	3.922 47.826 3.954 47.89 ;
			RECT	4.281 47.826 4.313 47.89 ;
			RECT	5.164 47.826 5.196 47.89 ;
			RECT	52.597 47.826 52.629 47.89 ;
			RECT	53.403 47.842 53.435 47.874 ;
			RECT	55.21 47.826 55.274 47.89 ;
			RECT	57.278 47.826 57.31 47.89 ;
			RECT	150.595 47.826 150.627 47.89 ;
			RECT	151.401 47.842 151.433 47.874 ;
			RECT	153.208 47.826 153.272 47.89 ;
			RECT	155.276 47.826 155.308 47.89 ;
			RECT	201.307 47.826 201.339 47.89 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 42.086 201.665 42.176 ;
			LAYER	J3 ;
			RECT	1.822 42.115 1.886 42.147 ;
			RECT	2.501 42.115 2.565 42.147 ;
			RECT	2.988 42.099 3.02 42.163 ;
			RECT	4.51 42.099 4.542 42.163 ;
			RECT	5.164 42.115 5.196 42.147 ;
			RECT	28.224 42.099 28.256 42.163 ;
			RECT	28.896 42.099 28.928 42.163 ;
			RECT	31.248 42.099 31.28 42.163 ;
			RECT	32.256 42.099 32.288 42.163 ;
			RECT	32.928 42.099 32.96 42.163 ;
			RECT	33.6 42.099 33.632 42.163 ;
			RECT	33.936 42.099 33.968 42.163 ;
			RECT	34.944 42.099 34.976 42.163 ;
			RECT	36.624 42.099 36.656 42.163 ;
			RECT	38.976 42.099 39.008 42.163 ;
			RECT	39.648 42.099 39.68 42.163 ;
			RECT	40.992 42.099 41.024 42.163 ;
			RECT	42 42.099 42.032 42.163 ;
			RECT	42.336 42.099 42.368 42.163 ;
			RECT	43.008 42.099 43.04 42.163 ;
			RECT	43.344 42.099 43.376 42.163 ;
			RECT	44.352 42.099 44.384 42.163 ;
			RECT	45.024 42.099 45.056 42.163 ;
			RECT	46.368 42.099 46.4 42.163 ;
			RECT	49.531 42.099 49.563 42.163 ;
			RECT	51.274 42.099 51.306 42.163 ;
			RECT	51.794 42.099 51.826 42.163 ;
			RECT	52.597 42.099 52.629 42.163 ;
			RECT	53.406 42.099 53.438 42.163 ;
			RECT	55.204 42.115 55.268 42.147 ;
			RECT	56.144 42.099 56.176 42.163 ;
			RECT	56.664 42.099 56.696 42.163 ;
			RECT	57.507 42.115 57.571 42.147 ;
			RECT	58.641 42.099 58.673 42.163 ;
			RECT	61.804 42.099 61.836 42.163 ;
			RECT	63.148 42.099 63.18 42.163 ;
			RECT	63.82 42.099 63.852 42.163 ;
			RECT	64.828 42.099 64.86 42.163 ;
			RECT	65.164 42.099 65.196 42.163 ;
			RECT	65.836 42.099 65.868 42.163 ;
			RECT	66.172 42.099 66.204 42.163 ;
			RECT	67.18 42.099 67.212 42.163 ;
			RECT	68.524 42.099 68.556 42.163 ;
			RECT	69.196 42.099 69.228 42.163 ;
			RECT	71.548 42.099 71.58 42.163 ;
			RECT	73.228 42.099 73.26 42.163 ;
			RECT	74.236 42.099 74.268 42.163 ;
			RECT	74.572 42.099 74.604 42.163 ;
			RECT	75.244 42.099 75.276 42.163 ;
			RECT	75.916 42.099 75.948 42.163 ;
			RECT	76.924 42.099 76.956 42.163 ;
			RECT	79.276 42.099 79.308 42.163 ;
			RECT	79.948 42.099 79.98 42.163 ;
			RECT	126.222 42.099 126.254 42.163 ;
			RECT	126.894 42.099 126.926 42.163 ;
			RECT	129.246 42.099 129.278 42.163 ;
			RECT	130.254 42.099 130.286 42.163 ;
			RECT	130.926 42.099 130.958 42.163 ;
			RECT	131.598 42.099 131.63 42.163 ;
			RECT	131.934 42.099 131.966 42.163 ;
			RECT	132.942 42.099 132.974 42.163 ;
			RECT	134.622 42.099 134.654 42.163 ;
			RECT	136.974 42.099 137.006 42.163 ;
			RECT	137.646 42.099 137.678 42.163 ;
			RECT	138.99 42.099 139.022 42.163 ;
			RECT	139.998 42.099 140.03 42.163 ;
			RECT	140.334 42.099 140.366 42.163 ;
			RECT	141.006 42.099 141.038 42.163 ;
			RECT	141.342 42.099 141.374 42.163 ;
			RECT	142.35 42.099 142.382 42.163 ;
			RECT	143.022 42.099 143.054 42.163 ;
			RECT	144.366 42.099 144.398 42.163 ;
			RECT	147.529 42.099 147.561 42.163 ;
			RECT	149.272 42.099 149.304 42.163 ;
			RECT	149.792 42.099 149.824 42.163 ;
			RECT	150.595 42.099 150.627 42.163 ;
			RECT	151.404 42.099 151.436 42.163 ;
			RECT	153.202 42.115 153.266 42.147 ;
			RECT	154.142 42.099 154.174 42.163 ;
			RECT	154.662 42.099 154.694 42.163 ;
			RECT	155.505 42.115 155.569 42.147 ;
			RECT	156.639 42.099 156.671 42.163 ;
			RECT	159.802 42.099 159.834 42.163 ;
			RECT	161.146 42.099 161.178 42.163 ;
			RECT	161.818 42.099 161.85 42.163 ;
			RECT	162.826 42.099 162.858 42.163 ;
			RECT	163.162 42.099 163.194 42.163 ;
			RECT	163.834 42.099 163.866 42.163 ;
			RECT	164.17 42.099 164.202 42.163 ;
			RECT	165.178 42.099 165.21 42.163 ;
			RECT	166.522 42.099 166.554 42.163 ;
			RECT	167.194 42.099 167.226 42.163 ;
			RECT	169.546 42.099 169.578 42.163 ;
			RECT	171.226 42.099 171.258 42.163 ;
			RECT	172.234 42.099 172.266 42.163 ;
			RECT	172.57 42.099 172.602 42.163 ;
			RECT	173.242 42.099 173.274 42.163 ;
			RECT	173.914 42.099 173.946 42.163 ;
			RECT	174.922 42.099 174.954 42.163 ;
			RECT	177.274 42.099 177.306 42.163 ;
			RECT	177.946 42.099 177.978 42.163 ;
			RECT	201.307 42.099 201.339 42.163 ;
		END

	END VDDPE

	PIN VSSE
		USE GROUND ;
		DIRECTION INOUT ;
		PORT
			LAYER	C4 ;
			RECT	0.294 81.843 201.665 81.933 ;
			LAYER	J3 ;
			RECT	0.908 81.856 0.94 81.92 ;
			RECT	5.927 81.856 5.959 81.92 ;
			RECT	6.095 81.856 6.127 81.92 ;
			RECT	49.271 81.856 49.303 81.92 ;
			RECT	49.439 81.856 49.471 81.92 ;
			RECT	51.881 81.856 51.913 81.92 ;
			RECT	53.534 81.872 53.598 81.904 ;
			RECT	58.733 81.856 58.765 81.92 ;
			RECT	58.901 81.856 58.933 81.92 ;
			RECT	102.077 81.856 102.109 81.92 ;
			RECT	102.245 81.856 102.277 81.92 ;
			RECT	103.925 81.856 103.957 81.92 ;
			RECT	104.093 81.856 104.125 81.92 ;
			RECT	147.269 81.856 147.301 81.92 ;
			RECT	147.437 81.856 147.469 81.92 ;
			RECT	149.879 81.856 149.911 81.92 ;
			RECT	151.532 81.872 151.596 81.904 ;
			RECT	156.731 81.856 156.763 81.92 ;
			RECT	156.899 81.856 156.931 81.92 ;
			RECT	200.075 81.856 200.107 81.92 ;
			RECT	200.243 81.856 200.275 81.92 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 0.243 201.665 0.333 ;
			LAYER	J3 ;
			RECT	0.908 0.256 0.94 0.32 ;
			RECT	5.927 0.256 5.959 0.32 ;
			RECT	6.095 0.256 6.127 0.32 ;
			RECT	49.271 0.256 49.303 0.32 ;
			RECT	49.439 0.256 49.471 0.32 ;
			RECT	51.881 0.256 51.913 0.32 ;
			RECT	53.534 0.272 53.598 0.304 ;
			RECT	58.733 0.256 58.765 0.32 ;
			RECT	58.901 0.256 58.933 0.32 ;
			RECT	102.077 0.256 102.109 0.32 ;
			RECT	102.245 0.256 102.277 0.32 ;
			RECT	103.925 0.256 103.957 0.32 ;
			RECT	104.093 0.256 104.125 0.32 ;
			RECT	147.269 0.256 147.301 0.32 ;
			RECT	147.437 0.256 147.469 0.32 ;
			RECT	149.879 0.256 149.911 0.32 ;
			RECT	151.532 0.272 151.596 0.304 ;
			RECT	156.731 0.256 156.763 0.32 ;
			RECT	156.899 0.256 156.931 0.32 ;
			RECT	200.075 0.256 200.107 0.32 ;
			RECT	200.243 0.256 200.275 0.32 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 31.538 201.665 31.648 ;
			LAYER	J3 ;
			RECT	0.755 31.561 0.787 31.625 ;
			RECT	1.645 31.561 1.709 31.625 ;
			RECT	2.323 31.577 2.387 31.609 ;
			RECT	3.438 31.561 3.47 31.625 ;
			RECT	3.585 31.561 3.617 31.625 ;
			RECT	3.755 31.561 3.787 31.625 ;
			RECT	4.195 31.561 4.227 31.625 ;
			RECT	4.944 31.561 5.008 31.625 ;
			RECT	5.409 31.561 5.441 31.625 ;
			RECT	49.311 31.561 49.375 31.625 ;
			RECT	52.124 31.561 52.156 31.625 ;
			RECT	52.578 31.561 52.61 31.625 ;
			RECT	53.132 31.561 53.196 31.625 ;
			RECT	53.91 31.561 53.942 31.625 ;
			RECT	54.251 31.561 54.283 31.625 ;
			RECT	55.562 31.561 55.626 31.625 ;
			RECT	55.803 31.561 55.835 31.625 ;
			RECT	58.829 31.561 58.893 31.625 ;
			RECT	102.763 31.561 102.795 31.625 ;
			RECT	102.995 31.561 103.027 31.625 ;
			RECT	103.175 31.561 103.207 31.625 ;
			RECT	103.407 31.561 103.439 31.625 ;
			RECT	147.309 31.561 147.373 31.625 ;
			RECT	150.122 31.561 150.154 31.625 ;
			RECT	150.576 31.561 150.608 31.625 ;
			RECT	151.13 31.561 151.194 31.625 ;
			RECT	151.908 31.561 151.94 31.625 ;
			RECT	152.249 31.561 152.281 31.625 ;
			RECT	153.56 31.561 153.624 31.625 ;
			RECT	153.801 31.561 153.833 31.625 ;
			RECT	156.827 31.561 156.891 31.625 ;
			RECT	200.761 31.561 200.793 31.625 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 32.248 201.665 32.358 ;
			LAYER	J3 ;
			RECT	1.645 32.271 1.709 32.335 ;
			RECT	2.129 32.271 2.161 32.335 ;
			RECT	2.323 32.271 2.387 32.335 ;
			RECT	3.438 32.271 3.47 32.335 ;
			RECT	3.755 32.271 3.787 32.335 ;
			RECT	4.195 32.271 4.227 32.335 ;
			RECT	4.944 32.271 5.008 32.335 ;
			RECT	6.347 32.271 6.379 32.335 ;
			RECT	6.683 32.271 6.715 32.335 ;
			RECT	7.019 32.271 7.051 32.335 ;
			RECT	7.355 32.271 7.387 32.335 ;
			RECT	7.691 32.271 7.723 32.335 ;
			RECT	8.027 32.271 8.059 32.335 ;
			RECT	8.363 32.271 8.395 32.335 ;
			RECT	8.699 32.271 8.731 32.335 ;
			RECT	9.035 32.271 9.067 32.335 ;
			RECT	9.371 32.271 9.403 32.335 ;
			RECT	9.707 32.271 9.739 32.335 ;
			RECT	10.043 32.271 10.075 32.335 ;
			RECT	10.379 32.271 10.411 32.335 ;
			RECT	10.715 32.271 10.747 32.335 ;
			RECT	11.051 32.271 11.083 32.335 ;
			RECT	11.387 32.271 11.419 32.335 ;
			RECT	11.723 32.271 11.755 32.335 ;
			RECT	12.059 32.271 12.091 32.335 ;
			RECT	12.395 32.271 12.427 32.335 ;
			RECT	12.731 32.271 12.763 32.335 ;
			RECT	13.067 32.271 13.099 32.335 ;
			RECT	13.403 32.271 13.435 32.335 ;
			RECT	13.739 32.271 13.771 32.335 ;
			RECT	14.075 32.271 14.107 32.335 ;
			RECT	14.411 32.271 14.443 32.335 ;
			RECT	14.747 32.271 14.779 32.335 ;
			RECT	15.083 32.271 15.115 32.335 ;
			RECT	15.419 32.271 15.451 32.335 ;
			RECT	15.755 32.271 15.787 32.335 ;
			RECT	16.091 32.271 16.123 32.335 ;
			RECT	16.427 32.271 16.459 32.335 ;
			RECT	16.763 32.271 16.795 32.335 ;
			RECT	17.099 32.271 17.131 32.335 ;
			RECT	17.435 32.271 17.467 32.335 ;
			RECT	17.771 32.271 17.803 32.335 ;
			RECT	18.107 32.271 18.139 32.335 ;
			RECT	18.443 32.271 18.475 32.335 ;
			RECT	18.779 32.271 18.811 32.335 ;
			RECT	19.115 32.271 19.147 32.335 ;
			RECT	19.451 32.271 19.483 32.335 ;
			RECT	19.787 32.271 19.819 32.335 ;
			RECT	20.123 32.271 20.155 32.335 ;
			RECT	20.459 32.271 20.491 32.335 ;
			RECT	20.795 32.271 20.827 32.335 ;
			RECT	21.131 32.271 21.163 32.335 ;
			RECT	21.467 32.271 21.499 32.335 ;
			RECT	21.803 32.271 21.835 32.335 ;
			RECT	22.139 32.271 22.171 32.335 ;
			RECT	22.475 32.271 22.507 32.335 ;
			RECT	22.811 32.271 22.843 32.335 ;
			RECT	23.147 32.271 23.179 32.335 ;
			RECT	23.483 32.271 23.515 32.335 ;
			RECT	23.819 32.271 23.851 32.335 ;
			RECT	24.155 32.271 24.187 32.335 ;
			RECT	24.491 32.271 24.523 32.335 ;
			RECT	24.827 32.271 24.859 32.335 ;
			RECT	25.163 32.271 25.195 32.335 ;
			RECT	25.499 32.271 25.531 32.335 ;
			RECT	25.835 32.271 25.867 32.335 ;
			RECT	26.171 32.271 26.203 32.335 ;
			RECT	26.507 32.271 26.539 32.335 ;
			RECT	26.843 32.271 26.875 32.335 ;
			RECT	27.179 32.271 27.211 32.335 ;
			RECT	27.515 32.271 27.547 32.335 ;
			RECT	49.311 32.271 49.375 32.335 ;
			RECT	52.124 32.271 52.156 32.335 ;
			RECT	52.578 32.271 52.61 32.335 ;
			RECT	52.968 32.271 53.032 32.335 ;
			RECT	54.251 32.271 54.283 32.335 ;
			RECT	55.562 32.271 55.626 32.335 ;
			RECT	55.803 32.271 55.835 32.335 ;
			RECT	58.829 32.271 58.893 32.335 ;
			RECT	80.657 32.271 80.689 32.335 ;
			RECT	80.993 32.271 81.025 32.335 ;
			RECT	81.329 32.271 81.361 32.335 ;
			RECT	81.665 32.271 81.697 32.335 ;
			RECT	82.001 32.271 82.033 32.335 ;
			RECT	82.337 32.271 82.369 32.335 ;
			RECT	82.673 32.271 82.705 32.335 ;
			RECT	83.009 32.271 83.041 32.335 ;
			RECT	83.345 32.271 83.377 32.335 ;
			RECT	83.681 32.271 83.713 32.335 ;
			RECT	84.017 32.271 84.049 32.335 ;
			RECT	84.353 32.271 84.385 32.335 ;
			RECT	84.689 32.271 84.721 32.335 ;
			RECT	85.025 32.271 85.057 32.335 ;
			RECT	85.361 32.271 85.393 32.335 ;
			RECT	85.697 32.271 85.729 32.335 ;
			RECT	86.033 32.271 86.065 32.335 ;
			RECT	86.369 32.271 86.401 32.335 ;
			RECT	86.705 32.271 86.737 32.335 ;
			RECT	87.041 32.271 87.073 32.335 ;
			RECT	87.377 32.271 87.409 32.335 ;
			RECT	87.713 32.271 87.745 32.335 ;
			RECT	88.049 32.271 88.081 32.335 ;
			RECT	88.385 32.271 88.417 32.335 ;
			RECT	88.721 32.271 88.753 32.335 ;
			RECT	89.057 32.271 89.089 32.335 ;
			RECT	89.393 32.271 89.425 32.335 ;
			RECT	89.729 32.271 89.761 32.335 ;
			RECT	90.065 32.271 90.097 32.335 ;
			RECT	90.401 32.271 90.433 32.335 ;
			RECT	90.737 32.271 90.769 32.335 ;
			RECT	91.073 32.271 91.105 32.335 ;
			RECT	91.409 32.271 91.441 32.335 ;
			RECT	91.745 32.271 91.777 32.335 ;
			RECT	92.081 32.271 92.113 32.335 ;
			RECT	92.417 32.271 92.449 32.335 ;
			RECT	92.753 32.271 92.785 32.335 ;
			RECT	93.089 32.271 93.121 32.335 ;
			RECT	93.425 32.271 93.457 32.335 ;
			RECT	93.761 32.271 93.793 32.335 ;
			RECT	94.097 32.271 94.129 32.335 ;
			RECT	94.433 32.271 94.465 32.335 ;
			RECT	94.769 32.271 94.801 32.335 ;
			RECT	95.105 32.271 95.137 32.335 ;
			RECT	95.441 32.271 95.473 32.335 ;
			RECT	95.777 32.271 95.809 32.335 ;
			RECT	96.113 32.271 96.145 32.335 ;
			RECT	96.449 32.271 96.481 32.335 ;
			RECT	96.785 32.271 96.817 32.335 ;
			RECT	97.121 32.271 97.153 32.335 ;
			RECT	97.457 32.271 97.489 32.335 ;
			RECT	97.793 32.271 97.825 32.335 ;
			RECT	98.129 32.271 98.161 32.335 ;
			RECT	98.465 32.271 98.497 32.335 ;
			RECT	98.801 32.271 98.833 32.335 ;
			RECT	99.137 32.271 99.169 32.335 ;
			RECT	99.473 32.271 99.505 32.335 ;
			RECT	99.809 32.271 99.841 32.335 ;
			RECT	100.145 32.271 100.177 32.335 ;
			RECT	100.481 32.271 100.513 32.335 ;
			RECT	100.817 32.271 100.849 32.335 ;
			RECT	101.153 32.271 101.185 32.335 ;
			RECT	101.489 32.271 101.521 32.335 ;
			RECT	101.825 32.271 101.857 32.335 ;
			RECT	104.345 32.271 104.377 32.335 ;
			RECT	104.681 32.271 104.713 32.335 ;
			RECT	105.017 32.271 105.049 32.335 ;
			RECT	105.353 32.271 105.385 32.335 ;
			RECT	105.689 32.271 105.721 32.335 ;
			RECT	106.025 32.271 106.057 32.335 ;
			RECT	106.361 32.271 106.393 32.335 ;
			RECT	106.697 32.271 106.729 32.335 ;
			RECT	107.033 32.271 107.065 32.335 ;
			RECT	107.369 32.271 107.401 32.335 ;
			RECT	107.705 32.271 107.737 32.335 ;
			RECT	108.041 32.271 108.073 32.335 ;
			RECT	108.377 32.271 108.409 32.335 ;
			RECT	108.713 32.271 108.745 32.335 ;
			RECT	109.049 32.271 109.081 32.335 ;
			RECT	109.385 32.271 109.417 32.335 ;
			RECT	109.721 32.271 109.753 32.335 ;
			RECT	110.057 32.271 110.089 32.335 ;
			RECT	110.393 32.271 110.425 32.335 ;
			RECT	110.729 32.271 110.761 32.335 ;
			RECT	111.065 32.271 111.097 32.335 ;
			RECT	111.401 32.271 111.433 32.335 ;
			RECT	111.737 32.271 111.769 32.335 ;
			RECT	112.073 32.271 112.105 32.335 ;
			RECT	112.409 32.271 112.441 32.335 ;
			RECT	112.745 32.271 112.777 32.335 ;
			RECT	113.081 32.271 113.113 32.335 ;
			RECT	113.417 32.271 113.449 32.335 ;
			RECT	113.753 32.271 113.785 32.335 ;
			RECT	114.089 32.271 114.121 32.335 ;
			RECT	114.425 32.271 114.457 32.335 ;
			RECT	114.761 32.271 114.793 32.335 ;
			RECT	115.097 32.271 115.129 32.335 ;
			RECT	115.433 32.271 115.465 32.335 ;
			RECT	115.769 32.271 115.801 32.335 ;
			RECT	116.105 32.271 116.137 32.335 ;
			RECT	116.441 32.271 116.473 32.335 ;
			RECT	116.777 32.271 116.809 32.335 ;
			RECT	117.113 32.271 117.145 32.335 ;
			RECT	117.449 32.271 117.481 32.335 ;
			RECT	117.785 32.271 117.817 32.335 ;
			RECT	118.121 32.271 118.153 32.335 ;
			RECT	118.457 32.271 118.489 32.335 ;
			RECT	118.793 32.271 118.825 32.335 ;
			RECT	119.129 32.271 119.161 32.335 ;
			RECT	119.465 32.271 119.497 32.335 ;
			RECT	119.801 32.271 119.833 32.335 ;
			RECT	120.137 32.271 120.169 32.335 ;
			RECT	120.473 32.271 120.505 32.335 ;
			RECT	120.809 32.271 120.841 32.335 ;
			RECT	121.145 32.271 121.177 32.335 ;
			RECT	121.481 32.271 121.513 32.335 ;
			RECT	121.817 32.271 121.849 32.335 ;
			RECT	122.153 32.271 122.185 32.335 ;
			RECT	122.489 32.271 122.521 32.335 ;
			RECT	122.825 32.271 122.857 32.335 ;
			RECT	123.161 32.271 123.193 32.335 ;
			RECT	123.497 32.271 123.529 32.335 ;
			RECT	123.833 32.271 123.865 32.335 ;
			RECT	124.169 32.271 124.201 32.335 ;
			RECT	124.505 32.271 124.537 32.335 ;
			RECT	124.841 32.271 124.873 32.335 ;
			RECT	125.177 32.271 125.209 32.335 ;
			RECT	125.513 32.271 125.545 32.335 ;
			RECT	147.309 32.271 147.373 32.335 ;
			RECT	150.122 32.271 150.154 32.335 ;
			RECT	150.576 32.271 150.608 32.335 ;
			RECT	150.966 32.271 151.03 32.335 ;
			RECT	152.249 32.271 152.281 32.335 ;
			RECT	153.56 32.271 153.624 32.335 ;
			RECT	153.801 32.271 153.833 32.335 ;
			RECT	156.827 32.271 156.891 32.335 ;
			RECT	178.655 32.271 178.687 32.335 ;
			RECT	178.991 32.271 179.023 32.335 ;
			RECT	179.327 32.271 179.359 32.335 ;
			RECT	179.663 32.271 179.695 32.335 ;
			RECT	179.999 32.271 180.031 32.335 ;
			RECT	180.335 32.271 180.367 32.335 ;
			RECT	180.671 32.271 180.703 32.335 ;
			RECT	181.007 32.271 181.039 32.335 ;
			RECT	181.343 32.271 181.375 32.335 ;
			RECT	181.679 32.271 181.711 32.335 ;
			RECT	182.015 32.271 182.047 32.335 ;
			RECT	182.351 32.271 182.383 32.335 ;
			RECT	182.687 32.271 182.719 32.335 ;
			RECT	183.023 32.271 183.055 32.335 ;
			RECT	183.359 32.271 183.391 32.335 ;
			RECT	183.695 32.271 183.727 32.335 ;
			RECT	184.031 32.271 184.063 32.335 ;
			RECT	184.367 32.271 184.399 32.335 ;
			RECT	184.703 32.271 184.735 32.335 ;
			RECT	185.039 32.271 185.071 32.335 ;
			RECT	185.375 32.271 185.407 32.335 ;
			RECT	185.711 32.271 185.743 32.335 ;
			RECT	186.047 32.271 186.079 32.335 ;
			RECT	186.383 32.271 186.415 32.335 ;
			RECT	186.719 32.271 186.751 32.335 ;
			RECT	187.055 32.271 187.087 32.335 ;
			RECT	187.391 32.271 187.423 32.335 ;
			RECT	187.727 32.271 187.759 32.335 ;
			RECT	188.063 32.271 188.095 32.335 ;
			RECT	188.399 32.271 188.431 32.335 ;
			RECT	188.735 32.271 188.767 32.335 ;
			RECT	189.071 32.271 189.103 32.335 ;
			RECT	189.407 32.271 189.439 32.335 ;
			RECT	189.743 32.271 189.775 32.335 ;
			RECT	190.079 32.271 190.111 32.335 ;
			RECT	190.415 32.271 190.447 32.335 ;
			RECT	190.751 32.271 190.783 32.335 ;
			RECT	191.087 32.271 191.119 32.335 ;
			RECT	191.423 32.271 191.455 32.335 ;
			RECT	191.759 32.271 191.791 32.335 ;
			RECT	192.095 32.271 192.127 32.335 ;
			RECT	192.431 32.271 192.463 32.335 ;
			RECT	192.767 32.271 192.799 32.335 ;
			RECT	193.103 32.271 193.135 32.335 ;
			RECT	193.439 32.271 193.471 32.335 ;
			RECT	193.775 32.271 193.807 32.335 ;
			RECT	194.111 32.271 194.143 32.335 ;
			RECT	194.447 32.271 194.479 32.335 ;
			RECT	194.783 32.271 194.815 32.335 ;
			RECT	195.119 32.271 195.151 32.335 ;
			RECT	195.455 32.271 195.487 32.335 ;
			RECT	195.791 32.271 195.823 32.335 ;
			RECT	196.127 32.271 196.159 32.335 ;
			RECT	196.463 32.271 196.495 32.335 ;
			RECT	196.799 32.271 196.831 32.335 ;
			RECT	197.135 32.271 197.167 32.335 ;
			RECT	197.471 32.271 197.503 32.335 ;
			RECT	197.807 32.271 197.839 32.335 ;
			RECT	198.143 32.271 198.175 32.335 ;
			RECT	198.479 32.271 198.511 32.335 ;
			RECT	198.815 32.271 198.847 32.335 ;
			RECT	199.151 32.271 199.183 32.335 ;
			RECT	199.487 32.271 199.519 32.335 ;
			RECT	199.823 32.271 199.855 32.335 ;
			RECT	201.403 32.271 201.435 32.335 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 33.238 201.665 33.348 ;
			LAYER	J3 ;
			RECT	0.755 33.261 0.787 33.325 ;
			RECT	1.645 33.261 1.709 33.325 ;
			RECT	2.124 33.261 2.156 33.325 ;
			RECT	2.323 33.277 2.387 33.309 ;
			RECT	3.438 33.261 3.47 33.325 ;
			RECT	4.195 33.261 4.227 33.325 ;
			RECT	4.944 33.261 5.008 33.325 ;
			RECT	6.347 33.261 6.379 33.325 ;
			RECT	6.683 33.261 6.715 33.325 ;
			RECT	7.019 33.261 7.051 33.325 ;
			RECT	7.355 33.261 7.387 33.325 ;
			RECT	7.691 33.261 7.723 33.325 ;
			RECT	8.027 33.261 8.059 33.325 ;
			RECT	8.363 33.261 8.395 33.325 ;
			RECT	8.699 33.261 8.731 33.325 ;
			RECT	9.035 33.261 9.067 33.325 ;
			RECT	9.371 33.261 9.403 33.325 ;
			RECT	9.707 33.261 9.739 33.325 ;
			RECT	10.043 33.261 10.075 33.325 ;
			RECT	10.379 33.261 10.411 33.325 ;
			RECT	10.715 33.261 10.747 33.325 ;
			RECT	11.051 33.261 11.083 33.325 ;
			RECT	11.387 33.261 11.419 33.325 ;
			RECT	11.723 33.261 11.755 33.325 ;
			RECT	12.059 33.261 12.091 33.325 ;
			RECT	12.395 33.261 12.427 33.325 ;
			RECT	12.731 33.261 12.763 33.325 ;
			RECT	13.067 33.261 13.099 33.325 ;
			RECT	13.403 33.261 13.435 33.325 ;
			RECT	13.739 33.261 13.771 33.325 ;
			RECT	14.075 33.261 14.107 33.325 ;
			RECT	14.411 33.261 14.443 33.325 ;
			RECT	14.747 33.261 14.779 33.325 ;
			RECT	15.083 33.261 15.115 33.325 ;
			RECT	15.419 33.261 15.451 33.325 ;
			RECT	15.755 33.261 15.787 33.325 ;
			RECT	16.091 33.261 16.123 33.325 ;
			RECT	16.427 33.261 16.459 33.325 ;
			RECT	16.763 33.261 16.795 33.325 ;
			RECT	17.099 33.261 17.131 33.325 ;
			RECT	17.435 33.261 17.467 33.325 ;
			RECT	17.771 33.261 17.803 33.325 ;
			RECT	18.107 33.261 18.139 33.325 ;
			RECT	18.443 33.261 18.475 33.325 ;
			RECT	18.779 33.261 18.811 33.325 ;
			RECT	19.115 33.261 19.147 33.325 ;
			RECT	19.451 33.261 19.483 33.325 ;
			RECT	19.787 33.261 19.819 33.325 ;
			RECT	20.123 33.261 20.155 33.325 ;
			RECT	20.459 33.261 20.491 33.325 ;
			RECT	20.795 33.261 20.827 33.325 ;
			RECT	21.131 33.261 21.163 33.325 ;
			RECT	21.467 33.261 21.499 33.325 ;
			RECT	21.803 33.261 21.835 33.325 ;
			RECT	22.139 33.261 22.171 33.325 ;
			RECT	22.475 33.261 22.507 33.325 ;
			RECT	22.811 33.261 22.843 33.325 ;
			RECT	23.147 33.261 23.179 33.325 ;
			RECT	23.483 33.261 23.515 33.325 ;
			RECT	23.819 33.261 23.851 33.325 ;
			RECT	24.155 33.261 24.187 33.325 ;
			RECT	24.491 33.261 24.523 33.325 ;
			RECT	24.827 33.261 24.859 33.325 ;
			RECT	25.163 33.261 25.195 33.325 ;
			RECT	25.499 33.261 25.531 33.325 ;
			RECT	25.835 33.261 25.867 33.325 ;
			RECT	26.171 33.261 26.203 33.325 ;
			RECT	26.507 33.261 26.539 33.325 ;
			RECT	26.843 33.261 26.875 33.325 ;
			RECT	27.179 33.261 27.211 33.325 ;
			RECT	27.515 33.261 27.547 33.325 ;
			RECT	27.851 33.261 27.883 33.325 ;
			RECT	28.019 33.261 28.051 33.325 ;
			RECT	28.187 33.261 28.219 33.325 ;
			RECT	28.355 33.261 28.387 33.325 ;
			RECT	28.523 33.261 28.555 33.325 ;
			RECT	28.691 33.261 28.723 33.325 ;
			RECT	28.859 33.261 28.891 33.325 ;
			RECT	29.027 33.261 29.059 33.325 ;
			RECT	29.195 33.261 29.227 33.325 ;
			RECT	29.363 33.261 29.395 33.325 ;
			RECT	29.531 33.261 29.563 33.325 ;
			RECT	29.699 33.261 29.731 33.325 ;
			RECT	29.867 33.261 29.899 33.325 ;
			RECT	30.035 33.261 30.067 33.325 ;
			RECT	30.203 33.261 30.235 33.325 ;
			RECT	30.371 33.261 30.403 33.325 ;
			RECT	30.539 33.261 30.571 33.325 ;
			RECT	30.707 33.261 30.739 33.325 ;
			RECT	30.875 33.261 30.907 33.325 ;
			RECT	31.043 33.261 31.075 33.325 ;
			RECT	31.211 33.261 31.243 33.325 ;
			RECT	31.379 33.261 31.411 33.325 ;
			RECT	31.547 33.261 31.579 33.325 ;
			RECT	31.715 33.261 31.747 33.325 ;
			RECT	31.883 33.261 31.915 33.325 ;
			RECT	32.051 33.261 32.083 33.325 ;
			RECT	32.219 33.261 32.251 33.325 ;
			RECT	32.387 33.261 32.419 33.325 ;
			RECT	32.555 33.261 32.587 33.325 ;
			RECT	32.723 33.261 32.755 33.325 ;
			RECT	32.891 33.261 32.923 33.325 ;
			RECT	33.059 33.261 33.091 33.325 ;
			RECT	33.227 33.261 33.259 33.325 ;
			RECT	33.395 33.261 33.427 33.325 ;
			RECT	33.563 33.261 33.595 33.325 ;
			RECT	33.731 33.261 33.763 33.325 ;
			RECT	33.899 33.261 33.931 33.325 ;
			RECT	34.067 33.261 34.099 33.325 ;
			RECT	34.235 33.261 34.267 33.325 ;
			RECT	34.403 33.261 34.435 33.325 ;
			RECT	34.571 33.261 34.603 33.325 ;
			RECT	34.739 33.261 34.771 33.325 ;
			RECT	34.907 33.261 34.939 33.325 ;
			RECT	35.075 33.261 35.107 33.325 ;
			RECT	35.243 33.261 35.275 33.325 ;
			RECT	35.411 33.261 35.443 33.325 ;
			RECT	35.579 33.261 35.611 33.325 ;
			RECT	35.747 33.261 35.779 33.325 ;
			RECT	35.915 33.261 35.947 33.325 ;
			RECT	36.083 33.261 36.115 33.325 ;
			RECT	36.251 33.261 36.283 33.325 ;
			RECT	36.419 33.261 36.451 33.325 ;
			RECT	36.587 33.261 36.619 33.325 ;
			RECT	36.755 33.261 36.787 33.325 ;
			RECT	36.923 33.261 36.955 33.325 ;
			RECT	37.091 33.261 37.123 33.325 ;
			RECT	37.259 33.261 37.291 33.325 ;
			RECT	37.427 33.261 37.459 33.325 ;
			RECT	37.595 33.261 37.627 33.325 ;
			RECT	37.763 33.261 37.795 33.325 ;
			RECT	37.931 33.261 37.963 33.325 ;
			RECT	38.099 33.261 38.131 33.325 ;
			RECT	38.267 33.261 38.299 33.325 ;
			RECT	38.435 33.261 38.467 33.325 ;
			RECT	38.603 33.261 38.635 33.325 ;
			RECT	38.771 33.261 38.803 33.325 ;
			RECT	38.939 33.261 38.971 33.325 ;
			RECT	39.107 33.261 39.139 33.325 ;
			RECT	39.275 33.261 39.307 33.325 ;
			RECT	39.443 33.261 39.475 33.325 ;
			RECT	39.611 33.261 39.643 33.325 ;
			RECT	39.779 33.261 39.811 33.325 ;
			RECT	39.947 33.261 39.979 33.325 ;
			RECT	40.115 33.261 40.147 33.325 ;
			RECT	40.283 33.261 40.315 33.325 ;
			RECT	40.451 33.261 40.483 33.325 ;
			RECT	40.619 33.261 40.651 33.325 ;
			RECT	40.787 33.261 40.819 33.325 ;
			RECT	40.955 33.261 40.987 33.325 ;
			RECT	41.123 33.261 41.155 33.325 ;
			RECT	41.291 33.261 41.323 33.325 ;
			RECT	41.459 33.261 41.491 33.325 ;
			RECT	41.627 33.261 41.659 33.325 ;
			RECT	41.795 33.261 41.827 33.325 ;
			RECT	41.963 33.261 41.995 33.325 ;
			RECT	42.131 33.261 42.163 33.325 ;
			RECT	42.299 33.261 42.331 33.325 ;
			RECT	42.467 33.261 42.499 33.325 ;
			RECT	42.635 33.261 42.667 33.325 ;
			RECT	42.803 33.261 42.835 33.325 ;
			RECT	42.971 33.261 43.003 33.325 ;
			RECT	43.139 33.261 43.171 33.325 ;
			RECT	43.307 33.261 43.339 33.325 ;
			RECT	43.475 33.261 43.507 33.325 ;
			RECT	43.643 33.261 43.675 33.325 ;
			RECT	43.811 33.261 43.843 33.325 ;
			RECT	43.979 33.261 44.011 33.325 ;
			RECT	44.147 33.261 44.179 33.325 ;
			RECT	44.315 33.261 44.347 33.325 ;
			RECT	44.483 33.261 44.515 33.325 ;
			RECT	44.651 33.261 44.683 33.325 ;
			RECT	44.819 33.261 44.851 33.325 ;
			RECT	44.987 33.261 45.019 33.325 ;
			RECT	45.155 33.261 45.187 33.325 ;
			RECT	45.323 33.261 45.355 33.325 ;
			RECT	45.491 33.261 45.523 33.325 ;
			RECT	45.659 33.261 45.691 33.325 ;
			RECT	45.827 33.261 45.859 33.325 ;
			RECT	45.995 33.261 46.027 33.325 ;
			RECT	46.163 33.261 46.195 33.325 ;
			RECT	46.331 33.261 46.363 33.325 ;
			RECT	46.499 33.261 46.531 33.325 ;
			RECT	46.667 33.261 46.699 33.325 ;
			RECT	46.835 33.261 46.867 33.325 ;
			RECT	47.003 33.261 47.035 33.325 ;
			RECT	47.171 33.261 47.203 33.325 ;
			RECT	47.339 33.261 47.371 33.325 ;
			RECT	47.507 33.261 47.539 33.325 ;
			RECT	47.675 33.261 47.707 33.325 ;
			RECT	47.843 33.261 47.875 33.325 ;
			RECT	48.011 33.261 48.043 33.325 ;
			RECT	48.179 33.261 48.211 33.325 ;
			RECT	48.347 33.261 48.379 33.325 ;
			RECT	48.515 33.261 48.547 33.325 ;
			RECT	48.683 33.261 48.715 33.325 ;
			RECT	48.851 33.261 48.883 33.325 ;
			RECT	49.019 33.261 49.051 33.325 ;
			RECT	49.327 33.261 49.359 33.325 ;
			RECT	49.613 33.261 49.645 33.325 ;
			RECT	52.578 33.261 52.61 33.325 ;
			RECT	52.968 33.261 53.032 33.325 ;
			RECT	53.91 33.261 53.942 33.325 ;
			RECT	54.251 33.261 54.283 33.325 ;
			RECT	55.562 33.261 55.626 33.325 ;
			RECT	55.803 33.261 55.835 33.325 ;
			RECT	55.969 33.261 56.033 33.325 ;
			RECT	58.559 33.261 58.591 33.325 ;
			RECT	58.845 33.261 58.877 33.325 ;
			RECT	59.153 33.261 59.185 33.325 ;
			RECT	59.321 33.261 59.353 33.325 ;
			RECT	59.489 33.261 59.521 33.325 ;
			RECT	59.657 33.261 59.689 33.325 ;
			RECT	59.825 33.261 59.857 33.325 ;
			RECT	59.993 33.261 60.025 33.325 ;
			RECT	60.161 33.261 60.193 33.325 ;
			RECT	60.329 33.261 60.361 33.325 ;
			RECT	60.497 33.261 60.529 33.325 ;
			RECT	60.665 33.261 60.697 33.325 ;
			RECT	60.833 33.261 60.865 33.325 ;
			RECT	61.001 33.261 61.033 33.325 ;
			RECT	61.169 33.261 61.201 33.325 ;
			RECT	61.337 33.261 61.369 33.325 ;
			RECT	61.505 33.261 61.537 33.325 ;
			RECT	61.673 33.261 61.705 33.325 ;
			RECT	61.841 33.261 61.873 33.325 ;
			RECT	62.009 33.261 62.041 33.325 ;
			RECT	62.177 33.261 62.209 33.325 ;
			RECT	62.345 33.261 62.377 33.325 ;
			RECT	62.513 33.261 62.545 33.325 ;
			RECT	62.681 33.261 62.713 33.325 ;
			RECT	62.849 33.261 62.881 33.325 ;
			RECT	63.017 33.261 63.049 33.325 ;
			RECT	63.185 33.261 63.217 33.325 ;
			RECT	63.353 33.261 63.385 33.325 ;
			RECT	63.521 33.261 63.553 33.325 ;
			RECT	63.689 33.261 63.721 33.325 ;
			RECT	63.857 33.261 63.889 33.325 ;
			RECT	64.025 33.261 64.057 33.325 ;
			RECT	64.193 33.261 64.225 33.325 ;
			RECT	64.361 33.261 64.393 33.325 ;
			RECT	64.529 33.261 64.561 33.325 ;
			RECT	64.697 33.261 64.729 33.325 ;
			RECT	64.865 33.261 64.897 33.325 ;
			RECT	65.033 33.261 65.065 33.325 ;
			RECT	65.201 33.261 65.233 33.325 ;
			RECT	65.369 33.261 65.401 33.325 ;
			RECT	65.537 33.261 65.569 33.325 ;
			RECT	65.705 33.261 65.737 33.325 ;
			RECT	65.873 33.261 65.905 33.325 ;
			RECT	66.041 33.261 66.073 33.325 ;
			RECT	66.209 33.261 66.241 33.325 ;
			RECT	66.377 33.261 66.409 33.325 ;
			RECT	66.545 33.261 66.577 33.325 ;
			RECT	66.713 33.261 66.745 33.325 ;
			RECT	66.881 33.261 66.913 33.325 ;
			RECT	67.049 33.261 67.081 33.325 ;
			RECT	67.217 33.261 67.249 33.325 ;
			RECT	67.385 33.261 67.417 33.325 ;
			RECT	67.553 33.261 67.585 33.325 ;
			RECT	67.721 33.261 67.753 33.325 ;
			RECT	67.889 33.261 67.921 33.325 ;
			RECT	68.057 33.261 68.089 33.325 ;
			RECT	68.225 33.261 68.257 33.325 ;
			RECT	68.393 33.261 68.425 33.325 ;
			RECT	68.561 33.261 68.593 33.325 ;
			RECT	68.729 33.261 68.761 33.325 ;
			RECT	68.897 33.261 68.929 33.325 ;
			RECT	69.065 33.261 69.097 33.325 ;
			RECT	69.233 33.261 69.265 33.325 ;
			RECT	69.401 33.261 69.433 33.325 ;
			RECT	69.569 33.261 69.601 33.325 ;
			RECT	69.737 33.261 69.769 33.325 ;
			RECT	69.905 33.261 69.937 33.325 ;
			RECT	70.073 33.261 70.105 33.325 ;
			RECT	70.241 33.261 70.273 33.325 ;
			RECT	70.409 33.261 70.441 33.325 ;
			RECT	70.577 33.261 70.609 33.325 ;
			RECT	70.745 33.261 70.777 33.325 ;
			RECT	70.913 33.261 70.945 33.325 ;
			RECT	71.081 33.261 71.113 33.325 ;
			RECT	71.249 33.261 71.281 33.325 ;
			RECT	71.417 33.261 71.449 33.325 ;
			RECT	71.585 33.261 71.617 33.325 ;
			RECT	71.753 33.261 71.785 33.325 ;
			RECT	71.921 33.261 71.953 33.325 ;
			RECT	72.089 33.261 72.121 33.325 ;
			RECT	72.257 33.261 72.289 33.325 ;
			RECT	72.425 33.261 72.457 33.325 ;
			RECT	72.593 33.261 72.625 33.325 ;
			RECT	72.761 33.261 72.793 33.325 ;
			RECT	72.929 33.261 72.961 33.325 ;
			RECT	73.097 33.261 73.129 33.325 ;
			RECT	73.265 33.261 73.297 33.325 ;
			RECT	73.433 33.261 73.465 33.325 ;
			RECT	73.601 33.261 73.633 33.325 ;
			RECT	73.769 33.261 73.801 33.325 ;
			RECT	73.937 33.261 73.969 33.325 ;
			RECT	74.105 33.261 74.137 33.325 ;
			RECT	74.273 33.261 74.305 33.325 ;
			RECT	74.441 33.261 74.473 33.325 ;
			RECT	74.609 33.261 74.641 33.325 ;
			RECT	74.777 33.261 74.809 33.325 ;
			RECT	74.945 33.261 74.977 33.325 ;
			RECT	75.113 33.261 75.145 33.325 ;
			RECT	75.281 33.261 75.313 33.325 ;
			RECT	75.449 33.261 75.481 33.325 ;
			RECT	75.617 33.261 75.649 33.325 ;
			RECT	75.785 33.261 75.817 33.325 ;
			RECT	75.953 33.261 75.985 33.325 ;
			RECT	76.121 33.261 76.153 33.325 ;
			RECT	76.289 33.261 76.321 33.325 ;
			RECT	76.457 33.261 76.489 33.325 ;
			RECT	76.625 33.261 76.657 33.325 ;
			RECT	76.793 33.261 76.825 33.325 ;
			RECT	76.961 33.261 76.993 33.325 ;
			RECT	77.129 33.261 77.161 33.325 ;
			RECT	77.297 33.261 77.329 33.325 ;
			RECT	77.465 33.261 77.497 33.325 ;
			RECT	77.633 33.261 77.665 33.325 ;
			RECT	77.801 33.261 77.833 33.325 ;
			RECT	77.969 33.261 78.001 33.325 ;
			RECT	78.137 33.261 78.169 33.325 ;
			RECT	78.305 33.261 78.337 33.325 ;
			RECT	78.473 33.261 78.505 33.325 ;
			RECT	78.641 33.261 78.673 33.325 ;
			RECT	78.809 33.261 78.841 33.325 ;
			RECT	78.977 33.261 79.009 33.325 ;
			RECT	79.145 33.261 79.177 33.325 ;
			RECT	79.313 33.261 79.345 33.325 ;
			RECT	79.481 33.261 79.513 33.325 ;
			RECT	79.649 33.261 79.681 33.325 ;
			RECT	79.817 33.261 79.849 33.325 ;
			RECT	79.985 33.261 80.017 33.325 ;
			RECT	80.153 33.261 80.185 33.325 ;
			RECT	80.321 33.261 80.353 33.325 ;
			RECT	80.657 33.261 80.689 33.325 ;
			RECT	80.993 33.261 81.025 33.325 ;
			RECT	81.329 33.261 81.361 33.325 ;
			RECT	81.665 33.261 81.697 33.325 ;
			RECT	82.001 33.261 82.033 33.325 ;
			RECT	82.337 33.261 82.369 33.325 ;
			RECT	82.673 33.261 82.705 33.325 ;
			RECT	83.009 33.261 83.041 33.325 ;
			RECT	83.345 33.261 83.377 33.325 ;
			RECT	83.681 33.261 83.713 33.325 ;
			RECT	84.017 33.261 84.049 33.325 ;
			RECT	84.353 33.261 84.385 33.325 ;
			RECT	84.689 33.261 84.721 33.325 ;
			RECT	85.025 33.261 85.057 33.325 ;
			RECT	85.361 33.261 85.393 33.325 ;
			RECT	85.697 33.261 85.729 33.325 ;
			RECT	86.033 33.261 86.065 33.325 ;
			RECT	86.369 33.261 86.401 33.325 ;
			RECT	86.705 33.261 86.737 33.325 ;
			RECT	87.041 33.261 87.073 33.325 ;
			RECT	87.377 33.261 87.409 33.325 ;
			RECT	87.713 33.261 87.745 33.325 ;
			RECT	88.049 33.261 88.081 33.325 ;
			RECT	88.385 33.261 88.417 33.325 ;
			RECT	88.721 33.261 88.753 33.325 ;
			RECT	89.057 33.261 89.089 33.325 ;
			RECT	89.393 33.261 89.425 33.325 ;
			RECT	89.729 33.261 89.761 33.325 ;
			RECT	90.065 33.261 90.097 33.325 ;
			RECT	90.401 33.261 90.433 33.325 ;
			RECT	90.737 33.261 90.769 33.325 ;
			RECT	91.073 33.261 91.105 33.325 ;
			RECT	91.409 33.261 91.441 33.325 ;
			RECT	91.745 33.261 91.777 33.325 ;
			RECT	92.081 33.261 92.113 33.325 ;
			RECT	92.417 33.261 92.449 33.325 ;
			RECT	92.753 33.261 92.785 33.325 ;
			RECT	93.089 33.261 93.121 33.325 ;
			RECT	93.425 33.261 93.457 33.325 ;
			RECT	93.761 33.261 93.793 33.325 ;
			RECT	94.097 33.261 94.129 33.325 ;
			RECT	94.433 33.261 94.465 33.325 ;
			RECT	94.769 33.261 94.801 33.325 ;
			RECT	95.105 33.261 95.137 33.325 ;
			RECT	95.441 33.261 95.473 33.325 ;
			RECT	95.777 33.261 95.809 33.325 ;
			RECT	96.113 33.261 96.145 33.325 ;
			RECT	96.449 33.261 96.481 33.325 ;
			RECT	96.785 33.261 96.817 33.325 ;
			RECT	97.121 33.261 97.153 33.325 ;
			RECT	97.457 33.261 97.489 33.325 ;
			RECT	97.793 33.261 97.825 33.325 ;
			RECT	98.129 33.261 98.161 33.325 ;
			RECT	98.465 33.261 98.497 33.325 ;
			RECT	98.801 33.261 98.833 33.325 ;
			RECT	99.137 33.261 99.169 33.325 ;
			RECT	99.473 33.261 99.505 33.325 ;
			RECT	99.809 33.261 99.841 33.325 ;
			RECT	100.145 33.261 100.177 33.325 ;
			RECT	100.481 33.261 100.513 33.325 ;
			RECT	100.817 33.261 100.849 33.325 ;
			RECT	101.153 33.261 101.185 33.325 ;
			RECT	101.489 33.261 101.521 33.325 ;
			RECT	101.825 33.261 101.857 33.325 ;
			RECT	102.995 33.261 103.027 33.325 ;
			RECT	103.175 33.261 103.207 33.325 ;
			RECT	104.345 33.261 104.377 33.325 ;
			RECT	104.681 33.261 104.713 33.325 ;
			RECT	105.017 33.261 105.049 33.325 ;
			RECT	105.353 33.261 105.385 33.325 ;
			RECT	105.689 33.261 105.721 33.325 ;
			RECT	106.025 33.261 106.057 33.325 ;
			RECT	106.361 33.261 106.393 33.325 ;
			RECT	106.697 33.261 106.729 33.325 ;
			RECT	107.033 33.261 107.065 33.325 ;
			RECT	107.369 33.261 107.401 33.325 ;
			RECT	107.705 33.261 107.737 33.325 ;
			RECT	108.041 33.261 108.073 33.325 ;
			RECT	108.377 33.261 108.409 33.325 ;
			RECT	108.713 33.261 108.745 33.325 ;
			RECT	109.049 33.261 109.081 33.325 ;
			RECT	109.385 33.261 109.417 33.325 ;
			RECT	109.721 33.261 109.753 33.325 ;
			RECT	110.057 33.261 110.089 33.325 ;
			RECT	110.393 33.261 110.425 33.325 ;
			RECT	110.729 33.261 110.761 33.325 ;
			RECT	111.065 33.261 111.097 33.325 ;
			RECT	111.401 33.261 111.433 33.325 ;
			RECT	111.737 33.261 111.769 33.325 ;
			RECT	112.073 33.261 112.105 33.325 ;
			RECT	112.409 33.261 112.441 33.325 ;
			RECT	112.745 33.261 112.777 33.325 ;
			RECT	113.081 33.261 113.113 33.325 ;
			RECT	113.417 33.261 113.449 33.325 ;
			RECT	113.753 33.261 113.785 33.325 ;
			RECT	114.089 33.261 114.121 33.325 ;
			RECT	114.425 33.261 114.457 33.325 ;
			RECT	114.761 33.261 114.793 33.325 ;
			RECT	115.097 33.261 115.129 33.325 ;
			RECT	115.433 33.261 115.465 33.325 ;
			RECT	115.769 33.261 115.801 33.325 ;
			RECT	116.105 33.261 116.137 33.325 ;
			RECT	116.441 33.261 116.473 33.325 ;
			RECT	116.777 33.261 116.809 33.325 ;
			RECT	117.113 33.261 117.145 33.325 ;
			RECT	117.449 33.261 117.481 33.325 ;
			RECT	117.785 33.261 117.817 33.325 ;
			RECT	118.121 33.261 118.153 33.325 ;
			RECT	118.457 33.261 118.489 33.325 ;
			RECT	118.793 33.261 118.825 33.325 ;
			RECT	119.129 33.261 119.161 33.325 ;
			RECT	119.465 33.261 119.497 33.325 ;
			RECT	119.801 33.261 119.833 33.325 ;
			RECT	120.137 33.261 120.169 33.325 ;
			RECT	120.473 33.261 120.505 33.325 ;
			RECT	120.809 33.261 120.841 33.325 ;
			RECT	121.145 33.261 121.177 33.325 ;
			RECT	121.481 33.261 121.513 33.325 ;
			RECT	121.817 33.261 121.849 33.325 ;
			RECT	122.153 33.261 122.185 33.325 ;
			RECT	122.489 33.261 122.521 33.325 ;
			RECT	122.825 33.261 122.857 33.325 ;
			RECT	123.161 33.261 123.193 33.325 ;
			RECT	123.497 33.261 123.529 33.325 ;
			RECT	123.833 33.261 123.865 33.325 ;
			RECT	124.169 33.261 124.201 33.325 ;
			RECT	124.505 33.261 124.537 33.325 ;
			RECT	124.841 33.261 124.873 33.325 ;
			RECT	125.177 33.261 125.209 33.325 ;
			RECT	125.513 33.261 125.545 33.325 ;
			RECT	125.849 33.261 125.881 33.325 ;
			RECT	126.017 33.261 126.049 33.325 ;
			RECT	126.185 33.261 126.217 33.325 ;
			RECT	126.353 33.261 126.385 33.325 ;
			RECT	126.521 33.261 126.553 33.325 ;
			RECT	126.689 33.261 126.721 33.325 ;
			RECT	126.857 33.261 126.889 33.325 ;
			RECT	127.025 33.261 127.057 33.325 ;
			RECT	127.193 33.261 127.225 33.325 ;
			RECT	127.361 33.261 127.393 33.325 ;
			RECT	127.529 33.261 127.561 33.325 ;
			RECT	127.697 33.261 127.729 33.325 ;
			RECT	127.865 33.261 127.897 33.325 ;
			RECT	128.033 33.261 128.065 33.325 ;
			RECT	128.201 33.261 128.233 33.325 ;
			RECT	128.369 33.261 128.401 33.325 ;
			RECT	128.537 33.261 128.569 33.325 ;
			RECT	128.705 33.261 128.737 33.325 ;
			RECT	128.873 33.261 128.905 33.325 ;
			RECT	129.041 33.261 129.073 33.325 ;
			RECT	129.209 33.261 129.241 33.325 ;
			RECT	129.377 33.261 129.409 33.325 ;
			RECT	129.545 33.261 129.577 33.325 ;
			RECT	129.713 33.261 129.745 33.325 ;
			RECT	129.881 33.261 129.913 33.325 ;
			RECT	130.049 33.261 130.081 33.325 ;
			RECT	130.217 33.261 130.249 33.325 ;
			RECT	130.385 33.261 130.417 33.325 ;
			RECT	130.553 33.261 130.585 33.325 ;
			RECT	130.721 33.261 130.753 33.325 ;
			RECT	130.889 33.261 130.921 33.325 ;
			RECT	131.057 33.261 131.089 33.325 ;
			RECT	131.225 33.261 131.257 33.325 ;
			RECT	131.393 33.261 131.425 33.325 ;
			RECT	131.561 33.261 131.593 33.325 ;
			RECT	131.729 33.261 131.761 33.325 ;
			RECT	131.897 33.261 131.929 33.325 ;
			RECT	132.065 33.261 132.097 33.325 ;
			RECT	132.233 33.261 132.265 33.325 ;
			RECT	132.401 33.261 132.433 33.325 ;
			RECT	132.569 33.261 132.601 33.325 ;
			RECT	132.737 33.261 132.769 33.325 ;
			RECT	132.905 33.261 132.937 33.325 ;
			RECT	133.073 33.261 133.105 33.325 ;
			RECT	133.241 33.261 133.273 33.325 ;
			RECT	133.409 33.261 133.441 33.325 ;
			RECT	133.577 33.261 133.609 33.325 ;
			RECT	133.745 33.261 133.777 33.325 ;
			RECT	133.913 33.261 133.945 33.325 ;
			RECT	134.081 33.261 134.113 33.325 ;
			RECT	134.249 33.261 134.281 33.325 ;
			RECT	134.417 33.261 134.449 33.325 ;
			RECT	134.585 33.261 134.617 33.325 ;
			RECT	134.753 33.261 134.785 33.325 ;
			RECT	134.921 33.261 134.953 33.325 ;
			RECT	135.089 33.261 135.121 33.325 ;
			RECT	135.257 33.261 135.289 33.325 ;
			RECT	135.425 33.261 135.457 33.325 ;
			RECT	135.593 33.261 135.625 33.325 ;
			RECT	135.761 33.261 135.793 33.325 ;
			RECT	135.929 33.261 135.961 33.325 ;
			RECT	136.097 33.261 136.129 33.325 ;
			RECT	136.265 33.261 136.297 33.325 ;
			RECT	136.433 33.261 136.465 33.325 ;
			RECT	136.601 33.261 136.633 33.325 ;
			RECT	136.769 33.261 136.801 33.325 ;
			RECT	136.937 33.261 136.969 33.325 ;
			RECT	137.105 33.261 137.137 33.325 ;
			RECT	137.273 33.261 137.305 33.325 ;
			RECT	137.441 33.261 137.473 33.325 ;
			RECT	137.609 33.261 137.641 33.325 ;
			RECT	137.777 33.261 137.809 33.325 ;
			RECT	137.945 33.261 137.977 33.325 ;
			RECT	138.113 33.261 138.145 33.325 ;
			RECT	138.281 33.261 138.313 33.325 ;
			RECT	138.449 33.261 138.481 33.325 ;
			RECT	138.617 33.261 138.649 33.325 ;
			RECT	138.785 33.261 138.817 33.325 ;
			RECT	138.953 33.261 138.985 33.325 ;
			RECT	139.121 33.261 139.153 33.325 ;
			RECT	139.289 33.261 139.321 33.325 ;
			RECT	139.457 33.261 139.489 33.325 ;
			RECT	139.625 33.261 139.657 33.325 ;
			RECT	139.793 33.261 139.825 33.325 ;
			RECT	139.961 33.261 139.993 33.325 ;
			RECT	140.129 33.261 140.161 33.325 ;
			RECT	140.297 33.261 140.329 33.325 ;
			RECT	140.465 33.261 140.497 33.325 ;
			RECT	140.633 33.261 140.665 33.325 ;
			RECT	140.801 33.261 140.833 33.325 ;
			RECT	140.969 33.261 141.001 33.325 ;
			RECT	141.137 33.261 141.169 33.325 ;
			RECT	141.305 33.261 141.337 33.325 ;
			RECT	141.473 33.261 141.505 33.325 ;
			RECT	141.641 33.261 141.673 33.325 ;
			RECT	141.809 33.261 141.841 33.325 ;
			RECT	141.977 33.261 142.009 33.325 ;
			RECT	142.145 33.261 142.177 33.325 ;
			RECT	142.313 33.261 142.345 33.325 ;
			RECT	142.481 33.261 142.513 33.325 ;
			RECT	142.649 33.261 142.681 33.325 ;
			RECT	142.817 33.261 142.849 33.325 ;
			RECT	142.985 33.261 143.017 33.325 ;
			RECT	143.153 33.261 143.185 33.325 ;
			RECT	143.321 33.261 143.353 33.325 ;
			RECT	143.489 33.261 143.521 33.325 ;
			RECT	143.657 33.261 143.689 33.325 ;
			RECT	143.825 33.261 143.857 33.325 ;
			RECT	143.993 33.261 144.025 33.325 ;
			RECT	144.161 33.261 144.193 33.325 ;
			RECT	144.329 33.261 144.361 33.325 ;
			RECT	144.497 33.261 144.529 33.325 ;
			RECT	144.665 33.261 144.697 33.325 ;
			RECT	144.833 33.261 144.865 33.325 ;
			RECT	145.001 33.261 145.033 33.325 ;
			RECT	145.169 33.261 145.201 33.325 ;
			RECT	145.337 33.261 145.369 33.325 ;
			RECT	145.505 33.261 145.537 33.325 ;
			RECT	145.673 33.261 145.705 33.325 ;
			RECT	145.841 33.261 145.873 33.325 ;
			RECT	146.009 33.261 146.041 33.325 ;
			RECT	146.177 33.261 146.209 33.325 ;
			RECT	146.345 33.261 146.377 33.325 ;
			RECT	146.513 33.261 146.545 33.325 ;
			RECT	146.681 33.261 146.713 33.325 ;
			RECT	146.849 33.261 146.881 33.325 ;
			RECT	147.017 33.261 147.049 33.325 ;
			RECT	147.325 33.261 147.357 33.325 ;
			RECT	147.611 33.261 147.643 33.325 ;
			RECT	150.576 33.261 150.608 33.325 ;
			RECT	150.966 33.261 151.03 33.325 ;
			RECT	151.908 33.261 151.94 33.325 ;
			RECT	152.249 33.261 152.281 33.325 ;
			RECT	153.56 33.261 153.624 33.325 ;
			RECT	153.801 33.261 153.833 33.325 ;
			RECT	153.967 33.261 154.031 33.325 ;
			RECT	156.557 33.261 156.589 33.325 ;
			RECT	156.843 33.261 156.875 33.325 ;
			RECT	157.151 33.261 157.183 33.325 ;
			RECT	157.319 33.261 157.351 33.325 ;
			RECT	157.487 33.261 157.519 33.325 ;
			RECT	157.655 33.261 157.687 33.325 ;
			RECT	157.823 33.261 157.855 33.325 ;
			RECT	157.991 33.261 158.023 33.325 ;
			RECT	158.159 33.261 158.191 33.325 ;
			RECT	158.327 33.261 158.359 33.325 ;
			RECT	158.495 33.261 158.527 33.325 ;
			RECT	158.663 33.261 158.695 33.325 ;
			RECT	158.831 33.261 158.863 33.325 ;
			RECT	158.999 33.261 159.031 33.325 ;
			RECT	159.167 33.261 159.199 33.325 ;
			RECT	159.335 33.261 159.367 33.325 ;
			RECT	159.503 33.261 159.535 33.325 ;
			RECT	159.671 33.261 159.703 33.325 ;
			RECT	159.839 33.261 159.871 33.325 ;
			RECT	160.007 33.261 160.039 33.325 ;
			RECT	160.175 33.261 160.207 33.325 ;
			RECT	160.343 33.261 160.375 33.325 ;
			RECT	160.511 33.261 160.543 33.325 ;
			RECT	160.679 33.261 160.711 33.325 ;
			RECT	160.847 33.261 160.879 33.325 ;
			RECT	161.015 33.261 161.047 33.325 ;
			RECT	161.183 33.261 161.215 33.325 ;
			RECT	161.351 33.261 161.383 33.325 ;
			RECT	161.519 33.261 161.551 33.325 ;
			RECT	161.687 33.261 161.719 33.325 ;
			RECT	161.855 33.261 161.887 33.325 ;
			RECT	162.023 33.261 162.055 33.325 ;
			RECT	162.191 33.261 162.223 33.325 ;
			RECT	162.359 33.261 162.391 33.325 ;
			RECT	162.527 33.261 162.559 33.325 ;
			RECT	162.695 33.261 162.727 33.325 ;
			RECT	162.863 33.261 162.895 33.325 ;
			RECT	163.031 33.261 163.063 33.325 ;
			RECT	163.199 33.261 163.231 33.325 ;
			RECT	163.367 33.261 163.399 33.325 ;
			RECT	163.535 33.261 163.567 33.325 ;
			RECT	163.703 33.261 163.735 33.325 ;
			RECT	163.871 33.261 163.903 33.325 ;
			RECT	164.039 33.261 164.071 33.325 ;
			RECT	164.207 33.261 164.239 33.325 ;
			RECT	164.375 33.261 164.407 33.325 ;
			RECT	164.543 33.261 164.575 33.325 ;
			RECT	164.711 33.261 164.743 33.325 ;
			RECT	164.879 33.261 164.911 33.325 ;
			RECT	165.047 33.261 165.079 33.325 ;
			RECT	165.215 33.261 165.247 33.325 ;
			RECT	165.383 33.261 165.415 33.325 ;
			RECT	165.551 33.261 165.583 33.325 ;
			RECT	165.719 33.261 165.751 33.325 ;
			RECT	165.887 33.261 165.919 33.325 ;
			RECT	166.055 33.261 166.087 33.325 ;
			RECT	166.223 33.261 166.255 33.325 ;
			RECT	166.391 33.261 166.423 33.325 ;
			RECT	166.559 33.261 166.591 33.325 ;
			RECT	166.727 33.261 166.759 33.325 ;
			RECT	166.895 33.261 166.927 33.325 ;
			RECT	167.063 33.261 167.095 33.325 ;
			RECT	167.231 33.261 167.263 33.325 ;
			RECT	167.399 33.261 167.431 33.325 ;
			RECT	167.567 33.261 167.599 33.325 ;
			RECT	167.735 33.261 167.767 33.325 ;
			RECT	167.903 33.261 167.935 33.325 ;
			RECT	168.071 33.261 168.103 33.325 ;
			RECT	168.239 33.261 168.271 33.325 ;
			RECT	168.407 33.261 168.439 33.325 ;
			RECT	168.575 33.261 168.607 33.325 ;
			RECT	168.743 33.261 168.775 33.325 ;
			RECT	168.911 33.261 168.943 33.325 ;
			RECT	169.079 33.261 169.111 33.325 ;
			RECT	169.247 33.261 169.279 33.325 ;
			RECT	169.415 33.261 169.447 33.325 ;
			RECT	169.583 33.261 169.615 33.325 ;
			RECT	169.751 33.261 169.783 33.325 ;
			RECT	169.919 33.261 169.951 33.325 ;
			RECT	170.087 33.261 170.119 33.325 ;
			RECT	170.255 33.261 170.287 33.325 ;
			RECT	170.423 33.261 170.455 33.325 ;
			RECT	170.591 33.261 170.623 33.325 ;
			RECT	170.759 33.261 170.791 33.325 ;
			RECT	170.927 33.261 170.959 33.325 ;
			RECT	171.095 33.261 171.127 33.325 ;
			RECT	171.263 33.261 171.295 33.325 ;
			RECT	171.431 33.261 171.463 33.325 ;
			RECT	171.599 33.261 171.631 33.325 ;
			RECT	171.767 33.261 171.799 33.325 ;
			RECT	171.935 33.261 171.967 33.325 ;
			RECT	172.103 33.261 172.135 33.325 ;
			RECT	172.271 33.261 172.303 33.325 ;
			RECT	172.439 33.261 172.471 33.325 ;
			RECT	172.607 33.261 172.639 33.325 ;
			RECT	172.775 33.261 172.807 33.325 ;
			RECT	172.943 33.261 172.975 33.325 ;
			RECT	173.111 33.261 173.143 33.325 ;
			RECT	173.279 33.261 173.311 33.325 ;
			RECT	173.447 33.261 173.479 33.325 ;
			RECT	173.615 33.261 173.647 33.325 ;
			RECT	173.783 33.261 173.815 33.325 ;
			RECT	173.951 33.261 173.983 33.325 ;
			RECT	174.119 33.261 174.151 33.325 ;
			RECT	174.287 33.261 174.319 33.325 ;
			RECT	174.455 33.261 174.487 33.325 ;
			RECT	174.623 33.261 174.655 33.325 ;
			RECT	174.791 33.261 174.823 33.325 ;
			RECT	174.959 33.261 174.991 33.325 ;
			RECT	175.127 33.261 175.159 33.325 ;
			RECT	175.295 33.261 175.327 33.325 ;
			RECT	175.463 33.261 175.495 33.325 ;
			RECT	175.631 33.261 175.663 33.325 ;
			RECT	175.799 33.261 175.831 33.325 ;
			RECT	175.967 33.261 175.999 33.325 ;
			RECT	176.135 33.261 176.167 33.325 ;
			RECT	176.303 33.261 176.335 33.325 ;
			RECT	176.471 33.261 176.503 33.325 ;
			RECT	176.639 33.261 176.671 33.325 ;
			RECT	176.807 33.261 176.839 33.325 ;
			RECT	176.975 33.261 177.007 33.325 ;
			RECT	177.143 33.261 177.175 33.325 ;
			RECT	177.311 33.261 177.343 33.325 ;
			RECT	177.479 33.261 177.511 33.325 ;
			RECT	177.647 33.261 177.679 33.325 ;
			RECT	177.815 33.261 177.847 33.325 ;
			RECT	177.983 33.261 178.015 33.325 ;
			RECT	178.151 33.261 178.183 33.325 ;
			RECT	178.319 33.261 178.351 33.325 ;
			RECT	178.655 33.261 178.687 33.325 ;
			RECT	178.991 33.261 179.023 33.325 ;
			RECT	179.327 33.261 179.359 33.325 ;
			RECT	179.663 33.261 179.695 33.325 ;
			RECT	179.999 33.261 180.031 33.325 ;
			RECT	180.335 33.261 180.367 33.325 ;
			RECT	180.671 33.261 180.703 33.325 ;
			RECT	181.007 33.261 181.039 33.325 ;
			RECT	181.343 33.261 181.375 33.325 ;
			RECT	181.679 33.261 181.711 33.325 ;
			RECT	182.015 33.261 182.047 33.325 ;
			RECT	182.351 33.261 182.383 33.325 ;
			RECT	182.687 33.261 182.719 33.325 ;
			RECT	183.023 33.261 183.055 33.325 ;
			RECT	183.359 33.261 183.391 33.325 ;
			RECT	183.695 33.261 183.727 33.325 ;
			RECT	184.031 33.261 184.063 33.325 ;
			RECT	184.367 33.261 184.399 33.325 ;
			RECT	184.703 33.261 184.735 33.325 ;
			RECT	185.039 33.261 185.071 33.325 ;
			RECT	185.375 33.261 185.407 33.325 ;
			RECT	185.711 33.261 185.743 33.325 ;
			RECT	186.047 33.261 186.079 33.325 ;
			RECT	186.383 33.261 186.415 33.325 ;
			RECT	186.719 33.261 186.751 33.325 ;
			RECT	187.055 33.261 187.087 33.325 ;
			RECT	187.391 33.261 187.423 33.325 ;
			RECT	187.727 33.261 187.759 33.325 ;
			RECT	188.063 33.261 188.095 33.325 ;
			RECT	188.399 33.261 188.431 33.325 ;
			RECT	188.735 33.261 188.767 33.325 ;
			RECT	189.071 33.261 189.103 33.325 ;
			RECT	189.407 33.261 189.439 33.325 ;
			RECT	189.743 33.261 189.775 33.325 ;
			RECT	190.079 33.261 190.111 33.325 ;
			RECT	190.415 33.261 190.447 33.325 ;
			RECT	190.751 33.261 190.783 33.325 ;
			RECT	191.087 33.261 191.119 33.325 ;
			RECT	191.423 33.261 191.455 33.325 ;
			RECT	191.759 33.261 191.791 33.325 ;
			RECT	192.095 33.261 192.127 33.325 ;
			RECT	192.431 33.261 192.463 33.325 ;
			RECT	192.767 33.261 192.799 33.325 ;
			RECT	193.103 33.261 193.135 33.325 ;
			RECT	193.439 33.261 193.471 33.325 ;
			RECT	193.775 33.261 193.807 33.325 ;
			RECT	194.111 33.261 194.143 33.325 ;
			RECT	194.447 33.261 194.479 33.325 ;
			RECT	194.783 33.261 194.815 33.325 ;
			RECT	195.119 33.261 195.151 33.325 ;
			RECT	195.455 33.261 195.487 33.325 ;
			RECT	195.791 33.261 195.823 33.325 ;
			RECT	196.127 33.261 196.159 33.325 ;
			RECT	196.463 33.261 196.495 33.325 ;
			RECT	196.799 33.261 196.831 33.325 ;
			RECT	197.135 33.261 197.167 33.325 ;
			RECT	197.471 33.261 197.503 33.325 ;
			RECT	197.807 33.261 197.839 33.325 ;
			RECT	198.143 33.261 198.175 33.325 ;
			RECT	198.479 33.261 198.511 33.325 ;
			RECT	198.815 33.261 198.847 33.325 ;
			RECT	199.151 33.261 199.183 33.325 ;
			RECT	199.487 33.261 199.519 33.325 ;
			RECT	199.823 33.261 199.855 33.325 ;
			RECT	201.403 33.261 201.435 33.325 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 38.477 201.665 38.567 ;
			LAYER	J3 ;
			RECT	1.645 38.506 1.709 38.538 ;
			RECT	2.197 38.49 2.229 38.554 ;
			RECT	2.339 38.49 2.371 38.554 ;
			RECT	4.354 38.49 4.386 38.554 ;
			RECT	4.805 38.49 4.837 38.554 ;
			RECT	5.567 38.49 5.599 38.554 ;
			RECT	6.389 38.49 6.421 38.554 ;
			RECT	6.725 38.49 6.757 38.554 ;
			RECT	7.061 38.49 7.093 38.554 ;
			RECT	7.397 38.49 7.429 38.554 ;
			RECT	7.733 38.49 7.765 38.554 ;
			RECT	8.069 38.49 8.101 38.554 ;
			RECT	8.405 38.49 8.437 38.554 ;
			RECT	8.741 38.49 8.773 38.554 ;
			RECT	9.077 38.49 9.109 38.554 ;
			RECT	9.413 38.49 9.445 38.554 ;
			RECT	9.749 38.49 9.781 38.554 ;
			RECT	10.085 38.49 10.117 38.554 ;
			RECT	10.421 38.49 10.453 38.554 ;
			RECT	10.757 38.49 10.789 38.554 ;
			RECT	11.093 38.49 11.125 38.554 ;
			RECT	11.429 38.49 11.461 38.554 ;
			RECT	11.765 38.49 11.797 38.554 ;
			RECT	12.101 38.49 12.133 38.554 ;
			RECT	12.437 38.49 12.469 38.554 ;
			RECT	12.773 38.49 12.805 38.554 ;
			RECT	13.109 38.49 13.141 38.554 ;
			RECT	13.445 38.49 13.477 38.554 ;
			RECT	13.781 38.49 13.813 38.554 ;
			RECT	14.117 38.49 14.149 38.554 ;
			RECT	14.453 38.49 14.485 38.554 ;
			RECT	14.789 38.49 14.821 38.554 ;
			RECT	15.125 38.49 15.157 38.554 ;
			RECT	15.461 38.49 15.493 38.554 ;
			RECT	15.797 38.49 15.829 38.554 ;
			RECT	16.133 38.49 16.165 38.554 ;
			RECT	16.469 38.49 16.501 38.554 ;
			RECT	16.805 38.49 16.837 38.554 ;
			RECT	17.141 38.49 17.173 38.554 ;
			RECT	17.477 38.49 17.509 38.554 ;
			RECT	17.813 38.49 17.845 38.554 ;
			RECT	18.149 38.49 18.181 38.554 ;
			RECT	18.485 38.49 18.517 38.554 ;
			RECT	18.821 38.49 18.853 38.554 ;
			RECT	19.157 38.49 19.189 38.554 ;
			RECT	19.493 38.49 19.525 38.554 ;
			RECT	19.829 38.49 19.861 38.554 ;
			RECT	20.165 38.49 20.197 38.554 ;
			RECT	20.501 38.49 20.533 38.554 ;
			RECT	20.837 38.49 20.869 38.554 ;
			RECT	21.173 38.49 21.205 38.554 ;
			RECT	21.509 38.49 21.541 38.554 ;
			RECT	21.845 38.49 21.877 38.554 ;
			RECT	22.181 38.49 22.213 38.554 ;
			RECT	22.517 38.49 22.549 38.554 ;
			RECT	22.853 38.49 22.885 38.554 ;
			RECT	23.189 38.49 23.221 38.554 ;
			RECT	23.525 38.49 23.557 38.554 ;
			RECT	23.861 38.49 23.893 38.554 ;
			RECT	24.197 38.49 24.229 38.554 ;
			RECT	24.533 38.49 24.565 38.554 ;
			RECT	24.869 38.49 24.901 38.554 ;
			RECT	25.205 38.49 25.237 38.554 ;
			RECT	25.541 38.49 25.573 38.554 ;
			RECT	25.877 38.49 25.909 38.554 ;
			RECT	26.213 38.49 26.245 38.554 ;
			RECT	26.549 38.49 26.581 38.554 ;
			RECT	26.885 38.49 26.917 38.554 ;
			RECT	27.221 38.49 27.253 38.554 ;
			RECT	27.557 38.49 27.589 38.554 ;
			RECT	28.224 38.49 28.256 38.554 ;
			RECT	28.896 38.49 28.928 38.554 ;
			RECT	29.568 38.49 29.6 38.554 ;
			RECT	30.24 38.49 30.272 38.554 ;
			RECT	30.576 38.49 30.608 38.554 ;
			RECT	31.248 38.49 31.28 38.554 ;
			RECT	31.92 38.49 31.952 38.554 ;
			RECT	32.256 38.49 32.288 38.554 ;
			RECT	32.592 38.49 32.624 38.554 ;
			RECT	32.928 38.49 32.96 38.554 ;
			RECT	33.264 38.49 33.296 38.554 ;
			RECT	33.6 38.49 33.632 38.554 ;
			RECT	33.926 38.49 33.958 38.554 ;
			RECT	34.272 38.49 34.304 38.554 ;
			RECT	35.28 38.49 35.312 38.554 ;
			RECT	35.952 38.49 35.984 38.554 ;
			RECT	37.296 38.49 37.328 38.554 ;
			RECT	37.632 38.49 37.664 38.554 ;
			RECT	38.64 38.49 38.672 38.554 ;
			RECT	39.648 38.49 39.68 38.554 ;
			RECT	41.328 38.49 41.36 38.554 ;
			RECT	42 38.49 42.032 38.554 ;
			RECT	42.336 38.49 42.368 38.554 ;
			RECT	42.672 38.49 42.704 38.554 ;
			RECT	43.008 38.49 43.04 38.554 ;
			RECT	43.68 38.49 43.712 38.554 ;
			RECT	44.016 38.49 44.048 38.554 ;
			RECT	44.688 38.49 44.72 38.554 ;
			RECT	45.696 38.49 45.728 38.554 ;
			RECT	46.368 38.49 46.4 38.554 ;
			RECT	47.04 38.49 47.072 38.554 ;
			RECT	48.384 38.49 48.416 38.554 ;
			RECT	48.536 38.49 48.568 38.554 ;
			RECT	49.091 38.49 49.123 38.554 ;
			RECT	49.327 38.49 49.359 38.554 ;
			RECT	51.92 38.49 51.952 38.554 ;
			RECT	52.968 38.506 53.032 38.538 ;
			RECT	53.878 38.506 53.942 38.538 ;
			RECT	54.804 38.49 54.836 38.554 ;
			RECT	55.53 38.49 55.562 38.554 ;
			RECT	55.969 38.506 56.033 38.538 ;
			RECT	57.18 38.49 57.212 38.554 ;
			RECT	57.363 38.49 57.395 38.554 ;
			RECT	58.845 38.49 58.877 38.554 ;
			RECT	59.081 38.49 59.113 38.554 ;
			RECT	59.636 38.49 59.668 38.554 ;
			RECT	59.788 38.49 59.82 38.554 ;
			RECT	61.132 38.49 61.164 38.554 ;
			RECT	61.804 38.49 61.836 38.554 ;
			RECT	62.476 38.49 62.508 38.554 ;
			RECT	63.484 38.49 63.516 38.554 ;
			RECT	64.156 38.49 64.188 38.554 ;
			RECT	64.492 38.49 64.524 38.554 ;
			RECT	65.164 38.49 65.196 38.554 ;
			RECT	65.5 38.49 65.532 38.554 ;
			RECT	65.836 38.49 65.868 38.554 ;
			RECT	66.172 38.49 66.204 38.554 ;
			RECT	66.844 38.49 66.876 38.554 ;
			RECT	68.524 38.49 68.556 38.554 ;
			RECT	69.532 38.49 69.564 38.554 ;
			RECT	70.54 38.49 70.572 38.554 ;
			RECT	70.876 38.49 70.908 38.554 ;
			RECT	72.22 38.49 72.252 38.554 ;
			RECT	72.892 38.49 72.924 38.554 ;
			RECT	73.9 38.49 73.932 38.554 ;
			RECT	74.246 38.49 74.278 38.554 ;
			RECT	74.572 38.49 74.604 38.554 ;
			RECT	74.908 38.49 74.94 38.554 ;
			RECT	75.244 38.49 75.276 38.554 ;
			RECT	75.58 38.49 75.612 38.554 ;
			RECT	75.916 38.49 75.948 38.554 ;
			RECT	76.252 38.49 76.284 38.554 ;
			RECT	76.924 38.49 76.956 38.554 ;
			RECT	77.596 38.49 77.628 38.554 ;
			RECT	77.932 38.49 77.964 38.554 ;
			RECT	78.604 38.49 78.636 38.554 ;
			RECT	79.276 38.49 79.308 38.554 ;
			RECT	79.948 38.49 79.98 38.554 ;
			RECT	80.615 38.49 80.647 38.554 ;
			RECT	80.951 38.49 80.983 38.554 ;
			RECT	81.287 38.49 81.319 38.554 ;
			RECT	81.623 38.49 81.655 38.554 ;
			RECT	81.959 38.49 81.991 38.554 ;
			RECT	82.295 38.49 82.327 38.554 ;
			RECT	82.631 38.49 82.663 38.554 ;
			RECT	82.967 38.49 82.999 38.554 ;
			RECT	83.303 38.49 83.335 38.554 ;
			RECT	83.639 38.49 83.671 38.554 ;
			RECT	83.975 38.49 84.007 38.554 ;
			RECT	84.311 38.49 84.343 38.554 ;
			RECT	84.647 38.49 84.679 38.554 ;
			RECT	84.983 38.49 85.015 38.554 ;
			RECT	85.319 38.49 85.351 38.554 ;
			RECT	85.655 38.49 85.687 38.554 ;
			RECT	85.991 38.49 86.023 38.554 ;
			RECT	86.327 38.49 86.359 38.554 ;
			RECT	86.663 38.49 86.695 38.554 ;
			RECT	86.999 38.49 87.031 38.554 ;
			RECT	87.335 38.49 87.367 38.554 ;
			RECT	87.671 38.49 87.703 38.554 ;
			RECT	88.007 38.49 88.039 38.554 ;
			RECT	88.343 38.49 88.375 38.554 ;
			RECT	88.679 38.49 88.711 38.554 ;
			RECT	89.015 38.49 89.047 38.554 ;
			RECT	89.351 38.49 89.383 38.554 ;
			RECT	89.687 38.49 89.719 38.554 ;
			RECT	90.023 38.49 90.055 38.554 ;
			RECT	90.359 38.49 90.391 38.554 ;
			RECT	90.695 38.49 90.727 38.554 ;
			RECT	91.031 38.49 91.063 38.554 ;
			RECT	91.367 38.49 91.399 38.554 ;
			RECT	91.703 38.49 91.735 38.554 ;
			RECT	92.039 38.49 92.071 38.554 ;
			RECT	92.375 38.49 92.407 38.554 ;
			RECT	92.711 38.49 92.743 38.554 ;
			RECT	93.047 38.49 93.079 38.554 ;
			RECT	93.383 38.49 93.415 38.554 ;
			RECT	93.719 38.49 93.751 38.554 ;
			RECT	94.055 38.49 94.087 38.554 ;
			RECT	94.391 38.49 94.423 38.554 ;
			RECT	94.727 38.49 94.759 38.554 ;
			RECT	95.063 38.49 95.095 38.554 ;
			RECT	95.399 38.49 95.431 38.554 ;
			RECT	95.735 38.49 95.767 38.554 ;
			RECT	96.071 38.49 96.103 38.554 ;
			RECT	96.407 38.49 96.439 38.554 ;
			RECT	96.743 38.49 96.775 38.554 ;
			RECT	97.079 38.49 97.111 38.554 ;
			RECT	97.415 38.49 97.447 38.554 ;
			RECT	97.751 38.49 97.783 38.554 ;
			RECT	98.087 38.49 98.119 38.554 ;
			RECT	98.423 38.49 98.455 38.554 ;
			RECT	98.759 38.49 98.791 38.554 ;
			RECT	99.095 38.49 99.127 38.554 ;
			RECT	99.431 38.49 99.463 38.554 ;
			RECT	99.767 38.49 99.799 38.554 ;
			RECT	100.103 38.49 100.135 38.554 ;
			RECT	100.439 38.49 100.471 38.554 ;
			RECT	100.775 38.49 100.807 38.554 ;
			RECT	101.111 38.49 101.143 38.554 ;
			RECT	101.447 38.49 101.479 38.554 ;
			RECT	101.783 38.49 101.815 38.554 ;
			RECT	102.605 38.49 102.637 38.554 ;
			RECT	102.995 38.49 103.027 38.554 ;
			RECT	103.175 38.49 103.207 38.554 ;
			RECT	103.565 38.49 103.597 38.554 ;
			RECT	104.387 38.49 104.419 38.554 ;
			RECT	104.723 38.49 104.755 38.554 ;
			RECT	105.059 38.49 105.091 38.554 ;
			RECT	105.395 38.49 105.427 38.554 ;
			RECT	105.731 38.49 105.763 38.554 ;
			RECT	106.067 38.49 106.099 38.554 ;
			RECT	106.403 38.49 106.435 38.554 ;
			RECT	106.739 38.49 106.771 38.554 ;
			RECT	107.075 38.49 107.107 38.554 ;
			RECT	107.411 38.49 107.443 38.554 ;
			RECT	107.747 38.49 107.779 38.554 ;
			RECT	108.083 38.49 108.115 38.554 ;
			RECT	108.419 38.49 108.451 38.554 ;
			RECT	108.755 38.49 108.787 38.554 ;
			RECT	109.091 38.49 109.123 38.554 ;
			RECT	109.427 38.49 109.459 38.554 ;
			RECT	109.763 38.49 109.795 38.554 ;
			RECT	110.099 38.49 110.131 38.554 ;
			RECT	110.435 38.49 110.467 38.554 ;
			RECT	110.771 38.49 110.803 38.554 ;
			RECT	111.107 38.49 111.139 38.554 ;
			RECT	111.443 38.49 111.475 38.554 ;
			RECT	111.779 38.49 111.811 38.554 ;
			RECT	112.115 38.49 112.147 38.554 ;
			RECT	112.451 38.49 112.483 38.554 ;
			RECT	112.787 38.49 112.819 38.554 ;
			RECT	113.123 38.49 113.155 38.554 ;
			RECT	113.459 38.49 113.491 38.554 ;
			RECT	113.795 38.49 113.827 38.554 ;
			RECT	114.131 38.49 114.163 38.554 ;
			RECT	114.467 38.49 114.499 38.554 ;
			RECT	114.803 38.49 114.835 38.554 ;
			RECT	115.139 38.49 115.171 38.554 ;
			RECT	115.475 38.49 115.507 38.554 ;
			RECT	115.811 38.49 115.843 38.554 ;
			RECT	116.147 38.49 116.179 38.554 ;
			RECT	116.483 38.49 116.515 38.554 ;
			RECT	116.819 38.49 116.851 38.554 ;
			RECT	117.155 38.49 117.187 38.554 ;
			RECT	117.491 38.49 117.523 38.554 ;
			RECT	117.827 38.49 117.859 38.554 ;
			RECT	118.163 38.49 118.195 38.554 ;
			RECT	118.499 38.49 118.531 38.554 ;
			RECT	118.835 38.49 118.867 38.554 ;
			RECT	119.171 38.49 119.203 38.554 ;
			RECT	119.507 38.49 119.539 38.554 ;
			RECT	119.843 38.49 119.875 38.554 ;
			RECT	120.179 38.49 120.211 38.554 ;
			RECT	120.515 38.49 120.547 38.554 ;
			RECT	120.851 38.49 120.883 38.554 ;
			RECT	121.187 38.49 121.219 38.554 ;
			RECT	121.523 38.49 121.555 38.554 ;
			RECT	121.859 38.49 121.891 38.554 ;
			RECT	122.195 38.49 122.227 38.554 ;
			RECT	122.531 38.49 122.563 38.554 ;
			RECT	122.867 38.49 122.899 38.554 ;
			RECT	123.203 38.49 123.235 38.554 ;
			RECT	123.539 38.49 123.571 38.554 ;
			RECT	123.875 38.49 123.907 38.554 ;
			RECT	124.211 38.49 124.243 38.554 ;
			RECT	124.547 38.49 124.579 38.554 ;
			RECT	124.883 38.49 124.915 38.554 ;
			RECT	125.219 38.49 125.251 38.554 ;
			RECT	125.555 38.49 125.587 38.554 ;
			RECT	126.222 38.49 126.254 38.554 ;
			RECT	126.894 38.49 126.926 38.554 ;
			RECT	127.566 38.49 127.598 38.554 ;
			RECT	128.238 38.49 128.27 38.554 ;
			RECT	128.574 38.49 128.606 38.554 ;
			RECT	129.246 38.49 129.278 38.554 ;
			RECT	129.918 38.49 129.95 38.554 ;
			RECT	130.254 38.49 130.286 38.554 ;
			RECT	130.59 38.49 130.622 38.554 ;
			RECT	130.926 38.49 130.958 38.554 ;
			RECT	131.262 38.49 131.294 38.554 ;
			RECT	131.598 38.49 131.63 38.554 ;
			RECT	131.924 38.49 131.956 38.554 ;
			RECT	132.27 38.49 132.302 38.554 ;
			RECT	133.278 38.49 133.31 38.554 ;
			RECT	133.95 38.49 133.982 38.554 ;
			RECT	135.294 38.49 135.326 38.554 ;
			RECT	135.63 38.49 135.662 38.554 ;
			RECT	136.638 38.49 136.67 38.554 ;
			RECT	137.646 38.49 137.678 38.554 ;
			RECT	139.326 38.49 139.358 38.554 ;
			RECT	139.998 38.49 140.03 38.554 ;
			RECT	140.334 38.49 140.366 38.554 ;
			RECT	140.67 38.49 140.702 38.554 ;
			RECT	141.006 38.49 141.038 38.554 ;
			RECT	141.678 38.49 141.71 38.554 ;
			RECT	142.014 38.49 142.046 38.554 ;
			RECT	142.686 38.49 142.718 38.554 ;
			RECT	143.694 38.49 143.726 38.554 ;
			RECT	144.366 38.49 144.398 38.554 ;
			RECT	145.038 38.49 145.07 38.554 ;
			RECT	146.382 38.49 146.414 38.554 ;
			RECT	146.534 38.49 146.566 38.554 ;
			RECT	147.089 38.49 147.121 38.554 ;
			RECT	147.325 38.49 147.357 38.554 ;
			RECT	149.918 38.49 149.95 38.554 ;
			RECT	150.966 38.506 151.03 38.538 ;
			RECT	151.876 38.506 151.94 38.538 ;
			RECT	152.802 38.49 152.834 38.554 ;
			RECT	153.528 38.49 153.56 38.554 ;
			RECT	153.967 38.506 154.031 38.538 ;
			RECT	155.178 38.49 155.21 38.554 ;
			RECT	155.361 38.49 155.393 38.554 ;
			RECT	156.843 38.49 156.875 38.554 ;
			RECT	157.079 38.49 157.111 38.554 ;
			RECT	157.634 38.49 157.666 38.554 ;
			RECT	157.786 38.49 157.818 38.554 ;
			RECT	159.13 38.49 159.162 38.554 ;
			RECT	159.802 38.49 159.834 38.554 ;
			RECT	160.474 38.49 160.506 38.554 ;
			RECT	161.482 38.49 161.514 38.554 ;
			RECT	162.154 38.49 162.186 38.554 ;
			RECT	162.49 38.49 162.522 38.554 ;
			RECT	163.162 38.49 163.194 38.554 ;
			RECT	163.498 38.49 163.53 38.554 ;
			RECT	163.834 38.49 163.866 38.554 ;
			RECT	164.17 38.49 164.202 38.554 ;
			RECT	164.842 38.49 164.874 38.554 ;
			RECT	166.522 38.49 166.554 38.554 ;
			RECT	167.53 38.49 167.562 38.554 ;
			RECT	168.538 38.49 168.57 38.554 ;
			RECT	168.874 38.49 168.906 38.554 ;
			RECT	170.218 38.49 170.25 38.554 ;
			RECT	170.89 38.49 170.922 38.554 ;
			RECT	171.898 38.49 171.93 38.554 ;
			RECT	172.244 38.49 172.276 38.554 ;
			RECT	172.57 38.49 172.602 38.554 ;
			RECT	172.906 38.49 172.938 38.554 ;
			RECT	173.242 38.49 173.274 38.554 ;
			RECT	173.578 38.49 173.61 38.554 ;
			RECT	173.914 38.49 173.946 38.554 ;
			RECT	174.25 38.49 174.282 38.554 ;
			RECT	174.922 38.49 174.954 38.554 ;
			RECT	175.594 38.49 175.626 38.554 ;
			RECT	175.93 38.49 175.962 38.554 ;
			RECT	176.602 38.49 176.634 38.554 ;
			RECT	177.274 38.49 177.306 38.554 ;
			RECT	177.946 38.49 177.978 38.554 ;
			RECT	178.613 38.49 178.645 38.554 ;
			RECT	178.949 38.49 178.981 38.554 ;
			RECT	179.285 38.49 179.317 38.554 ;
			RECT	179.621 38.49 179.653 38.554 ;
			RECT	179.957 38.49 179.989 38.554 ;
			RECT	180.293 38.49 180.325 38.554 ;
			RECT	180.629 38.49 180.661 38.554 ;
			RECT	180.965 38.49 180.997 38.554 ;
			RECT	181.301 38.49 181.333 38.554 ;
			RECT	181.637 38.49 181.669 38.554 ;
			RECT	181.973 38.49 182.005 38.554 ;
			RECT	182.309 38.49 182.341 38.554 ;
			RECT	182.645 38.49 182.677 38.554 ;
			RECT	182.981 38.49 183.013 38.554 ;
			RECT	183.317 38.49 183.349 38.554 ;
			RECT	183.653 38.49 183.685 38.554 ;
			RECT	183.989 38.49 184.021 38.554 ;
			RECT	184.325 38.49 184.357 38.554 ;
			RECT	184.661 38.49 184.693 38.554 ;
			RECT	184.997 38.49 185.029 38.554 ;
			RECT	185.333 38.49 185.365 38.554 ;
			RECT	185.669 38.49 185.701 38.554 ;
			RECT	186.005 38.49 186.037 38.554 ;
			RECT	186.341 38.49 186.373 38.554 ;
			RECT	186.677 38.49 186.709 38.554 ;
			RECT	187.013 38.49 187.045 38.554 ;
			RECT	187.349 38.49 187.381 38.554 ;
			RECT	187.685 38.49 187.717 38.554 ;
			RECT	188.021 38.49 188.053 38.554 ;
			RECT	188.357 38.49 188.389 38.554 ;
			RECT	188.693 38.49 188.725 38.554 ;
			RECT	189.029 38.49 189.061 38.554 ;
			RECT	189.365 38.49 189.397 38.554 ;
			RECT	189.701 38.49 189.733 38.554 ;
			RECT	190.037 38.49 190.069 38.554 ;
			RECT	190.373 38.49 190.405 38.554 ;
			RECT	190.709 38.49 190.741 38.554 ;
			RECT	191.045 38.49 191.077 38.554 ;
			RECT	191.381 38.49 191.413 38.554 ;
			RECT	191.717 38.49 191.749 38.554 ;
			RECT	192.053 38.49 192.085 38.554 ;
			RECT	192.389 38.49 192.421 38.554 ;
			RECT	192.725 38.49 192.757 38.554 ;
			RECT	193.061 38.49 193.093 38.554 ;
			RECT	193.397 38.49 193.429 38.554 ;
			RECT	193.733 38.49 193.765 38.554 ;
			RECT	194.069 38.49 194.101 38.554 ;
			RECT	194.405 38.49 194.437 38.554 ;
			RECT	194.741 38.49 194.773 38.554 ;
			RECT	195.077 38.49 195.109 38.554 ;
			RECT	195.413 38.49 195.445 38.554 ;
			RECT	195.749 38.49 195.781 38.554 ;
			RECT	196.085 38.49 196.117 38.554 ;
			RECT	196.421 38.49 196.453 38.554 ;
			RECT	196.757 38.49 196.789 38.554 ;
			RECT	197.093 38.49 197.125 38.554 ;
			RECT	197.429 38.49 197.461 38.554 ;
			RECT	197.765 38.49 197.797 38.554 ;
			RECT	198.101 38.49 198.133 38.554 ;
			RECT	198.437 38.49 198.469 38.554 ;
			RECT	198.773 38.49 198.805 38.554 ;
			RECT	199.109 38.49 199.141 38.554 ;
			RECT	199.445 38.49 199.477 38.554 ;
			RECT	199.781 38.49 199.813 38.554 ;
			RECT	200.603 38.49 200.635 38.554 ;
			RECT	201.403 38.49 201.435 38.554 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 40.729 201.665 40.819 ;
			LAYER	J3 ;
			RECT	1.164 40.742 1.196 40.806 ;
			RECT	1.645 40.758 1.709 40.79 ;
			RECT	2.197 40.758 2.229 40.79 ;
			RECT	2.339 40.758 2.371 40.79 ;
			RECT	3.438 40.742 3.47 40.806 ;
			RECT	4.354 40.758 4.386 40.79 ;
			RECT	4.554 40.742 4.586 40.806 ;
			RECT	5.567 40.742 5.599 40.806 ;
			RECT	5.758 40.742 5.79 40.806 ;
			RECT	6.389 40.742 6.421 40.806 ;
			RECT	6.725 40.742 6.757 40.806 ;
			RECT	7.061 40.742 7.093 40.806 ;
			RECT	7.397 40.742 7.429 40.806 ;
			RECT	7.733 40.742 7.765 40.806 ;
			RECT	8.069 40.742 8.101 40.806 ;
			RECT	8.405 40.742 8.437 40.806 ;
			RECT	8.741 40.742 8.773 40.806 ;
			RECT	9.077 40.742 9.109 40.806 ;
			RECT	9.413 40.742 9.445 40.806 ;
			RECT	9.749 40.742 9.781 40.806 ;
			RECT	10.085 40.742 10.117 40.806 ;
			RECT	10.421 40.742 10.453 40.806 ;
			RECT	10.757 40.742 10.789 40.806 ;
			RECT	11.093 40.742 11.125 40.806 ;
			RECT	11.429 40.742 11.461 40.806 ;
			RECT	11.765 40.742 11.797 40.806 ;
			RECT	12.101 40.742 12.133 40.806 ;
			RECT	12.437 40.742 12.469 40.806 ;
			RECT	12.773 40.742 12.805 40.806 ;
			RECT	13.109 40.742 13.141 40.806 ;
			RECT	13.445 40.742 13.477 40.806 ;
			RECT	13.781 40.742 13.813 40.806 ;
			RECT	14.117 40.742 14.149 40.806 ;
			RECT	14.453 40.742 14.485 40.806 ;
			RECT	14.789 40.742 14.821 40.806 ;
			RECT	15.125 40.742 15.157 40.806 ;
			RECT	15.461 40.742 15.493 40.806 ;
			RECT	15.797 40.742 15.829 40.806 ;
			RECT	16.133 40.742 16.165 40.806 ;
			RECT	16.469 40.742 16.501 40.806 ;
			RECT	16.805 40.742 16.837 40.806 ;
			RECT	17.141 40.742 17.173 40.806 ;
			RECT	17.477 40.742 17.509 40.806 ;
			RECT	17.813 40.742 17.845 40.806 ;
			RECT	18.149 40.742 18.181 40.806 ;
			RECT	18.485 40.742 18.517 40.806 ;
			RECT	18.821 40.742 18.853 40.806 ;
			RECT	19.157 40.742 19.189 40.806 ;
			RECT	19.493 40.742 19.525 40.806 ;
			RECT	19.829 40.742 19.861 40.806 ;
			RECT	20.165 40.742 20.197 40.806 ;
			RECT	20.501 40.742 20.533 40.806 ;
			RECT	20.837 40.742 20.869 40.806 ;
			RECT	21.173 40.742 21.205 40.806 ;
			RECT	21.509 40.742 21.541 40.806 ;
			RECT	21.845 40.742 21.877 40.806 ;
			RECT	22.181 40.742 22.213 40.806 ;
			RECT	22.517 40.742 22.549 40.806 ;
			RECT	22.853 40.742 22.885 40.806 ;
			RECT	23.189 40.742 23.221 40.806 ;
			RECT	23.525 40.742 23.557 40.806 ;
			RECT	23.861 40.742 23.893 40.806 ;
			RECT	24.197 40.742 24.229 40.806 ;
			RECT	24.533 40.742 24.565 40.806 ;
			RECT	24.869 40.742 24.901 40.806 ;
			RECT	25.205 40.742 25.237 40.806 ;
			RECT	25.541 40.742 25.573 40.806 ;
			RECT	25.877 40.742 25.909 40.806 ;
			RECT	26.213 40.742 26.245 40.806 ;
			RECT	26.549 40.742 26.581 40.806 ;
			RECT	26.885 40.742 26.917 40.806 ;
			RECT	27.221 40.742 27.253 40.806 ;
			RECT	27.557 40.742 27.589 40.806 ;
			RECT	28.224 40.742 28.256 40.806 ;
			RECT	28.56 40.742 28.592 40.806 ;
			RECT	28.896 40.742 28.928 40.806 ;
			RECT	29.232 40.742 29.264 40.806 ;
			RECT	29.568 40.742 29.6 40.806 ;
			RECT	29.904 40.742 29.936 40.806 ;
			RECT	30.24 40.742 30.272 40.806 ;
			RECT	30.576 40.742 30.608 40.806 ;
			RECT	30.912 40.742 30.944 40.806 ;
			RECT	31.248 40.742 31.28 40.806 ;
			RECT	31.584 40.742 31.616 40.806 ;
			RECT	31.92 40.742 31.952 40.806 ;
			RECT	32.256 40.742 32.288 40.806 ;
			RECT	32.592 40.742 32.624 40.806 ;
			RECT	32.928 40.742 32.96 40.806 ;
			RECT	33.264 40.742 33.296 40.806 ;
			RECT	33.6 40.742 33.632 40.806 ;
			RECT	33.936 40.742 33.968 40.806 ;
			RECT	34.272 40.742 34.304 40.806 ;
			RECT	34.608 40.742 34.64 40.806 ;
			RECT	34.944 40.742 34.976 40.806 ;
			RECT	35.28 40.742 35.312 40.806 ;
			RECT	35.616 40.742 35.648 40.806 ;
			RECT	35.952 40.742 35.984 40.806 ;
			RECT	36.288 40.742 36.32 40.806 ;
			RECT	36.624 40.742 36.656 40.806 ;
			RECT	36.96 40.742 36.992 40.806 ;
			RECT	37.296 40.742 37.328 40.806 ;
			RECT	37.632 40.742 37.664 40.806 ;
			RECT	37.968 40.742 38 40.806 ;
			RECT	38.64 40.742 38.672 40.806 ;
			RECT	38.976 40.742 39.008 40.806 ;
			RECT	39.648 40.742 39.68 40.806 ;
			RECT	39.984 40.742 40.016 40.806 ;
			RECT	40.32 40.742 40.352 40.806 ;
			RECT	40.656 40.742 40.688 40.806 ;
			RECT	40.992 40.742 41.024 40.806 ;
			RECT	41.328 40.742 41.36 40.806 ;
			RECT	41.664 40.742 41.696 40.806 ;
			RECT	42 40.742 42.032 40.806 ;
			RECT	42.336 40.742 42.368 40.806 ;
			RECT	42.672 40.742 42.704 40.806 ;
			RECT	43.008 40.742 43.04 40.806 ;
			RECT	43.344 40.742 43.376 40.806 ;
			RECT	43.68 40.742 43.712 40.806 ;
			RECT	44.016 40.742 44.048 40.806 ;
			RECT	44.352 40.742 44.384 40.806 ;
			RECT	44.688 40.742 44.72 40.806 ;
			RECT	45.024 40.742 45.056 40.806 ;
			RECT	45.696 40.742 45.728 40.806 ;
			RECT	46.032 40.742 46.064 40.806 ;
			RECT	46.368 40.742 46.4 40.806 ;
			RECT	46.704 40.742 46.736 40.806 ;
			RECT	47.04 40.742 47.072 40.806 ;
			RECT	47.376 40.742 47.408 40.806 ;
			RECT	47.712 40.742 47.744 40.806 ;
			RECT	48.384 40.742 48.416 40.806 ;
			RECT	49.091 40.742 49.123 40.806 ;
			RECT	49.327 40.742 49.359 40.806 ;
			RECT	49.711 40.742 49.743 40.806 ;
			RECT	50.33 40.742 50.362 40.806 ;
			RECT	50.648 40.742 50.68 40.806 ;
			RECT	51.92 40.742 51.952 40.806 ;
			RECT	52.968 40.758 53.032 40.79 ;
			RECT	53.91 40.742 53.942 40.806 ;
			RECT	54.363 40.758 54.427 40.79 ;
			RECT	54.804 40.742 54.836 40.806 ;
			RECT	55.562 40.758 55.626 40.79 ;
			RECT	55.969 40.758 56.033 40.79 ;
			RECT	57.363 40.742 57.395 40.806 ;
			RECT	58.461 40.742 58.493 40.806 ;
			RECT	58.845 40.742 58.877 40.806 ;
			RECT	59.081 40.742 59.113 40.806 ;
			RECT	59.788 40.742 59.82 40.806 ;
			RECT	60.46 40.742 60.492 40.806 ;
			RECT	60.796 40.742 60.828 40.806 ;
			RECT	61.132 40.742 61.164 40.806 ;
			RECT	61.468 40.742 61.5 40.806 ;
			RECT	61.804 40.742 61.836 40.806 ;
			RECT	62.14 40.742 62.172 40.806 ;
			RECT	62.476 40.742 62.508 40.806 ;
			RECT	63.148 40.742 63.18 40.806 ;
			RECT	63.484 40.742 63.516 40.806 ;
			RECT	63.82 40.742 63.852 40.806 ;
			RECT	64.156 40.742 64.188 40.806 ;
			RECT	64.492 40.742 64.524 40.806 ;
			RECT	64.828 40.742 64.86 40.806 ;
			RECT	65.164 40.742 65.196 40.806 ;
			RECT	65.5 40.742 65.532 40.806 ;
			RECT	65.836 40.742 65.868 40.806 ;
			RECT	66.172 40.742 66.204 40.806 ;
			RECT	66.508 40.742 66.54 40.806 ;
			RECT	66.844 40.742 66.876 40.806 ;
			RECT	67.18 40.742 67.212 40.806 ;
			RECT	67.516 40.742 67.548 40.806 ;
			RECT	67.852 40.742 67.884 40.806 ;
			RECT	68.188 40.742 68.22 40.806 ;
			RECT	68.524 40.742 68.556 40.806 ;
			RECT	69.196 40.742 69.228 40.806 ;
			RECT	69.532 40.742 69.564 40.806 ;
			RECT	70.204 40.742 70.236 40.806 ;
			RECT	70.54 40.742 70.572 40.806 ;
			RECT	70.876 40.742 70.908 40.806 ;
			RECT	71.212 40.742 71.244 40.806 ;
			RECT	71.548 40.742 71.58 40.806 ;
			RECT	71.884 40.742 71.916 40.806 ;
			RECT	72.22 40.742 72.252 40.806 ;
			RECT	72.556 40.742 72.588 40.806 ;
			RECT	72.892 40.742 72.924 40.806 ;
			RECT	73.228 40.742 73.26 40.806 ;
			RECT	73.564 40.742 73.596 40.806 ;
			RECT	73.9 40.742 73.932 40.806 ;
			RECT	74.236 40.742 74.268 40.806 ;
			RECT	74.572 40.742 74.604 40.806 ;
			RECT	74.908 40.742 74.94 40.806 ;
			RECT	75.244 40.742 75.276 40.806 ;
			RECT	75.58 40.742 75.612 40.806 ;
			RECT	75.916 40.742 75.948 40.806 ;
			RECT	76.252 40.742 76.284 40.806 ;
			RECT	76.588 40.742 76.62 40.806 ;
			RECT	76.924 40.742 76.956 40.806 ;
			RECT	77.26 40.742 77.292 40.806 ;
			RECT	77.596 40.742 77.628 40.806 ;
			RECT	77.932 40.742 77.964 40.806 ;
			RECT	78.268 40.742 78.3 40.806 ;
			RECT	78.604 40.742 78.636 40.806 ;
			RECT	78.94 40.742 78.972 40.806 ;
			RECT	79.276 40.742 79.308 40.806 ;
			RECT	79.612 40.742 79.644 40.806 ;
			RECT	79.948 40.742 79.98 40.806 ;
			RECT	80.615 40.742 80.647 40.806 ;
			RECT	80.951 40.742 80.983 40.806 ;
			RECT	81.287 40.742 81.319 40.806 ;
			RECT	81.623 40.742 81.655 40.806 ;
			RECT	81.959 40.742 81.991 40.806 ;
			RECT	82.295 40.742 82.327 40.806 ;
			RECT	82.631 40.742 82.663 40.806 ;
			RECT	82.967 40.742 82.999 40.806 ;
			RECT	83.303 40.742 83.335 40.806 ;
			RECT	83.639 40.742 83.671 40.806 ;
			RECT	83.975 40.742 84.007 40.806 ;
			RECT	84.311 40.742 84.343 40.806 ;
			RECT	84.647 40.742 84.679 40.806 ;
			RECT	84.983 40.742 85.015 40.806 ;
			RECT	85.319 40.742 85.351 40.806 ;
			RECT	85.655 40.742 85.687 40.806 ;
			RECT	85.991 40.742 86.023 40.806 ;
			RECT	86.327 40.742 86.359 40.806 ;
			RECT	86.663 40.742 86.695 40.806 ;
			RECT	86.999 40.742 87.031 40.806 ;
			RECT	87.335 40.742 87.367 40.806 ;
			RECT	87.671 40.742 87.703 40.806 ;
			RECT	88.007 40.742 88.039 40.806 ;
			RECT	88.343 40.742 88.375 40.806 ;
			RECT	88.679 40.742 88.711 40.806 ;
			RECT	89.015 40.742 89.047 40.806 ;
			RECT	89.351 40.742 89.383 40.806 ;
			RECT	89.687 40.742 89.719 40.806 ;
			RECT	90.023 40.742 90.055 40.806 ;
			RECT	90.359 40.742 90.391 40.806 ;
			RECT	90.695 40.742 90.727 40.806 ;
			RECT	91.031 40.742 91.063 40.806 ;
			RECT	91.367 40.742 91.399 40.806 ;
			RECT	91.703 40.742 91.735 40.806 ;
			RECT	92.039 40.742 92.071 40.806 ;
			RECT	92.375 40.742 92.407 40.806 ;
			RECT	92.711 40.742 92.743 40.806 ;
			RECT	93.047 40.742 93.079 40.806 ;
			RECT	93.383 40.742 93.415 40.806 ;
			RECT	93.719 40.742 93.751 40.806 ;
			RECT	94.055 40.742 94.087 40.806 ;
			RECT	94.391 40.742 94.423 40.806 ;
			RECT	94.727 40.742 94.759 40.806 ;
			RECT	95.063 40.742 95.095 40.806 ;
			RECT	95.399 40.742 95.431 40.806 ;
			RECT	95.735 40.742 95.767 40.806 ;
			RECT	96.071 40.742 96.103 40.806 ;
			RECT	96.407 40.742 96.439 40.806 ;
			RECT	96.743 40.742 96.775 40.806 ;
			RECT	97.079 40.742 97.111 40.806 ;
			RECT	97.415 40.742 97.447 40.806 ;
			RECT	97.751 40.742 97.783 40.806 ;
			RECT	98.087 40.742 98.119 40.806 ;
			RECT	98.423 40.742 98.455 40.806 ;
			RECT	98.759 40.742 98.791 40.806 ;
			RECT	99.095 40.742 99.127 40.806 ;
			RECT	99.431 40.742 99.463 40.806 ;
			RECT	99.767 40.742 99.799 40.806 ;
			RECT	100.103 40.742 100.135 40.806 ;
			RECT	100.439 40.742 100.471 40.806 ;
			RECT	100.775 40.742 100.807 40.806 ;
			RECT	101.111 40.742 101.143 40.806 ;
			RECT	101.447 40.742 101.479 40.806 ;
			RECT	101.783 40.742 101.815 40.806 ;
			RECT	102.414 40.742 102.446 40.806 ;
			RECT	102.605 40.742 102.637 40.806 ;
			RECT	102.995 40.742 103.027 40.806 ;
			RECT	103.175 40.742 103.207 40.806 ;
			RECT	103.565 40.742 103.597 40.806 ;
			RECT	103.756 40.742 103.788 40.806 ;
			RECT	104.387 40.742 104.419 40.806 ;
			RECT	104.723 40.742 104.755 40.806 ;
			RECT	105.059 40.742 105.091 40.806 ;
			RECT	105.395 40.742 105.427 40.806 ;
			RECT	105.731 40.742 105.763 40.806 ;
			RECT	106.067 40.742 106.099 40.806 ;
			RECT	106.403 40.742 106.435 40.806 ;
			RECT	106.739 40.742 106.771 40.806 ;
			RECT	107.075 40.742 107.107 40.806 ;
			RECT	107.411 40.742 107.443 40.806 ;
			RECT	107.747 40.742 107.779 40.806 ;
			RECT	108.083 40.742 108.115 40.806 ;
			RECT	108.419 40.742 108.451 40.806 ;
			RECT	108.755 40.742 108.787 40.806 ;
			RECT	109.091 40.742 109.123 40.806 ;
			RECT	109.427 40.742 109.459 40.806 ;
			RECT	109.763 40.742 109.795 40.806 ;
			RECT	110.099 40.742 110.131 40.806 ;
			RECT	110.435 40.742 110.467 40.806 ;
			RECT	110.771 40.742 110.803 40.806 ;
			RECT	111.107 40.742 111.139 40.806 ;
			RECT	111.443 40.742 111.475 40.806 ;
			RECT	111.779 40.742 111.811 40.806 ;
			RECT	112.115 40.742 112.147 40.806 ;
			RECT	112.451 40.742 112.483 40.806 ;
			RECT	112.787 40.742 112.819 40.806 ;
			RECT	113.123 40.742 113.155 40.806 ;
			RECT	113.459 40.742 113.491 40.806 ;
			RECT	113.795 40.742 113.827 40.806 ;
			RECT	114.131 40.742 114.163 40.806 ;
			RECT	114.467 40.742 114.499 40.806 ;
			RECT	114.803 40.742 114.835 40.806 ;
			RECT	115.139 40.742 115.171 40.806 ;
			RECT	115.475 40.742 115.507 40.806 ;
			RECT	115.811 40.742 115.843 40.806 ;
			RECT	116.147 40.742 116.179 40.806 ;
			RECT	116.483 40.742 116.515 40.806 ;
			RECT	116.819 40.742 116.851 40.806 ;
			RECT	117.155 40.742 117.187 40.806 ;
			RECT	117.491 40.742 117.523 40.806 ;
			RECT	117.827 40.742 117.859 40.806 ;
			RECT	118.163 40.742 118.195 40.806 ;
			RECT	118.499 40.742 118.531 40.806 ;
			RECT	118.835 40.742 118.867 40.806 ;
			RECT	119.171 40.742 119.203 40.806 ;
			RECT	119.507 40.742 119.539 40.806 ;
			RECT	119.843 40.742 119.875 40.806 ;
			RECT	120.179 40.742 120.211 40.806 ;
			RECT	120.515 40.742 120.547 40.806 ;
			RECT	120.851 40.742 120.883 40.806 ;
			RECT	121.187 40.742 121.219 40.806 ;
			RECT	121.523 40.742 121.555 40.806 ;
			RECT	121.859 40.742 121.891 40.806 ;
			RECT	122.195 40.742 122.227 40.806 ;
			RECT	122.531 40.742 122.563 40.806 ;
			RECT	122.867 40.742 122.899 40.806 ;
			RECT	123.203 40.742 123.235 40.806 ;
			RECT	123.539 40.742 123.571 40.806 ;
			RECT	123.875 40.742 123.907 40.806 ;
			RECT	124.211 40.742 124.243 40.806 ;
			RECT	124.547 40.742 124.579 40.806 ;
			RECT	124.883 40.742 124.915 40.806 ;
			RECT	125.219 40.742 125.251 40.806 ;
			RECT	125.555 40.742 125.587 40.806 ;
			RECT	126.222 40.742 126.254 40.806 ;
			RECT	126.558 40.742 126.59 40.806 ;
			RECT	126.894 40.742 126.926 40.806 ;
			RECT	127.23 40.742 127.262 40.806 ;
			RECT	127.566 40.742 127.598 40.806 ;
			RECT	127.902 40.742 127.934 40.806 ;
			RECT	128.238 40.742 128.27 40.806 ;
			RECT	128.574 40.742 128.606 40.806 ;
			RECT	128.91 40.742 128.942 40.806 ;
			RECT	129.246 40.742 129.278 40.806 ;
			RECT	129.582 40.742 129.614 40.806 ;
			RECT	129.918 40.742 129.95 40.806 ;
			RECT	130.254 40.742 130.286 40.806 ;
			RECT	130.59 40.742 130.622 40.806 ;
			RECT	130.926 40.742 130.958 40.806 ;
			RECT	131.262 40.742 131.294 40.806 ;
			RECT	131.598 40.742 131.63 40.806 ;
			RECT	131.934 40.742 131.966 40.806 ;
			RECT	132.27 40.742 132.302 40.806 ;
			RECT	132.606 40.742 132.638 40.806 ;
			RECT	132.942 40.742 132.974 40.806 ;
			RECT	133.278 40.742 133.31 40.806 ;
			RECT	133.614 40.742 133.646 40.806 ;
			RECT	133.95 40.742 133.982 40.806 ;
			RECT	134.286 40.742 134.318 40.806 ;
			RECT	134.622 40.742 134.654 40.806 ;
			RECT	134.958 40.742 134.99 40.806 ;
			RECT	135.294 40.742 135.326 40.806 ;
			RECT	135.63 40.742 135.662 40.806 ;
			RECT	135.966 40.742 135.998 40.806 ;
			RECT	136.638 40.742 136.67 40.806 ;
			RECT	136.974 40.742 137.006 40.806 ;
			RECT	137.646 40.742 137.678 40.806 ;
			RECT	137.982 40.742 138.014 40.806 ;
			RECT	138.318 40.742 138.35 40.806 ;
			RECT	138.654 40.742 138.686 40.806 ;
			RECT	138.99 40.742 139.022 40.806 ;
			RECT	139.326 40.742 139.358 40.806 ;
			RECT	139.662 40.742 139.694 40.806 ;
			RECT	139.998 40.742 140.03 40.806 ;
			RECT	140.334 40.742 140.366 40.806 ;
			RECT	140.67 40.742 140.702 40.806 ;
			RECT	141.006 40.742 141.038 40.806 ;
			RECT	141.342 40.742 141.374 40.806 ;
			RECT	141.678 40.742 141.71 40.806 ;
			RECT	142.014 40.742 142.046 40.806 ;
			RECT	142.35 40.742 142.382 40.806 ;
			RECT	142.686 40.742 142.718 40.806 ;
			RECT	143.022 40.742 143.054 40.806 ;
			RECT	143.694 40.742 143.726 40.806 ;
			RECT	144.03 40.742 144.062 40.806 ;
			RECT	144.366 40.742 144.398 40.806 ;
			RECT	144.702 40.742 144.734 40.806 ;
			RECT	145.038 40.742 145.07 40.806 ;
			RECT	145.374 40.742 145.406 40.806 ;
			RECT	145.71 40.742 145.742 40.806 ;
			RECT	146.382 40.742 146.414 40.806 ;
			RECT	147.089 40.742 147.121 40.806 ;
			RECT	147.325 40.742 147.357 40.806 ;
			RECT	147.709 40.742 147.741 40.806 ;
			RECT	148.328 40.742 148.36 40.806 ;
			RECT	148.646 40.742 148.678 40.806 ;
			RECT	149.918 40.742 149.95 40.806 ;
			RECT	150.966 40.758 151.03 40.79 ;
			RECT	151.908 40.742 151.94 40.806 ;
			RECT	152.361 40.758 152.425 40.79 ;
			RECT	152.802 40.742 152.834 40.806 ;
			RECT	153.56 40.758 153.624 40.79 ;
			RECT	153.967 40.758 154.031 40.79 ;
			RECT	155.361 40.742 155.393 40.806 ;
			RECT	156.459 40.742 156.491 40.806 ;
			RECT	156.843 40.742 156.875 40.806 ;
			RECT	157.079 40.742 157.111 40.806 ;
			RECT	157.786 40.742 157.818 40.806 ;
			RECT	158.458 40.742 158.49 40.806 ;
			RECT	158.794 40.742 158.826 40.806 ;
			RECT	159.13 40.742 159.162 40.806 ;
			RECT	159.466 40.742 159.498 40.806 ;
			RECT	159.802 40.742 159.834 40.806 ;
			RECT	160.138 40.742 160.17 40.806 ;
			RECT	160.474 40.742 160.506 40.806 ;
			RECT	161.146 40.742 161.178 40.806 ;
			RECT	161.482 40.742 161.514 40.806 ;
			RECT	161.818 40.742 161.85 40.806 ;
			RECT	162.154 40.742 162.186 40.806 ;
			RECT	162.49 40.742 162.522 40.806 ;
			RECT	162.826 40.742 162.858 40.806 ;
			RECT	163.162 40.742 163.194 40.806 ;
			RECT	163.498 40.742 163.53 40.806 ;
			RECT	163.834 40.742 163.866 40.806 ;
			RECT	164.17 40.742 164.202 40.806 ;
			RECT	164.506 40.742 164.538 40.806 ;
			RECT	164.842 40.742 164.874 40.806 ;
			RECT	165.178 40.742 165.21 40.806 ;
			RECT	165.514 40.742 165.546 40.806 ;
			RECT	165.85 40.742 165.882 40.806 ;
			RECT	166.186 40.742 166.218 40.806 ;
			RECT	166.522 40.742 166.554 40.806 ;
			RECT	167.194 40.742 167.226 40.806 ;
			RECT	167.53 40.742 167.562 40.806 ;
			RECT	168.202 40.742 168.234 40.806 ;
			RECT	168.538 40.742 168.57 40.806 ;
			RECT	168.874 40.742 168.906 40.806 ;
			RECT	169.21 40.742 169.242 40.806 ;
			RECT	169.546 40.742 169.578 40.806 ;
			RECT	169.882 40.742 169.914 40.806 ;
			RECT	170.218 40.742 170.25 40.806 ;
			RECT	170.554 40.742 170.586 40.806 ;
			RECT	170.89 40.742 170.922 40.806 ;
			RECT	171.226 40.742 171.258 40.806 ;
			RECT	171.562 40.742 171.594 40.806 ;
			RECT	171.898 40.742 171.93 40.806 ;
			RECT	172.234 40.742 172.266 40.806 ;
			RECT	172.57 40.742 172.602 40.806 ;
			RECT	172.906 40.742 172.938 40.806 ;
			RECT	173.242 40.742 173.274 40.806 ;
			RECT	173.578 40.742 173.61 40.806 ;
			RECT	173.914 40.742 173.946 40.806 ;
			RECT	174.25 40.742 174.282 40.806 ;
			RECT	174.586 40.742 174.618 40.806 ;
			RECT	174.922 40.742 174.954 40.806 ;
			RECT	175.258 40.742 175.29 40.806 ;
			RECT	175.594 40.742 175.626 40.806 ;
			RECT	175.93 40.742 175.962 40.806 ;
			RECT	176.266 40.742 176.298 40.806 ;
			RECT	176.602 40.742 176.634 40.806 ;
			RECT	176.938 40.742 176.97 40.806 ;
			RECT	177.274 40.742 177.306 40.806 ;
			RECT	177.61 40.742 177.642 40.806 ;
			RECT	177.946 40.742 177.978 40.806 ;
			RECT	178.613 40.742 178.645 40.806 ;
			RECT	178.949 40.742 178.981 40.806 ;
			RECT	179.285 40.742 179.317 40.806 ;
			RECT	179.621 40.742 179.653 40.806 ;
			RECT	179.957 40.742 179.989 40.806 ;
			RECT	180.293 40.742 180.325 40.806 ;
			RECT	180.629 40.742 180.661 40.806 ;
			RECT	180.965 40.742 180.997 40.806 ;
			RECT	181.301 40.742 181.333 40.806 ;
			RECT	181.637 40.742 181.669 40.806 ;
			RECT	181.973 40.742 182.005 40.806 ;
			RECT	182.309 40.742 182.341 40.806 ;
			RECT	182.645 40.742 182.677 40.806 ;
			RECT	182.981 40.742 183.013 40.806 ;
			RECT	183.317 40.742 183.349 40.806 ;
			RECT	183.653 40.742 183.685 40.806 ;
			RECT	183.989 40.742 184.021 40.806 ;
			RECT	184.325 40.742 184.357 40.806 ;
			RECT	184.661 40.742 184.693 40.806 ;
			RECT	184.997 40.742 185.029 40.806 ;
			RECT	185.333 40.742 185.365 40.806 ;
			RECT	185.669 40.742 185.701 40.806 ;
			RECT	186.005 40.742 186.037 40.806 ;
			RECT	186.341 40.742 186.373 40.806 ;
			RECT	186.677 40.742 186.709 40.806 ;
			RECT	187.013 40.742 187.045 40.806 ;
			RECT	187.349 40.742 187.381 40.806 ;
			RECT	187.685 40.742 187.717 40.806 ;
			RECT	188.021 40.742 188.053 40.806 ;
			RECT	188.357 40.742 188.389 40.806 ;
			RECT	188.693 40.742 188.725 40.806 ;
			RECT	189.029 40.742 189.061 40.806 ;
			RECT	189.365 40.742 189.397 40.806 ;
			RECT	189.701 40.742 189.733 40.806 ;
			RECT	190.037 40.742 190.069 40.806 ;
			RECT	190.373 40.742 190.405 40.806 ;
			RECT	190.709 40.742 190.741 40.806 ;
			RECT	191.045 40.742 191.077 40.806 ;
			RECT	191.381 40.742 191.413 40.806 ;
			RECT	191.717 40.742 191.749 40.806 ;
			RECT	192.053 40.742 192.085 40.806 ;
			RECT	192.389 40.742 192.421 40.806 ;
			RECT	192.725 40.742 192.757 40.806 ;
			RECT	193.061 40.742 193.093 40.806 ;
			RECT	193.397 40.742 193.429 40.806 ;
			RECT	193.733 40.742 193.765 40.806 ;
			RECT	194.069 40.742 194.101 40.806 ;
			RECT	194.405 40.742 194.437 40.806 ;
			RECT	194.741 40.742 194.773 40.806 ;
			RECT	195.077 40.742 195.109 40.806 ;
			RECT	195.413 40.742 195.445 40.806 ;
			RECT	195.749 40.742 195.781 40.806 ;
			RECT	196.085 40.742 196.117 40.806 ;
			RECT	196.421 40.742 196.453 40.806 ;
			RECT	196.757 40.742 196.789 40.806 ;
			RECT	197.093 40.742 197.125 40.806 ;
			RECT	197.429 40.742 197.461 40.806 ;
			RECT	197.765 40.742 197.797 40.806 ;
			RECT	198.101 40.742 198.133 40.806 ;
			RECT	198.437 40.742 198.469 40.806 ;
			RECT	198.773 40.742 198.805 40.806 ;
			RECT	199.109 40.742 199.141 40.806 ;
			RECT	199.445 40.742 199.477 40.806 ;
			RECT	199.781 40.742 199.813 40.806 ;
			RECT	200.412 40.742 200.444 40.806 ;
			RECT	200.603 40.742 200.635 40.806 ;
			RECT	201.403 40.742 201.435 40.806 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 43.598 201.665 43.718 ;
			LAYER	J3 ;
			RECT	0.703 43.642 0.735 43.674 ;
			RECT	1.164 43.626 1.196 43.69 ;
			RECT	1.645 43.626 1.709 43.69 ;
			RECT	2.197 43.626 2.229 43.69 ;
			RECT	2.343 43.626 2.375 43.69 ;
			RECT	3.451 43.626 3.483 43.69 ;
			RECT	4.354 43.626 4.386 43.69 ;
			RECT	4.61 43.626 4.642 43.69 ;
			RECT	4.805 43.626 4.837 43.69 ;
			RECT	5.567 43.626 5.599 43.69 ;
			RECT	6.389 43.626 6.421 43.69 ;
			RECT	6.725 43.626 6.757 43.69 ;
			RECT	7.061 43.626 7.093 43.69 ;
			RECT	7.397 43.626 7.429 43.69 ;
			RECT	7.733 43.626 7.765 43.69 ;
			RECT	8.069 43.626 8.101 43.69 ;
			RECT	8.405 43.626 8.437 43.69 ;
			RECT	8.741 43.626 8.773 43.69 ;
			RECT	9.077 43.626 9.109 43.69 ;
			RECT	9.413 43.626 9.445 43.69 ;
			RECT	9.749 43.626 9.781 43.69 ;
			RECT	10.085 43.626 10.117 43.69 ;
			RECT	10.421 43.626 10.453 43.69 ;
			RECT	10.757 43.626 10.789 43.69 ;
			RECT	11.093 43.626 11.125 43.69 ;
			RECT	11.429 43.626 11.461 43.69 ;
			RECT	11.765 43.626 11.797 43.69 ;
			RECT	12.101 43.626 12.133 43.69 ;
			RECT	12.437 43.626 12.469 43.69 ;
			RECT	12.773 43.626 12.805 43.69 ;
			RECT	13.109 43.626 13.141 43.69 ;
			RECT	13.445 43.626 13.477 43.69 ;
			RECT	13.781 43.626 13.813 43.69 ;
			RECT	14.117 43.626 14.149 43.69 ;
			RECT	14.453 43.626 14.485 43.69 ;
			RECT	14.789 43.626 14.821 43.69 ;
			RECT	15.125 43.626 15.157 43.69 ;
			RECT	15.461 43.626 15.493 43.69 ;
			RECT	15.797 43.626 15.829 43.69 ;
			RECT	16.133 43.626 16.165 43.69 ;
			RECT	16.469 43.626 16.501 43.69 ;
			RECT	16.805 43.626 16.837 43.69 ;
			RECT	17.141 43.626 17.173 43.69 ;
			RECT	17.477 43.626 17.509 43.69 ;
			RECT	17.813 43.626 17.845 43.69 ;
			RECT	18.149 43.626 18.181 43.69 ;
			RECT	18.485 43.626 18.517 43.69 ;
			RECT	18.821 43.626 18.853 43.69 ;
			RECT	19.157 43.626 19.189 43.69 ;
			RECT	19.493 43.626 19.525 43.69 ;
			RECT	19.829 43.626 19.861 43.69 ;
			RECT	20.165 43.626 20.197 43.69 ;
			RECT	20.501 43.626 20.533 43.69 ;
			RECT	20.837 43.626 20.869 43.69 ;
			RECT	21.173 43.626 21.205 43.69 ;
			RECT	21.509 43.626 21.541 43.69 ;
			RECT	21.845 43.626 21.877 43.69 ;
			RECT	22.181 43.626 22.213 43.69 ;
			RECT	22.517 43.626 22.549 43.69 ;
			RECT	22.853 43.626 22.885 43.69 ;
			RECT	23.189 43.626 23.221 43.69 ;
			RECT	23.525 43.626 23.557 43.69 ;
			RECT	23.861 43.626 23.893 43.69 ;
			RECT	24.197 43.626 24.229 43.69 ;
			RECT	24.533 43.626 24.565 43.69 ;
			RECT	24.869 43.626 24.901 43.69 ;
			RECT	25.205 43.626 25.237 43.69 ;
			RECT	25.541 43.626 25.573 43.69 ;
			RECT	25.877 43.626 25.909 43.69 ;
			RECT	26.213 43.626 26.245 43.69 ;
			RECT	26.549 43.626 26.581 43.69 ;
			RECT	26.885 43.626 26.917 43.69 ;
			RECT	27.221 43.626 27.253 43.69 ;
			RECT	27.557 43.626 27.589 43.69 ;
			RECT	27.888 43.626 27.92 43.69 ;
			RECT	28.56 43.626 28.592 43.69 ;
			RECT	29.232 43.626 29.264 43.69 ;
			RECT	29.568 43.626 29.6 43.69 ;
			RECT	29.904 43.626 29.936 43.69 ;
			RECT	30.24 43.626 30.272 43.69 ;
			RECT	30.576 43.626 30.608 43.69 ;
			RECT	30.912 43.626 30.944 43.69 ;
			RECT	31.584 43.626 31.616 43.69 ;
			RECT	31.92 43.626 31.952 43.69 ;
			RECT	32.592 43.626 32.624 43.69 ;
			RECT	33.264 43.626 33.296 43.69 ;
			RECT	34.272 43.626 34.304 43.69 ;
			RECT	34.608 43.626 34.64 43.69 ;
			RECT	35.616 43.626 35.648 43.69 ;
			RECT	35.952 43.626 35.984 43.69 ;
			RECT	36.96 43.626 36.992 43.69 ;
			RECT	37.296 43.626 37.328 43.69 ;
			RECT	38.304 43.626 38.336 43.69 ;
			RECT	38.64 43.626 38.672 43.69 ;
			RECT	39.648 43.626 39.68 43.69 ;
			RECT	40.32 43.626 40.352 43.69 ;
			RECT	41.328 43.626 41.36 43.69 ;
			RECT	42.672 43.626 42.704 43.69 ;
			RECT	43.68 43.626 43.712 43.69 ;
			RECT	44.016 43.626 44.048 43.69 ;
			RECT	44.201 43.626 44.233 43.69 ;
			RECT	45.36 43.626 45.392 43.69 ;
			RECT	46.032 43.626 46.064 43.69 ;
			RECT	47.04 43.626 47.072 43.69 ;
			RECT	48.52 43.626 48.584 43.69 ;
			RECT	49.056 43.626 49.088 43.69 ;
			RECT	49.327 43.626 49.359 43.69 ;
			RECT	49.675 43.626 49.707 43.69 ;
			RECT	50.33 43.626 50.362 43.69 ;
			RECT	52.026 43.626 52.058 43.69 ;
			RECT	52.968 43.626 53.032 43.69 ;
			RECT	53.91 43.626 53.942 43.69 ;
			RECT	54.251 43.642 54.283 43.674 ;
			RECT	55.562 43.626 55.626 43.69 ;
			RECT	55.842 43.626 55.874 43.69 ;
			RECT	55.969 43.626 56.033 43.69 ;
			RECT	58.497 43.626 58.529 43.69 ;
			RECT	58.845 43.626 58.877 43.69 ;
			RECT	59.116 43.626 59.148 43.69 ;
			RECT	59.62 43.626 59.684 43.69 ;
			RECT	61.132 43.626 61.164 43.69 ;
			RECT	62.14 43.626 62.172 43.69 ;
			RECT	62.812 43.626 62.844 43.69 ;
			RECT	63.971 43.626 64.003 43.69 ;
			RECT	64.156 43.626 64.188 43.69 ;
			RECT	64.492 43.626 64.524 43.69 ;
			RECT	65.5 43.626 65.532 43.69 ;
			RECT	66.844 43.626 66.876 43.69 ;
			RECT	67.852 43.626 67.884 43.69 ;
			RECT	68.524 43.626 68.556 43.69 ;
			RECT	69.532 43.626 69.564 43.69 ;
			RECT	69.868 43.626 69.9 43.69 ;
			RECT	70.876 43.626 70.908 43.69 ;
			RECT	71.212 43.626 71.244 43.69 ;
			RECT	72.22 43.626 72.252 43.69 ;
			RECT	72.556 43.626 72.588 43.69 ;
			RECT	73.564 43.626 73.596 43.69 ;
			RECT	73.9 43.626 73.932 43.69 ;
			RECT	74.908 43.626 74.94 43.69 ;
			RECT	75.58 43.626 75.612 43.69 ;
			RECT	76.252 43.626 76.284 43.69 ;
			RECT	76.588 43.626 76.62 43.69 ;
			RECT	77.26 43.626 77.292 43.69 ;
			RECT	77.596 43.626 77.628 43.69 ;
			RECT	77.932 43.626 77.964 43.69 ;
			RECT	78.268 43.626 78.3 43.69 ;
			RECT	78.604 43.626 78.636 43.69 ;
			RECT	78.94 43.626 78.972 43.69 ;
			RECT	79.612 43.626 79.644 43.69 ;
			RECT	80.284 43.626 80.316 43.69 ;
			RECT	80.615 43.626 80.647 43.69 ;
			RECT	80.951 43.626 80.983 43.69 ;
			RECT	81.287 43.626 81.319 43.69 ;
			RECT	81.623 43.626 81.655 43.69 ;
			RECT	81.959 43.626 81.991 43.69 ;
			RECT	82.295 43.626 82.327 43.69 ;
			RECT	82.631 43.626 82.663 43.69 ;
			RECT	82.967 43.626 82.999 43.69 ;
			RECT	83.303 43.626 83.335 43.69 ;
			RECT	83.639 43.626 83.671 43.69 ;
			RECT	83.975 43.626 84.007 43.69 ;
			RECT	84.311 43.626 84.343 43.69 ;
			RECT	84.647 43.626 84.679 43.69 ;
			RECT	84.983 43.626 85.015 43.69 ;
			RECT	85.319 43.626 85.351 43.69 ;
			RECT	85.655 43.626 85.687 43.69 ;
			RECT	85.991 43.626 86.023 43.69 ;
			RECT	86.327 43.626 86.359 43.69 ;
			RECT	86.663 43.626 86.695 43.69 ;
			RECT	86.999 43.626 87.031 43.69 ;
			RECT	87.335 43.626 87.367 43.69 ;
			RECT	87.671 43.626 87.703 43.69 ;
			RECT	88.007 43.626 88.039 43.69 ;
			RECT	88.343 43.626 88.375 43.69 ;
			RECT	88.679 43.626 88.711 43.69 ;
			RECT	89.015 43.626 89.047 43.69 ;
			RECT	89.351 43.626 89.383 43.69 ;
			RECT	89.687 43.626 89.719 43.69 ;
			RECT	90.023 43.626 90.055 43.69 ;
			RECT	90.359 43.626 90.391 43.69 ;
			RECT	90.695 43.626 90.727 43.69 ;
			RECT	91.031 43.626 91.063 43.69 ;
			RECT	91.367 43.626 91.399 43.69 ;
			RECT	91.703 43.626 91.735 43.69 ;
			RECT	92.039 43.626 92.071 43.69 ;
			RECT	92.375 43.626 92.407 43.69 ;
			RECT	92.711 43.626 92.743 43.69 ;
			RECT	93.047 43.626 93.079 43.69 ;
			RECT	93.383 43.626 93.415 43.69 ;
			RECT	93.719 43.626 93.751 43.69 ;
			RECT	94.055 43.626 94.087 43.69 ;
			RECT	94.391 43.626 94.423 43.69 ;
			RECT	94.727 43.626 94.759 43.69 ;
			RECT	95.063 43.626 95.095 43.69 ;
			RECT	95.399 43.626 95.431 43.69 ;
			RECT	95.735 43.626 95.767 43.69 ;
			RECT	96.071 43.626 96.103 43.69 ;
			RECT	96.407 43.626 96.439 43.69 ;
			RECT	96.743 43.626 96.775 43.69 ;
			RECT	97.079 43.626 97.111 43.69 ;
			RECT	97.415 43.626 97.447 43.69 ;
			RECT	97.751 43.626 97.783 43.69 ;
			RECT	98.087 43.626 98.119 43.69 ;
			RECT	98.423 43.626 98.455 43.69 ;
			RECT	98.759 43.626 98.791 43.69 ;
			RECT	99.095 43.626 99.127 43.69 ;
			RECT	99.431 43.626 99.463 43.69 ;
			RECT	99.767 43.626 99.799 43.69 ;
			RECT	100.103 43.626 100.135 43.69 ;
			RECT	100.439 43.626 100.471 43.69 ;
			RECT	100.775 43.626 100.807 43.69 ;
			RECT	101.111 43.626 101.143 43.69 ;
			RECT	101.447 43.626 101.479 43.69 ;
			RECT	101.783 43.626 101.815 43.69 ;
			RECT	102.605 43.626 102.637 43.69 ;
			RECT	102.994 43.626 103.026 43.69 ;
			RECT	103.176 43.626 103.208 43.69 ;
			RECT	103.565 43.626 103.597 43.69 ;
			RECT	104.387 43.626 104.419 43.69 ;
			RECT	104.723 43.626 104.755 43.69 ;
			RECT	105.059 43.626 105.091 43.69 ;
			RECT	105.395 43.626 105.427 43.69 ;
			RECT	105.731 43.626 105.763 43.69 ;
			RECT	106.067 43.626 106.099 43.69 ;
			RECT	106.403 43.626 106.435 43.69 ;
			RECT	106.739 43.626 106.771 43.69 ;
			RECT	107.075 43.626 107.107 43.69 ;
			RECT	107.411 43.626 107.443 43.69 ;
			RECT	107.747 43.626 107.779 43.69 ;
			RECT	108.083 43.626 108.115 43.69 ;
			RECT	108.419 43.626 108.451 43.69 ;
			RECT	108.755 43.626 108.787 43.69 ;
			RECT	109.091 43.626 109.123 43.69 ;
			RECT	109.427 43.626 109.459 43.69 ;
			RECT	109.763 43.626 109.795 43.69 ;
			RECT	110.099 43.626 110.131 43.69 ;
			RECT	110.435 43.626 110.467 43.69 ;
			RECT	110.771 43.626 110.803 43.69 ;
			RECT	111.107 43.626 111.139 43.69 ;
			RECT	111.443 43.626 111.475 43.69 ;
			RECT	111.779 43.626 111.811 43.69 ;
			RECT	112.115 43.626 112.147 43.69 ;
			RECT	112.451 43.626 112.483 43.69 ;
			RECT	112.787 43.626 112.819 43.69 ;
			RECT	113.123 43.626 113.155 43.69 ;
			RECT	113.459 43.626 113.491 43.69 ;
			RECT	113.795 43.626 113.827 43.69 ;
			RECT	114.131 43.626 114.163 43.69 ;
			RECT	114.467 43.626 114.499 43.69 ;
			RECT	114.803 43.626 114.835 43.69 ;
			RECT	115.139 43.626 115.171 43.69 ;
			RECT	115.475 43.626 115.507 43.69 ;
			RECT	115.811 43.626 115.843 43.69 ;
			RECT	116.147 43.626 116.179 43.69 ;
			RECT	116.483 43.626 116.515 43.69 ;
			RECT	116.819 43.626 116.851 43.69 ;
			RECT	117.155 43.626 117.187 43.69 ;
			RECT	117.491 43.626 117.523 43.69 ;
			RECT	117.827 43.626 117.859 43.69 ;
			RECT	118.163 43.626 118.195 43.69 ;
			RECT	118.499 43.626 118.531 43.69 ;
			RECT	118.835 43.626 118.867 43.69 ;
			RECT	119.171 43.626 119.203 43.69 ;
			RECT	119.507 43.626 119.539 43.69 ;
			RECT	119.843 43.626 119.875 43.69 ;
			RECT	120.179 43.626 120.211 43.69 ;
			RECT	120.515 43.626 120.547 43.69 ;
			RECT	120.851 43.626 120.883 43.69 ;
			RECT	121.187 43.626 121.219 43.69 ;
			RECT	121.523 43.626 121.555 43.69 ;
			RECT	121.859 43.626 121.891 43.69 ;
			RECT	122.195 43.626 122.227 43.69 ;
			RECT	122.531 43.626 122.563 43.69 ;
			RECT	122.867 43.626 122.899 43.69 ;
			RECT	123.203 43.626 123.235 43.69 ;
			RECT	123.539 43.626 123.571 43.69 ;
			RECT	123.875 43.626 123.907 43.69 ;
			RECT	124.211 43.626 124.243 43.69 ;
			RECT	124.547 43.626 124.579 43.69 ;
			RECT	124.883 43.626 124.915 43.69 ;
			RECT	125.219 43.626 125.251 43.69 ;
			RECT	125.555 43.626 125.587 43.69 ;
			RECT	125.886 43.626 125.918 43.69 ;
			RECT	126.558 43.626 126.59 43.69 ;
			RECT	127.23 43.626 127.262 43.69 ;
			RECT	127.566 43.626 127.598 43.69 ;
			RECT	127.902 43.626 127.934 43.69 ;
			RECT	128.238 43.626 128.27 43.69 ;
			RECT	128.574 43.626 128.606 43.69 ;
			RECT	128.91 43.626 128.942 43.69 ;
			RECT	129.582 43.626 129.614 43.69 ;
			RECT	129.918 43.626 129.95 43.69 ;
			RECT	130.59 43.626 130.622 43.69 ;
			RECT	131.262 43.626 131.294 43.69 ;
			RECT	132.27 43.626 132.302 43.69 ;
			RECT	132.606 43.626 132.638 43.69 ;
			RECT	133.614 43.626 133.646 43.69 ;
			RECT	133.95 43.626 133.982 43.69 ;
			RECT	134.958 43.626 134.99 43.69 ;
			RECT	135.294 43.626 135.326 43.69 ;
			RECT	136.302 43.626 136.334 43.69 ;
			RECT	136.638 43.626 136.67 43.69 ;
			RECT	137.646 43.626 137.678 43.69 ;
			RECT	138.318 43.626 138.35 43.69 ;
			RECT	139.326 43.626 139.358 43.69 ;
			RECT	140.67 43.626 140.702 43.69 ;
			RECT	141.678 43.626 141.71 43.69 ;
			RECT	142.014 43.626 142.046 43.69 ;
			RECT	142.199 43.626 142.231 43.69 ;
			RECT	143.358 43.626 143.39 43.69 ;
			RECT	144.03 43.626 144.062 43.69 ;
			RECT	145.038 43.626 145.07 43.69 ;
			RECT	146.518 43.626 146.582 43.69 ;
			RECT	147.054 43.626 147.086 43.69 ;
			RECT	147.325 43.626 147.357 43.69 ;
			RECT	147.673 43.626 147.705 43.69 ;
			RECT	148.328 43.626 148.36 43.69 ;
			RECT	150.024 43.626 150.056 43.69 ;
			RECT	150.966 43.626 151.03 43.69 ;
			RECT	151.908 43.626 151.94 43.69 ;
			RECT	152.249 43.642 152.281 43.674 ;
			RECT	153.56 43.626 153.624 43.69 ;
			RECT	153.84 43.626 153.872 43.69 ;
			RECT	153.967 43.626 154.031 43.69 ;
			RECT	156.495 43.626 156.527 43.69 ;
			RECT	156.843 43.626 156.875 43.69 ;
			RECT	157.114 43.626 157.146 43.69 ;
			RECT	157.618 43.626 157.682 43.69 ;
			RECT	159.13 43.626 159.162 43.69 ;
			RECT	160.138 43.626 160.17 43.69 ;
			RECT	160.81 43.626 160.842 43.69 ;
			RECT	161.969 43.626 162.001 43.69 ;
			RECT	162.154 43.626 162.186 43.69 ;
			RECT	162.49 43.626 162.522 43.69 ;
			RECT	163.498 43.626 163.53 43.69 ;
			RECT	164.842 43.626 164.874 43.69 ;
			RECT	165.85 43.626 165.882 43.69 ;
			RECT	166.522 43.626 166.554 43.69 ;
			RECT	167.53 43.626 167.562 43.69 ;
			RECT	167.866 43.626 167.898 43.69 ;
			RECT	168.874 43.626 168.906 43.69 ;
			RECT	169.21 43.626 169.242 43.69 ;
			RECT	170.218 43.626 170.25 43.69 ;
			RECT	170.554 43.626 170.586 43.69 ;
			RECT	171.562 43.626 171.594 43.69 ;
			RECT	171.898 43.626 171.93 43.69 ;
			RECT	172.906 43.626 172.938 43.69 ;
			RECT	173.578 43.626 173.61 43.69 ;
			RECT	174.25 43.626 174.282 43.69 ;
			RECT	174.586 43.626 174.618 43.69 ;
			RECT	175.258 43.626 175.29 43.69 ;
			RECT	175.594 43.626 175.626 43.69 ;
			RECT	175.93 43.626 175.962 43.69 ;
			RECT	176.266 43.626 176.298 43.69 ;
			RECT	176.602 43.626 176.634 43.69 ;
			RECT	176.938 43.626 176.97 43.69 ;
			RECT	177.61 43.626 177.642 43.69 ;
			RECT	178.282 43.626 178.314 43.69 ;
			RECT	178.613 43.626 178.645 43.69 ;
			RECT	178.949 43.626 178.981 43.69 ;
			RECT	179.285 43.626 179.317 43.69 ;
			RECT	179.621 43.626 179.653 43.69 ;
			RECT	179.957 43.626 179.989 43.69 ;
			RECT	180.293 43.626 180.325 43.69 ;
			RECT	180.629 43.626 180.661 43.69 ;
			RECT	180.965 43.626 180.997 43.69 ;
			RECT	181.301 43.626 181.333 43.69 ;
			RECT	181.637 43.626 181.669 43.69 ;
			RECT	181.973 43.626 182.005 43.69 ;
			RECT	182.309 43.626 182.341 43.69 ;
			RECT	182.645 43.626 182.677 43.69 ;
			RECT	182.981 43.626 183.013 43.69 ;
			RECT	183.317 43.626 183.349 43.69 ;
			RECT	183.653 43.626 183.685 43.69 ;
			RECT	183.989 43.626 184.021 43.69 ;
			RECT	184.325 43.626 184.357 43.69 ;
			RECT	184.661 43.626 184.693 43.69 ;
			RECT	184.997 43.626 185.029 43.69 ;
			RECT	185.333 43.626 185.365 43.69 ;
			RECT	185.669 43.626 185.701 43.69 ;
			RECT	186.005 43.626 186.037 43.69 ;
			RECT	186.341 43.626 186.373 43.69 ;
			RECT	186.677 43.626 186.709 43.69 ;
			RECT	187.013 43.626 187.045 43.69 ;
			RECT	187.349 43.626 187.381 43.69 ;
			RECT	187.685 43.626 187.717 43.69 ;
			RECT	188.021 43.626 188.053 43.69 ;
			RECT	188.357 43.626 188.389 43.69 ;
			RECT	188.693 43.626 188.725 43.69 ;
			RECT	189.029 43.626 189.061 43.69 ;
			RECT	189.365 43.626 189.397 43.69 ;
			RECT	189.701 43.626 189.733 43.69 ;
			RECT	190.037 43.626 190.069 43.69 ;
			RECT	190.373 43.626 190.405 43.69 ;
			RECT	190.709 43.626 190.741 43.69 ;
			RECT	191.045 43.626 191.077 43.69 ;
			RECT	191.381 43.626 191.413 43.69 ;
			RECT	191.717 43.626 191.749 43.69 ;
			RECT	192.053 43.626 192.085 43.69 ;
			RECT	192.389 43.626 192.421 43.69 ;
			RECT	192.725 43.626 192.757 43.69 ;
			RECT	193.061 43.626 193.093 43.69 ;
			RECT	193.397 43.626 193.429 43.69 ;
			RECT	193.733 43.626 193.765 43.69 ;
			RECT	194.069 43.626 194.101 43.69 ;
			RECT	194.405 43.626 194.437 43.69 ;
			RECT	194.741 43.626 194.773 43.69 ;
			RECT	195.077 43.626 195.109 43.69 ;
			RECT	195.413 43.626 195.445 43.69 ;
			RECT	195.749 43.626 195.781 43.69 ;
			RECT	196.085 43.626 196.117 43.69 ;
			RECT	196.421 43.626 196.453 43.69 ;
			RECT	196.757 43.626 196.789 43.69 ;
			RECT	197.093 43.626 197.125 43.69 ;
			RECT	197.429 43.626 197.461 43.69 ;
			RECT	197.765 43.626 197.797 43.69 ;
			RECT	198.101 43.626 198.133 43.69 ;
			RECT	198.437 43.626 198.469 43.69 ;
			RECT	198.773 43.626 198.805 43.69 ;
			RECT	199.109 43.626 199.141 43.69 ;
			RECT	199.445 43.626 199.477 43.69 ;
			RECT	199.781 43.626 199.813 43.69 ;
			RECT	200.603 43.626 200.635 43.69 ;
			RECT	201.403 43.626 201.435 43.69 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 48.828 201.665 48.938 ;
			LAYER	J3 ;
			RECT	0.755 48.851 0.787 48.915 ;
			RECT	1.164 48.851 1.196 48.915 ;
			RECT	1.645 48.851 1.709 48.915 ;
			RECT	2.339 48.851 2.371 48.915 ;
			RECT	4.195 48.851 4.227 48.915 ;
			RECT	4.944 48.851 5.008 48.915 ;
			RECT	5.809 48.851 5.841 48.915 ;
			RECT	6.095 48.851 6.127 48.915 ;
			RECT	6.347 48.851 6.379 48.915 ;
			RECT	6.683 48.851 6.715 48.915 ;
			RECT	7.019 48.851 7.051 48.915 ;
			RECT	7.355 48.851 7.387 48.915 ;
			RECT	7.691 48.851 7.723 48.915 ;
			RECT	8.027 48.851 8.059 48.915 ;
			RECT	8.363 48.851 8.395 48.915 ;
			RECT	8.699 48.851 8.731 48.915 ;
			RECT	9.035 48.851 9.067 48.915 ;
			RECT	9.371 48.851 9.403 48.915 ;
			RECT	9.707 48.851 9.739 48.915 ;
			RECT	10.043 48.851 10.075 48.915 ;
			RECT	10.379 48.851 10.411 48.915 ;
			RECT	10.715 48.851 10.747 48.915 ;
			RECT	11.051 48.851 11.083 48.915 ;
			RECT	11.387 48.851 11.419 48.915 ;
			RECT	11.723 48.851 11.755 48.915 ;
			RECT	12.059 48.851 12.091 48.915 ;
			RECT	12.395 48.851 12.427 48.915 ;
			RECT	12.731 48.851 12.763 48.915 ;
			RECT	13.067 48.851 13.099 48.915 ;
			RECT	13.403 48.851 13.435 48.915 ;
			RECT	13.739 48.851 13.771 48.915 ;
			RECT	14.075 48.851 14.107 48.915 ;
			RECT	14.411 48.851 14.443 48.915 ;
			RECT	14.747 48.851 14.779 48.915 ;
			RECT	15.083 48.851 15.115 48.915 ;
			RECT	15.419 48.851 15.451 48.915 ;
			RECT	15.755 48.851 15.787 48.915 ;
			RECT	16.091 48.851 16.123 48.915 ;
			RECT	16.427 48.851 16.459 48.915 ;
			RECT	16.763 48.851 16.795 48.915 ;
			RECT	17.099 48.851 17.131 48.915 ;
			RECT	17.435 48.851 17.467 48.915 ;
			RECT	17.771 48.851 17.803 48.915 ;
			RECT	18.107 48.851 18.139 48.915 ;
			RECT	18.443 48.851 18.475 48.915 ;
			RECT	18.779 48.851 18.811 48.915 ;
			RECT	19.115 48.851 19.147 48.915 ;
			RECT	19.451 48.851 19.483 48.915 ;
			RECT	19.787 48.851 19.819 48.915 ;
			RECT	20.123 48.851 20.155 48.915 ;
			RECT	20.459 48.851 20.491 48.915 ;
			RECT	20.795 48.851 20.827 48.915 ;
			RECT	21.131 48.851 21.163 48.915 ;
			RECT	21.467 48.851 21.499 48.915 ;
			RECT	21.803 48.851 21.835 48.915 ;
			RECT	22.139 48.851 22.171 48.915 ;
			RECT	22.475 48.851 22.507 48.915 ;
			RECT	22.811 48.851 22.843 48.915 ;
			RECT	23.147 48.851 23.179 48.915 ;
			RECT	23.483 48.851 23.515 48.915 ;
			RECT	23.819 48.851 23.851 48.915 ;
			RECT	24.155 48.851 24.187 48.915 ;
			RECT	24.491 48.851 24.523 48.915 ;
			RECT	24.827 48.851 24.859 48.915 ;
			RECT	25.163 48.851 25.195 48.915 ;
			RECT	25.499 48.851 25.531 48.915 ;
			RECT	25.835 48.851 25.867 48.915 ;
			RECT	26.171 48.851 26.203 48.915 ;
			RECT	26.507 48.851 26.539 48.915 ;
			RECT	26.843 48.851 26.875 48.915 ;
			RECT	27.179 48.851 27.211 48.915 ;
			RECT	27.515 48.851 27.547 48.915 ;
			RECT	27.851 48.851 27.883 48.915 ;
			RECT	28.019 48.851 28.051 48.915 ;
			RECT	28.187 48.851 28.219 48.915 ;
			RECT	28.355 48.851 28.387 48.915 ;
			RECT	28.523 48.851 28.555 48.915 ;
			RECT	28.691 48.851 28.723 48.915 ;
			RECT	28.859 48.851 28.891 48.915 ;
			RECT	29.027 48.851 29.059 48.915 ;
			RECT	29.195 48.851 29.227 48.915 ;
			RECT	29.363 48.851 29.395 48.915 ;
			RECT	29.531 48.851 29.563 48.915 ;
			RECT	29.699 48.851 29.731 48.915 ;
			RECT	29.867 48.851 29.899 48.915 ;
			RECT	30.035 48.851 30.067 48.915 ;
			RECT	30.203 48.851 30.235 48.915 ;
			RECT	30.371 48.851 30.403 48.915 ;
			RECT	30.539 48.851 30.571 48.915 ;
			RECT	30.707 48.851 30.739 48.915 ;
			RECT	30.875 48.851 30.907 48.915 ;
			RECT	31.043 48.851 31.075 48.915 ;
			RECT	31.211 48.851 31.243 48.915 ;
			RECT	31.379 48.851 31.411 48.915 ;
			RECT	31.547 48.851 31.579 48.915 ;
			RECT	31.715 48.851 31.747 48.915 ;
			RECT	31.883 48.851 31.915 48.915 ;
			RECT	32.051 48.851 32.083 48.915 ;
			RECT	32.219 48.851 32.251 48.915 ;
			RECT	32.387 48.851 32.419 48.915 ;
			RECT	32.555 48.851 32.587 48.915 ;
			RECT	32.723 48.851 32.755 48.915 ;
			RECT	32.891 48.851 32.923 48.915 ;
			RECT	33.059 48.851 33.091 48.915 ;
			RECT	33.227 48.851 33.259 48.915 ;
			RECT	33.395 48.851 33.427 48.915 ;
			RECT	33.563 48.851 33.595 48.915 ;
			RECT	33.731 48.851 33.763 48.915 ;
			RECT	33.899 48.851 33.931 48.915 ;
			RECT	34.067 48.851 34.099 48.915 ;
			RECT	34.235 48.851 34.267 48.915 ;
			RECT	34.403 48.851 34.435 48.915 ;
			RECT	34.571 48.851 34.603 48.915 ;
			RECT	34.739 48.851 34.771 48.915 ;
			RECT	34.907 48.851 34.939 48.915 ;
			RECT	35.075 48.851 35.107 48.915 ;
			RECT	35.243 48.851 35.275 48.915 ;
			RECT	35.411 48.851 35.443 48.915 ;
			RECT	35.579 48.851 35.611 48.915 ;
			RECT	35.747 48.851 35.779 48.915 ;
			RECT	35.915 48.851 35.947 48.915 ;
			RECT	36.083 48.851 36.115 48.915 ;
			RECT	36.251 48.851 36.283 48.915 ;
			RECT	36.419 48.851 36.451 48.915 ;
			RECT	36.587 48.851 36.619 48.915 ;
			RECT	36.755 48.851 36.787 48.915 ;
			RECT	36.923 48.851 36.955 48.915 ;
			RECT	37.091 48.851 37.123 48.915 ;
			RECT	37.259 48.851 37.291 48.915 ;
			RECT	37.427 48.851 37.459 48.915 ;
			RECT	37.595 48.851 37.627 48.915 ;
			RECT	37.763 48.851 37.795 48.915 ;
			RECT	37.931 48.851 37.963 48.915 ;
			RECT	38.099 48.851 38.131 48.915 ;
			RECT	38.267 48.851 38.299 48.915 ;
			RECT	38.435 48.851 38.467 48.915 ;
			RECT	38.603 48.851 38.635 48.915 ;
			RECT	38.771 48.851 38.803 48.915 ;
			RECT	38.939 48.851 38.971 48.915 ;
			RECT	39.107 48.851 39.139 48.915 ;
			RECT	39.275 48.851 39.307 48.915 ;
			RECT	39.443 48.851 39.475 48.915 ;
			RECT	39.611 48.851 39.643 48.915 ;
			RECT	39.779 48.851 39.811 48.915 ;
			RECT	39.947 48.851 39.979 48.915 ;
			RECT	40.115 48.851 40.147 48.915 ;
			RECT	40.283 48.851 40.315 48.915 ;
			RECT	40.451 48.851 40.483 48.915 ;
			RECT	40.619 48.851 40.651 48.915 ;
			RECT	40.787 48.851 40.819 48.915 ;
			RECT	40.955 48.851 40.987 48.915 ;
			RECT	41.123 48.851 41.155 48.915 ;
			RECT	41.291 48.851 41.323 48.915 ;
			RECT	41.459 48.851 41.491 48.915 ;
			RECT	41.627 48.851 41.659 48.915 ;
			RECT	41.795 48.851 41.827 48.915 ;
			RECT	41.963 48.851 41.995 48.915 ;
			RECT	42.131 48.851 42.163 48.915 ;
			RECT	42.299 48.851 42.331 48.915 ;
			RECT	42.467 48.851 42.499 48.915 ;
			RECT	42.635 48.851 42.667 48.915 ;
			RECT	42.803 48.851 42.835 48.915 ;
			RECT	42.971 48.851 43.003 48.915 ;
			RECT	43.139 48.851 43.171 48.915 ;
			RECT	43.307 48.851 43.339 48.915 ;
			RECT	43.475 48.851 43.507 48.915 ;
			RECT	43.643 48.851 43.675 48.915 ;
			RECT	43.811 48.851 43.843 48.915 ;
			RECT	43.979 48.851 44.011 48.915 ;
			RECT	44.147 48.851 44.179 48.915 ;
			RECT	44.315 48.851 44.347 48.915 ;
			RECT	44.483 48.851 44.515 48.915 ;
			RECT	44.651 48.851 44.683 48.915 ;
			RECT	44.819 48.851 44.851 48.915 ;
			RECT	44.987 48.851 45.019 48.915 ;
			RECT	45.155 48.851 45.187 48.915 ;
			RECT	45.323 48.851 45.355 48.915 ;
			RECT	45.491 48.851 45.523 48.915 ;
			RECT	45.659 48.851 45.691 48.915 ;
			RECT	45.827 48.851 45.859 48.915 ;
			RECT	45.995 48.851 46.027 48.915 ;
			RECT	46.163 48.851 46.195 48.915 ;
			RECT	46.331 48.851 46.363 48.915 ;
			RECT	46.499 48.851 46.531 48.915 ;
			RECT	46.667 48.851 46.699 48.915 ;
			RECT	46.835 48.851 46.867 48.915 ;
			RECT	47.003 48.851 47.035 48.915 ;
			RECT	47.171 48.851 47.203 48.915 ;
			RECT	47.339 48.851 47.371 48.915 ;
			RECT	47.507 48.851 47.539 48.915 ;
			RECT	47.675 48.851 47.707 48.915 ;
			RECT	47.843 48.851 47.875 48.915 ;
			RECT	48.011 48.851 48.043 48.915 ;
			RECT	48.179 48.851 48.211 48.915 ;
			RECT	48.347 48.851 48.379 48.915 ;
			RECT	48.515 48.851 48.547 48.915 ;
			RECT	48.683 48.851 48.715 48.915 ;
			RECT	48.851 48.851 48.883 48.915 ;
			RECT	49.019 48.851 49.051 48.915 ;
			RECT	49.311 48.851 49.375 48.915 ;
			RECT	49.566 48.851 49.598 48.915 ;
			RECT	52.03 48.851 52.062 48.915 ;
			RECT	52.578 48.851 52.61 48.915 ;
			RECT	52.976 48.854 53.008 48.918 ;
			RECT	53.91 48.851 53.942 48.915 ;
			RECT	54.251 48.851 54.283 48.915 ;
			RECT	54.812 48.851 54.844 48.915 ;
			RECT	55.562 48.867 55.626 48.899 ;
			RECT	55.803 48.851 55.835 48.915 ;
			RECT	55.969 48.851 56.033 48.915 ;
			RECT	57.844 48.851 57.876 48.915 ;
			RECT	58.606 48.851 58.638 48.915 ;
			RECT	58.829 48.851 58.893 48.915 ;
			RECT	59.153 48.851 59.185 48.915 ;
			RECT	59.321 48.851 59.353 48.915 ;
			RECT	59.489 48.851 59.521 48.915 ;
			RECT	59.657 48.851 59.689 48.915 ;
			RECT	59.825 48.851 59.857 48.915 ;
			RECT	59.993 48.851 60.025 48.915 ;
			RECT	60.161 48.851 60.193 48.915 ;
			RECT	60.329 48.851 60.361 48.915 ;
			RECT	60.497 48.851 60.529 48.915 ;
			RECT	60.665 48.851 60.697 48.915 ;
			RECT	60.833 48.851 60.865 48.915 ;
			RECT	61.001 48.851 61.033 48.915 ;
			RECT	61.169 48.851 61.201 48.915 ;
			RECT	61.337 48.851 61.369 48.915 ;
			RECT	61.505 48.851 61.537 48.915 ;
			RECT	61.673 48.851 61.705 48.915 ;
			RECT	61.841 48.851 61.873 48.915 ;
			RECT	62.009 48.851 62.041 48.915 ;
			RECT	62.177 48.851 62.209 48.915 ;
			RECT	62.345 48.851 62.377 48.915 ;
			RECT	62.513 48.851 62.545 48.915 ;
			RECT	62.681 48.851 62.713 48.915 ;
			RECT	62.849 48.851 62.881 48.915 ;
			RECT	63.017 48.851 63.049 48.915 ;
			RECT	63.185 48.851 63.217 48.915 ;
			RECT	63.353 48.851 63.385 48.915 ;
			RECT	63.521 48.851 63.553 48.915 ;
			RECT	63.689 48.851 63.721 48.915 ;
			RECT	63.857 48.851 63.889 48.915 ;
			RECT	64.025 48.851 64.057 48.915 ;
			RECT	64.193 48.851 64.225 48.915 ;
			RECT	64.361 48.851 64.393 48.915 ;
			RECT	64.529 48.851 64.561 48.915 ;
			RECT	64.697 48.851 64.729 48.915 ;
			RECT	64.865 48.851 64.897 48.915 ;
			RECT	65.033 48.851 65.065 48.915 ;
			RECT	65.201 48.851 65.233 48.915 ;
			RECT	65.369 48.851 65.401 48.915 ;
			RECT	65.537 48.851 65.569 48.915 ;
			RECT	65.705 48.851 65.737 48.915 ;
			RECT	65.873 48.851 65.905 48.915 ;
			RECT	66.041 48.851 66.073 48.915 ;
			RECT	66.209 48.851 66.241 48.915 ;
			RECT	66.377 48.851 66.409 48.915 ;
			RECT	66.545 48.851 66.577 48.915 ;
			RECT	66.713 48.851 66.745 48.915 ;
			RECT	66.881 48.851 66.913 48.915 ;
			RECT	67.049 48.851 67.081 48.915 ;
			RECT	67.217 48.851 67.249 48.915 ;
			RECT	67.385 48.851 67.417 48.915 ;
			RECT	67.553 48.851 67.585 48.915 ;
			RECT	67.721 48.851 67.753 48.915 ;
			RECT	67.889 48.851 67.921 48.915 ;
			RECT	68.057 48.851 68.089 48.915 ;
			RECT	68.225 48.851 68.257 48.915 ;
			RECT	68.393 48.851 68.425 48.915 ;
			RECT	68.561 48.851 68.593 48.915 ;
			RECT	68.729 48.851 68.761 48.915 ;
			RECT	68.897 48.851 68.929 48.915 ;
			RECT	69.065 48.851 69.097 48.915 ;
			RECT	69.233 48.851 69.265 48.915 ;
			RECT	69.401 48.851 69.433 48.915 ;
			RECT	69.569 48.851 69.601 48.915 ;
			RECT	69.737 48.851 69.769 48.915 ;
			RECT	69.905 48.851 69.937 48.915 ;
			RECT	70.073 48.851 70.105 48.915 ;
			RECT	70.241 48.851 70.273 48.915 ;
			RECT	70.409 48.851 70.441 48.915 ;
			RECT	70.577 48.851 70.609 48.915 ;
			RECT	70.745 48.851 70.777 48.915 ;
			RECT	70.913 48.851 70.945 48.915 ;
			RECT	71.081 48.851 71.113 48.915 ;
			RECT	71.249 48.851 71.281 48.915 ;
			RECT	71.417 48.851 71.449 48.915 ;
			RECT	71.585 48.851 71.617 48.915 ;
			RECT	71.753 48.851 71.785 48.915 ;
			RECT	71.921 48.851 71.953 48.915 ;
			RECT	72.089 48.851 72.121 48.915 ;
			RECT	72.257 48.851 72.289 48.915 ;
			RECT	72.425 48.851 72.457 48.915 ;
			RECT	72.593 48.851 72.625 48.915 ;
			RECT	72.761 48.851 72.793 48.915 ;
			RECT	72.929 48.851 72.961 48.915 ;
			RECT	73.097 48.851 73.129 48.915 ;
			RECT	73.265 48.851 73.297 48.915 ;
			RECT	73.433 48.851 73.465 48.915 ;
			RECT	73.601 48.851 73.633 48.915 ;
			RECT	73.769 48.851 73.801 48.915 ;
			RECT	73.937 48.851 73.969 48.915 ;
			RECT	74.105 48.851 74.137 48.915 ;
			RECT	74.273 48.851 74.305 48.915 ;
			RECT	74.441 48.851 74.473 48.915 ;
			RECT	74.609 48.851 74.641 48.915 ;
			RECT	74.777 48.851 74.809 48.915 ;
			RECT	74.945 48.851 74.977 48.915 ;
			RECT	75.113 48.851 75.145 48.915 ;
			RECT	75.281 48.851 75.313 48.915 ;
			RECT	75.449 48.851 75.481 48.915 ;
			RECT	75.617 48.851 75.649 48.915 ;
			RECT	75.785 48.851 75.817 48.915 ;
			RECT	75.953 48.851 75.985 48.915 ;
			RECT	76.121 48.851 76.153 48.915 ;
			RECT	76.289 48.851 76.321 48.915 ;
			RECT	76.457 48.851 76.489 48.915 ;
			RECT	76.625 48.851 76.657 48.915 ;
			RECT	76.793 48.851 76.825 48.915 ;
			RECT	76.961 48.851 76.993 48.915 ;
			RECT	77.129 48.851 77.161 48.915 ;
			RECT	77.297 48.851 77.329 48.915 ;
			RECT	77.465 48.851 77.497 48.915 ;
			RECT	77.633 48.851 77.665 48.915 ;
			RECT	77.801 48.851 77.833 48.915 ;
			RECT	77.969 48.851 78.001 48.915 ;
			RECT	78.137 48.851 78.169 48.915 ;
			RECT	78.305 48.851 78.337 48.915 ;
			RECT	78.473 48.851 78.505 48.915 ;
			RECT	78.641 48.851 78.673 48.915 ;
			RECT	78.809 48.851 78.841 48.915 ;
			RECT	78.977 48.851 79.009 48.915 ;
			RECT	79.145 48.851 79.177 48.915 ;
			RECT	79.313 48.851 79.345 48.915 ;
			RECT	79.481 48.851 79.513 48.915 ;
			RECT	79.649 48.851 79.681 48.915 ;
			RECT	79.817 48.851 79.849 48.915 ;
			RECT	79.985 48.851 80.017 48.915 ;
			RECT	80.153 48.851 80.185 48.915 ;
			RECT	80.321 48.851 80.353 48.915 ;
			RECT	80.657 48.851 80.689 48.915 ;
			RECT	80.993 48.851 81.025 48.915 ;
			RECT	81.329 48.851 81.361 48.915 ;
			RECT	81.665 48.851 81.697 48.915 ;
			RECT	82.001 48.851 82.033 48.915 ;
			RECT	82.337 48.851 82.369 48.915 ;
			RECT	82.673 48.851 82.705 48.915 ;
			RECT	83.009 48.851 83.041 48.915 ;
			RECT	83.345 48.851 83.377 48.915 ;
			RECT	83.681 48.851 83.713 48.915 ;
			RECT	84.017 48.851 84.049 48.915 ;
			RECT	84.353 48.851 84.385 48.915 ;
			RECT	84.689 48.851 84.721 48.915 ;
			RECT	85.025 48.851 85.057 48.915 ;
			RECT	85.361 48.851 85.393 48.915 ;
			RECT	85.697 48.851 85.729 48.915 ;
			RECT	86.033 48.851 86.065 48.915 ;
			RECT	86.369 48.851 86.401 48.915 ;
			RECT	86.705 48.851 86.737 48.915 ;
			RECT	87.041 48.851 87.073 48.915 ;
			RECT	87.377 48.851 87.409 48.915 ;
			RECT	87.713 48.851 87.745 48.915 ;
			RECT	88.049 48.851 88.081 48.915 ;
			RECT	88.385 48.851 88.417 48.915 ;
			RECT	88.721 48.851 88.753 48.915 ;
			RECT	89.057 48.851 89.089 48.915 ;
			RECT	89.393 48.851 89.425 48.915 ;
			RECT	89.729 48.851 89.761 48.915 ;
			RECT	90.065 48.851 90.097 48.915 ;
			RECT	90.401 48.851 90.433 48.915 ;
			RECT	90.737 48.851 90.769 48.915 ;
			RECT	91.073 48.851 91.105 48.915 ;
			RECT	91.409 48.851 91.441 48.915 ;
			RECT	91.745 48.851 91.777 48.915 ;
			RECT	92.081 48.851 92.113 48.915 ;
			RECT	92.417 48.851 92.449 48.915 ;
			RECT	92.753 48.851 92.785 48.915 ;
			RECT	93.089 48.851 93.121 48.915 ;
			RECT	93.425 48.851 93.457 48.915 ;
			RECT	93.761 48.851 93.793 48.915 ;
			RECT	94.097 48.851 94.129 48.915 ;
			RECT	94.433 48.851 94.465 48.915 ;
			RECT	94.769 48.851 94.801 48.915 ;
			RECT	95.105 48.851 95.137 48.915 ;
			RECT	95.441 48.851 95.473 48.915 ;
			RECT	95.777 48.851 95.809 48.915 ;
			RECT	96.113 48.851 96.145 48.915 ;
			RECT	96.449 48.851 96.481 48.915 ;
			RECT	96.785 48.851 96.817 48.915 ;
			RECT	97.121 48.851 97.153 48.915 ;
			RECT	97.457 48.851 97.489 48.915 ;
			RECT	97.793 48.851 97.825 48.915 ;
			RECT	98.129 48.851 98.161 48.915 ;
			RECT	98.465 48.851 98.497 48.915 ;
			RECT	98.801 48.851 98.833 48.915 ;
			RECT	99.137 48.851 99.169 48.915 ;
			RECT	99.473 48.851 99.505 48.915 ;
			RECT	99.809 48.851 99.841 48.915 ;
			RECT	100.145 48.851 100.177 48.915 ;
			RECT	100.481 48.851 100.513 48.915 ;
			RECT	100.817 48.851 100.849 48.915 ;
			RECT	101.153 48.851 101.185 48.915 ;
			RECT	101.489 48.851 101.521 48.915 ;
			RECT	101.825 48.851 101.857 48.915 ;
			RECT	102.077 48.851 102.109 48.915 ;
			RECT	102.363 48.851 102.395 48.915 ;
			RECT	102.995 48.851 103.027 48.915 ;
			RECT	103.175 48.851 103.207 48.915 ;
			RECT	103.807 48.851 103.839 48.915 ;
			RECT	104.093 48.851 104.125 48.915 ;
			RECT	104.345 48.851 104.377 48.915 ;
			RECT	104.681 48.851 104.713 48.915 ;
			RECT	105.017 48.851 105.049 48.915 ;
			RECT	105.353 48.851 105.385 48.915 ;
			RECT	105.689 48.851 105.721 48.915 ;
			RECT	106.025 48.851 106.057 48.915 ;
			RECT	106.361 48.851 106.393 48.915 ;
			RECT	106.697 48.851 106.729 48.915 ;
			RECT	107.033 48.851 107.065 48.915 ;
			RECT	107.369 48.851 107.401 48.915 ;
			RECT	107.705 48.851 107.737 48.915 ;
			RECT	108.041 48.851 108.073 48.915 ;
			RECT	108.377 48.851 108.409 48.915 ;
			RECT	108.713 48.851 108.745 48.915 ;
			RECT	109.049 48.851 109.081 48.915 ;
			RECT	109.385 48.851 109.417 48.915 ;
			RECT	109.721 48.851 109.753 48.915 ;
			RECT	110.057 48.851 110.089 48.915 ;
			RECT	110.393 48.851 110.425 48.915 ;
			RECT	110.729 48.851 110.761 48.915 ;
			RECT	111.065 48.851 111.097 48.915 ;
			RECT	111.401 48.851 111.433 48.915 ;
			RECT	111.737 48.851 111.769 48.915 ;
			RECT	112.073 48.851 112.105 48.915 ;
			RECT	112.409 48.851 112.441 48.915 ;
			RECT	112.745 48.851 112.777 48.915 ;
			RECT	113.081 48.851 113.113 48.915 ;
			RECT	113.417 48.851 113.449 48.915 ;
			RECT	113.753 48.851 113.785 48.915 ;
			RECT	114.089 48.851 114.121 48.915 ;
			RECT	114.425 48.851 114.457 48.915 ;
			RECT	114.761 48.851 114.793 48.915 ;
			RECT	115.097 48.851 115.129 48.915 ;
			RECT	115.433 48.851 115.465 48.915 ;
			RECT	115.769 48.851 115.801 48.915 ;
			RECT	116.105 48.851 116.137 48.915 ;
			RECT	116.441 48.851 116.473 48.915 ;
			RECT	116.777 48.851 116.809 48.915 ;
			RECT	117.113 48.851 117.145 48.915 ;
			RECT	117.449 48.851 117.481 48.915 ;
			RECT	117.785 48.851 117.817 48.915 ;
			RECT	118.121 48.851 118.153 48.915 ;
			RECT	118.457 48.851 118.489 48.915 ;
			RECT	118.793 48.851 118.825 48.915 ;
			RECT	119.129 48.851 119.161 48.915 ;
			RECT	119.465 48.851 119.497 48.915 ;
			RECT	119.801 48.851 119.833 48.915 ;
			RECT	120.137 48.851 120.169 48.915 ;
			RECT	120.473 48.851 120.505 48.915 ;
			RECT	120.809 48.851 120.841 48.915 ;
			RECT	121.145 48.851 121.177 48.915 ;
			RECT	121.481 48.851 121.513 48.915 ;
			RECT	121.817 48.851 121.849 48.915 ;
			RECT	122.153 48.851 122.185 48.915 ;
			RECT	122.489 48.851 122.521 48.915 ;
			RECT	122.825 48.851 122.857 48.915 ;
			RECT	123.161 48.851 123.193 48.915 ;
			RECT	123.497 48.851 123.529 48.915 ;
			RECT	123.833 48.851 123.865 48.915 ;
			RECT	124.169 48.851 124.201 48.915 ;
			RECT	124.505 48.851 124.537 48.915 ;
			RECT	124.841 48.851 124.873 48.915 ;
			RECT	125.177 48.851 125.209 48.915 ;
			RECT	125.513 48.851 125.545 48.915 ;
			RECT	125.849 48.851 125.881 48.915 ;
			RECT	126.017 48.851 126.049 48.915 ;
			RECT	126.185 48.851 126.217 48.915 ;
			RECT	126.353 48.851 126.385 48.915 ;
			RECT	126.521 48.851 126.553 48.915 ;
			RECT	126.689 48.851 126.721 48.915 ;
			RECT	126.857 48.851 126.889 48.915 ;
			RECT	127.025 48.851 127.057 48.915 ;
			RECT	127.193 48.851 127.225 48.915 ;
			RECT	127.361 48.851 127.393 48.915 ;
			RECT	127.529 48.851 127.561 48.915 ;
			RECT	127.697 48.851 127.729 48.915 ;
			RECT	127.865 48.851 127.897 48.915 ;
			RECT	128.033 48.851 128.065 48.915 ;
			RECT	128.201 48.851 128.233 48.915 ;
			RECT	128.369 48.851 128.401 48.915 ;
			RECT	128.537 48.851 128.569 48.915 ;
			RECT	128.705 48.851 128.737 48.915 ;
			RECT	128.873 48.851 128.905 48.915 ;
			RECT	129.041 48.851 129.073 48.915 ;
			RECT	129.209 48.851 129.241 48.915 ;
			RECT	129.377 48.851 129.409 48.915 ;
			RECT	129.545 48.851 129.577 48.915 ;
			RECT	129.713 48.851 129.745 48.915 ;
			RECT	129.881 48.851 129.913 48.915 ;
			RECT	130.049 48.851 130.081 48.915 ;
			RECT	130.217 48.851 130.249 48.915 ;
			RECT	130.385 48.851 130.417 48.915 ;
			RECT	130.553 48.851 130.585 48.915 ;
			RECT	130.721 48.851 130.753 48.915 ;
			RECT	130.889 48.851 130.921 48.915 ;
			RECT	131.057 48.851 131.089 48.915 ;
			RECT	131.225 48.851 131.257 48.915 ;
			RECT	131.393 48.851 131.425 48.915 ;
			RECT	131.561 48.851 131.593 48.915 ;
			RECT	131.729 48.851 131.761 48.915 ;
			RECT	131.897 48.851 131.929 48.915 ;
			RECT	132.065 48.851 132.097 48.915 ;
			RECT	132.233 48.851 132.265 48.915 ;
			RECT	132.401 48.851 132.433 48.915 ;
			RECT	132.569 48.851 132.601 48.915 ;
			RECT	132.737 48.851 132.769 48.915 ;
			RECT	132.905 48.851 132.937 48.915 ;
			RECT	133.073 48.851 133.105 48.915 ;
			RECT	133.241 48.851 133.273 48.915 ;
			RECT	133.409 48.851 133.441 48.915 ;
			RECT	133.577 48.851 133.609 48.915 ;
			RECT	133.745 48.851 133.777 48.915 ;
			RECT	133.913 48.851 133.945 48.915 ;
			RECT	134.081 48.851 134.113 48.915 ;
			RECT	134.249 48.851 134.281 48.915 ;
			RECT	134.417 48.851 134.449 48.915 ;
			RECT	134.585 48.851 134.617 48.915 ;
			RECT	134.753 48.851 134.785 48.915 ;
			RECT	134.921 48.851 134.953 48.915 ;
			RECT	135.089 48.851 135.121 48.915 ;
			RECT	135.257 48.851 135.289 48.915 ;
			RECT	135.425 48.851 135.457 48.915 ;
			RECT	135.593 48.851 135.625 48.915 ;
			RECT	135.761 48.851 135.793 48.915 ;
			RECT	135.929 48.851 135.961 48.915 ;
			RECT	136.097 48.851 136.129 48.915 ;
			RECT	136.265 48.851 136.297 48.915 ;
			RECT	136.433 48.851 136.465 48.915 ;
			RECT	136.601 48.851 136.633 48.915 ;
			RECT	136.769 48.851 136.801 48.915 ;
			RECT	136.937 48.851 136.969 48.915 ;
			RECT	137.105 48.851 137.137 48.915 ;
			RECT	137.273 48.851 137.305 48.915 ;
			RECT	137.441 48.851 137.473 48.915 ;
			RECT	137.609 48.851 137.641 48.915 ;
			RECT	137.777 48.851 137.809 48.915 ;
			RECT	137.945 48.851 137.977 48.915 ;
			RECT	138.113 48.851 138.145 48.915 ;
			RECT	138.281 48.851 138.313 48.915 ;
			RECT	138.449 48.851 138.481 48.915 ;
			RECT	138.617 48.851 138.649 48.915 ;
			RECT	138.785 48.851 138.817 48.915 ;
			RECT	138.953 48.851 138.985 48.915 ;
			RECT	139.121 48.851 139.153 48.915 ;
			RECT	139.289 48.851 139.321 48.915 ;
			RECT	139.457 48.851 139.489 48.915 ;
			RECT	139.625 48.851 139.657 48.915 ;
			RECT	139.793 48.851 139.825 48.915 ;
			RECT	139.961 48.851 139.993 48.915 ;
			RECT	140.129 48.851 140.161 48.915 ;
			RECT	140.297 48.851 140.329 48.915 ;
			RECT	140.465 48.851 140.497 48.915 ;
			RECT	140.633 48.851 140.665 48.915 ;
			RECT	140.801 48.851 140.833 48.915 ;
			RECT	140.969 48.851 141.001 48.915 ;
			RECT	141.137 48.851 141.169 48.915 ;
			RECT	141.305 48.851 141.337 48.915 ;
			RECT	141.473 48.851 141.505 48.915 ;
			RECT	141.641 48.851 141.673 48.915 ;
			RECT	141.809 48.851 141.841 48.915 ;
			RECT	141.977 48.851 142.009 48.915 ;
			RECT	142.145 48.851 142.177 48.915 ;
			RECT	142.313 48.851 142.345 48.915 ;
			RECT	142.481 48.851 142.513 48.915 ;
			RECT	142.649 48.851 142.681 48.915 ;
			RECT	142.817 48.851 142.849 48.915 ;
			RECT	142.985 48.851 143.017 48.915 ;
			RECT	143.153 48.851 143.185 48.915 ;
			RECT	143.321 48.851 143.353 48.915 ;
			RECT	143.489 48.851 143.521 48.915 ;
			RECT	143.657 48.851 143.689 48.915 ;
			RECT	143.825 48.851 143.857 48.915 ;
			RECT	143.993 48.851 144.025 48.915 ;
			RECT	144.161 48.851 144.193 48.915 ;
			RECT	144.329 48.851 144.361 48.915 ;
			RECT	144.497 48.851 144.529 48.915 ;
			RECT	144.665 48.851 144.697 48.915 ;
			RECT	144.833 48.851 144.865 48.915 ;
			RECT	145.001 48.851 145.033 48.915 ;
			RECT	145.169 48.851 145.201 48.915 ;
			RECT	145.337 48.851 145.369 48.915 ;
			RECT	145.505 48.851 145.537 48.915 ;
			RECT	145.673 48.851 145.705 48.915 ;
			RECT	145.841 48.851 145.873 48.915 ;
			RECT	146.009 48.851 146.041 48.915 ;
			RECT	146.177 48.851 146.209 48.915 ;
			RECT	146.345 48.851 146.377 48.915 ;
			RECT	146.513 48.851 146.545 48.915 ;
			RECT	146.681 48.851 146.713 48.915 ;
			RECT	146.849 48.851 146.881 48.915 ;
			RECT	147.017 48.851 147.049 48.915 ;
			RECT	147.309 48.851 147.373 48.915 ;
			RECT	147.564 48.851 147.596 48.915 ;
			RECT	150.028 48.851 150.06 48.915 ;
			RECT	150.576 48.851 150.608 48.915 ;
			RECT	150.974 48.854 151.006 48.918 ;
			RECT	151.908 48.851 151.94 48.915 ;
			RECT	152.249 48.851 152.281 48.915 ;
			RECT	152.81 48.851 152.842 48.915 ;
			RECT	153.56 48.867 153.624 48.899 ;
			RECT	153.801 48.851 153.833 48.915 ;
			RECT	153.967 48.851 154.031 48.915 ;
			RECT	155.842 48.851 155.874 48.915 ;
			RECT	156.604 48.851 156.636 48.915 ;
			RECT	156.827 48.851 156.891 48.915 ;
			RECT	157.151 48.851 157.183 48.915 ;
			RECT	157.319 48.851 157.351 48.915 ;
			RECT	157.487 48.851 157.519 48.915 ;
			RECT	157.655 48.851 157.687 48.915 ;
			RECT	157.823 48.851 157.855 48.915 ;
			RECT	157.991 48.851 158.023 48.915 ;
			RECT	158.159 48.851 158.191 48.915 ;
			RECT	158.327 48.851 158.359 48.915 ;
			RECT	158.495 48.851 158.527 48.915 ;
			RECT	158.663 48.851 158.695 48.915 ;
			RECT	158.831 48.851 158.863 48.915 ;
			RECT	158.999 48.851 159.031 48.915 ;
			RECT	159.167 48.851 159.199 48.915 ;
			RECT	159.335 48.851 159.367 48.915 ;
			RECT	159.503 48.851 159.535 48.915 ;
			RECT	159.671 48.851 159.703 48.915 ;
			RECT	159.839 48.851 159.871 48.915 ;
			RECT	160.007 48.851 160.039 48.915 ;
			RECT	160.175 48.851 160.207 48.915 ;
			RECT	160.343 48.851 160.375 48.915 ;
			RECT	160.511 48.851 160.543 48.915 ;
			RECT	160.679 48.851 160.711 48.915 ;
			RECT	160.847 48.851 160.879 48.915 ;
			RECT	161.015 48.851 161.047 48.915 ;
			RECT	161.183 48.851 161.215 48.915 ;
			RECT	161.351 48.851 161.383 48.915 ;
			RECT	161.519 48.851 161.551 48.915 ;
			RECT	161.687 48.851 161.719 48.915 ;
			RECT	161.855 48.851 161.887 48.915 ;
			RECT	162.023 48.851 162.055 48.915 ;
			RECT	162.191 48.851 162.223 48.915 ;
			RECT	162.359 48.851 162.391 48.915 ;
			RECT	162.527 48.851 162.559 48.915 ;
			RECT	162.695 48.851 162.727 48.915 ;
			RECT	162.863 48.851 162.895 48.915 ;
			RECT	163.031 48.851 163.063 48.915 ;
			RECT	163.199 48.851 163.231 48.915 ;
			RECT	163.367 48.851 163.399 48.915 ;
			RECT	163.535 48.851 163.567 48.915 ;
			RECT	163.703 48.851 163.735 48.915 ;
			RECT	163.871 48.851 163.903 48.915 ;
			RECT	164.039 48.851 164.071 48.915 ;
			RECT	164.207 48.851 164.239 48.915 ;
			RECT	164.375 48.851 164.407 48.915 ;
			RECT	164.543 48.851 164.575 48.915 ;
			RECT	164.711 48.851 164.743 48.915 ;
			RECT	164.879 48.851 164.911 48.915 ;
			RECT	165.047 48.851 165.079 48.915 ;
			RECT	165.215 48.851 165.247 48.915 ;
			RECT	165.383 48.851 165.415 48.915 ;
			RECT	165.551 48.851 165.583 48.915 ;
			RECT	165.719 48.851 165.751 48.915 ;
			RECT	165.887 48.851 165.919 48.915 ;
			RECT	166.055 48.851 166.087 48.915 ;
			RECT	166.223 48.851 166.255 48.915 ;
			RECT	166.391 48.851 166.423 48.915 ;
			RECT	166.559 48.851 166.591 48.915 ;
			RECT	166.727 48.851 166.759 48.915 ;
			RECT	166.895 48.851 166.927 48.915 ;
			RECT	167.063 48.851 167.095 48.915 ;
			RECT	167.231 48.851 167.263 48.915 ;
			RECT	167.399 48.851 167.431 48.915 ;
			RECT	167.567 48.851 167.599 48.915 ;
			RECT	167.735 48.851 167.767 48.915 ;
			RECT	167.903 48.851 167.935 48.915 ;
			RECT	168.071 48.851 168.103 48.915 ;
			RECT	168.239 48.851 168.271 48.915 ;
			RECT	168.407 48.851 168.439 48.915 ;
			RECT	168.575 48.851 168.607 48.915 ;
			RECT	168.743 48.851 168.775 48.915 ;
			RECT	168.911 48.851 168.943 48.915 ;
			RECT	169.079 48.851 169.111 48.915 ;
			RECT	169.247 48.851 169.279 48.915 ;
			RECT	169.415 48.851 169.447 48.915 ;
			RECT	169.583 48.851 169.615 48.915 ;
			RECT	169.751 48.851 169.783 48.915 ;
			RECT	169.919 48.851 169.951 48.915 ;
			RECT	170.087 48.851 170.119 48.915 ;
			RECT	170.255 48.851 170.287 48.915 ;
			RECT	170.423 48.851 170.455 48.915 ;
			RECT	170.591 48.851 170.623 48.915 ;
			RECT	170.759 48.851 170.791 48.915 ;
			RECT	170.927 48.851 170.959 48.915 ;
			RECT	171.095 48.851 171.127 48.915 ;
			RECT	171.263 48.851 171.295 48.915 ;
			RECT	171.431 48.851 171.463 48.915 ;
			RECT	171.599 48.851 171.631 48.915 ;
			RECT	171.767 48.851 171.799 48.915 ;
			RECT	171.935 48.851 171.967 48.915 ;
			RECT	172.103 48.851 172.135 48.915 ;
			RECT	172.271 48.851 172.303 48.915 ;
			RECT	172.439 48.851 172.471 48.915 ;
			RECT	172.607 48.851 172.639 48.915 ;
			RECT	172.775 48.851 172.807 48.915 ;
			RECT	172.943 48.851 172.975 48.915 ;
			RECT	173.111 48.851 173.143 48.915 ;
			RECT	173.279 48.851 173.311 48.915 ;
			RECT	173.447 48.851 173.479 48.915 ;
			RECT	173.615 48.851 173.647 48.915 ;
			RECT	173.783 48.851 173.815 48.915 ;
			RECT	173.951 48.851 173.983 48.915 ;
			RECT	174.119 48.851 174.151 48.915 ;
			RECT	174.287 48.851 174.319 48.915 ;
			RECT	174.455 48.851 174.487 48.915 ;
			RECT	174.623 48.851 174.655 48.915 ;
			RECT	174.791 48.851 174.823 48.915 ;
			RECT	174.959 48.851 174.991 48.915 ;
			RECT	175.127 48.851 175.159 48.915 ;
			RECT	175.295 48.851 175.327 48.915 ;
			RECT	175.463 48.851 175.495 48.915 ;
			RECT	175.631 48.851 175.663 48.915 ;
			RECT	175.799 48.851 175.831 48.915 ;
			RECT	175.967 48.851 175.999 48.915 ;
			RECT	176.135 48.851 176.167 48.915 ;
			RECT	176.303 48.851 176.335 48.915 ;
			RECT	176.471 48.851 176.503 48.915 ;
			RECT	176.639 48.851 176.671 48.915 ;
			RECT	176.807 48.851 176.839 48.915 ;
			RECT	176.975 48.851 177.007 48.915 ;
			RECT	177.143 48.851 177.175 48.915 ;
			RECT	177.311 48.851 177.343 48.915 ;
			RECT	177.479 48.851 177.511 48.915 ;
			RECT	177.647 48.851 177.679 48.915 ;
			RECT	177.815 48.851 177.847 48.915 ;
			RECT	177.983 48.851 178.015 48.915 ;
			RECT	178.151 48.851 178.183 48.915 ;
			RECT	178.319 48.851 178.351 48.915 ;
			RECT	178.655 48.851 178.687 48.915 ;
			RECT	178.991 48.851 179.023 48.915 ;
			RECT	179.327 48.851 179.359 48.915 ;
			RECT	179.663 48.851 179.695 48.915 ;
			RECT	179.999 48.851 180.031 48.915 ;
			RECT	180.335 48.851 180.367 48.915 ;
			RECT	180.671 48.851 180.703 48.915 ;
			RECT	181.007 48.851 181.039 48.915 ;
			RECT	181.343 48.851 181.375 48.915 ;
			RECT	181.679 48.851 181.711 48.915 ;
			RECT	182.015 48.851 182.047 48.915 ;
			RECT	182.351 48.851 182.383 48.915 ;
			RECT	182.687 48.851 182.719 48.915 ;
			RECT	183.023 48.851 183.055 48.915 ;
			RECT	183.359 48.851 183.391 48.915 ;
			RECT	183.695 48.851 183.727 48.915 ;
			RECT	184.031 48.851 184.063 48.915 ;
			RECT	184.367 48.851 184.399 48.915 ;
			RECT	184.703 48.851 184.735 48.915 ;
			RECT	185.039 48.851 185.071 48.915 ;
			RECT	185.375 48.851 185.407 48.915 ;
			RECT	185.711 48.851 185.743 48.915 ;
			RECT	186.047 48.851 186.079 48.915 ;
			RECT	186.383 48.851 186.415 48.915 ;
			RECT	186.719 48.851 186.751 48.915 ;
			RECT	187.055 48.851 187.087 48.915 ;
			RECT	187.391 48.851 187.423 48.915 ;
			RECT	187.727 48.851 187.759 48.915 ;
			RECT	188.063 48.851 188.095 48.915 ;
			RECT	188.399 48.851 188.431 48.915 ;
			RECT	188.735 48.851 188.767 48.915 ;
			RECT	189.071 48.851 189.103 48.915 ;
			RECT	189.407 48.851 189.439 48.915 ;
			RECT	189.743 48.851 189.775 48.915 ;
			RECT	190.079 48.851 190.111 48.915 ;
			RECT	190.415 48.851 190.447 48.915 ;
			RECT	190.751 48.851 190.783 48.915 ;
			RECT	191.087 48.851 191.119 48.915 ;
			RECT	191.423 48.851 191.455 48.915 ;
			RECT	191.759 48.851 191.791 48.915 ;
			RECT	192.095 48.851 192.127 48.915 ;
			RECT	192.431 48.851 192.463 48.915 ;
			RECT	192.767 48.851 192.799 48.915 ;
			RECT	193.103 48.851 193.135 48.915 ;
			RECT	193.439 48.851 193.471 48.915 ;
			RECT	193.775 48.851 193.807 48.915 ;
			RECT	194.111 48.851 194.143 48.915 ;
			RECT	194.447 48.851 194.479 48.915 ;
			RECT	194.783 48.851 194.815 48.915 ;
			RECT	195.119 48.851 195.151 48.915 ;
			RECT	195.455 48.851 195.487 48.915 ;
			RECT	195.791 48.851 195.823 48.915 ;
			RECT	196.127 48.851 196.159 48.915 ;
			RECT	196.463 48.851 196.495 48.915 ;
			RECT	196.799 48.851 196.831 48.915 ;
			RECT	197.135 48.851 197.167 48.915 ;
			RECT	197.471 48.851 197.503 48.915 ;
			RECT	197.807 48.851 197.839 48.915 ;
			RECT	198.143 48.851 198.175 48.915 ;
			RECT	198.479 48.851 198.511 48.915 ;
			RECT	198.815 48.851 198.847 48.915 ;
			RECT	199.151 48.851 199.183 48.915 ;
			RECT	199.487 48.851 199.519 48.915 ;
			RECT	199.823 48.851 199.855 48.915 ;
			RECT	200.075 48.851 200.107 48.915 ;
			RECT	200.361 48.851 200.393 48.915 ;
			RECT	201.403 48.851 201.435 48.915 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 49.42 201.665 49.51 ;
			LAYER	J3 ;
			RECT	0.755 49.433 0.787 49.497 ;
			RECT	1.164 49.433 1.196 49.497 ;
			RECT	1.645 49.449 1.709 49.481 ;
			RECT	2.339 49.433 2.371 49.497 ;
			RECT	3.438 49.433 3.47 49.497 ;
			RECT	4.195 49.433 4.227 49.497 ;
			RECT	4.944 49.449 5.008 49.481 ;
			RECT	6.347 49.433 6.379 49.497 ;
			RECT	6.683 49.433 6.715 49.497 ;
			RECT	7.019 49.433 7.051 49.497 ;
			RECT	7.355 49.433 7.387 49.497 ;
			RECT	7.691 49.433 7.723 49.497 ;
			RECT	8.027 49.433 8.059 49.497 ;
			RECT	8.363 49.433 8.395 49.497 ;
			RECT	8.699 49.433 8.731 49.497 ;
			RECT	9.035 49.433 9.067 49.497 ;
			RECT	9.371 49.433 9.403 49.497 ;
			RECT	9.707 49.433 9.739 49.497 ;
			RECT	10.043 49.433 10.075 49.497 ;
			RECT	10.379 49.433 10.411 49.497 ;
			RECT	10.715 49.433 10.747 49.497 ;
			RECT	11.051 49.433 11.083 49.497 ;
			RECT	11.387 49.433 11.419 49.497 ;
			RECT	11.723 49.433 11.755 49.497 ;
			RECT	12.059 49.433 12.091 49.497 ;
			RECT	12.395 49.433 12.427 49.497 ;
			RECT	12.731 49.433 12.763 49.497 ;
			RECT	13.067 49.433 13.099 49.497 ;
			RECT	13.403 49.433 13.435 49.497 ;
			RECT	13.739 49.433 13.771 49.497 ;
			RECT	14.075 49.433 14.107 49.497 ;
			RECT	14.411 49.433 14.443 49.497 ;
			RECT	14.747 49.433 14.779 49.497 ;
			RECT	15.083 49.433 15.115 49.497 ;
			RECT	15.419 49.433 15.451 49.497 ;
			RECT	15.755 49.433 15.787 49.497 ;
			RECT	16.091 49.433 16.123 49.497 ;
			RECT	16.427 49.433 16.459 49.497 ;
			RECT	16.763 49.433 16.795 49.497 ;
			RECT	17.099 49.433 17.131 49.497 ;
			RECT	17.435 49.433 17.467 49.497 ;
			RECT	17.771 49.433 17.803 49.497 ;
			RECT	18.107 49.433 18.139 49.497 ;
			RECT	18.443 49.433 18.475 49.497 ;
			RECT	18.779 49.433 18.811 49.497 ;
			RECT	19.115 49.433 19.147 49.497 ;
			RECT	19.451 49.433 19.483 49.497 ;
			RECT	19.787 49.433 19.819 49.497 ;
			RECT	20.123 49.433 20.155 49.497 ;
			RECT	20.459 49.433 20.491 49.497 ;
			RECT	20.795 49.433 20.827 49.497 ;
			RECT	21.131 49.433 21.163 49.497 ;
			RECT	21.467 49.433 21.499 49.497 ;
			RECT	21.803 49.433 21.835 49.497 ;
			RECT	22.139 49.433 22.171 49.497 ;
			RECT	22.475 49.433 22.507 49.497 ;
			RECT	22.811 49.433 22.843 49.497 ;
			RECT	23.147 49.433 23.179 49.497 ;
			RECT	23.483 49.433 23.515 49.497 ;
			RECT	23.819 49.433 23.851 49.497 ;
			RECT	24.155 49.433 24.187 49.497 ;
			RECT	24.491 49.433 24.523 49.497 ;
			RECT	24.827 49.433 24.859 49.497 ;
			RECT	25.163 49.433 25.195 49.497 ;
			RECT	25.499 49.433 25.531 49.497 ;
			RECT	25.835 49.433 25.867 49.497 ;
			RECT	26.171 49.433 26.203 49.497 ;
			RECT	26.507 49.433 26.539 49.497 ;
			RECT	26.843 49.433 26.875 49.497 ;
			RECT	27.179 49.433 27.211 49.497 ;
			RECT	27.515 49.433 27.547 49.497 ;
			RECT	49.327 49.433 49.359 49.497 ;
			RECT	52.124 49.433 52.156 49.497 ;
			RECT	52.578 49.433 52.61 49.497 ;
			RECT	53.148 49.433 53.18 49.497 ;
			RECT	54.251 49.433 54.283 49.497 ;
			RECT	55.578 49.433 55.61 49.497 ;
			RECT	55.803 49.433 55.835 49.497 ;
			RECT	57.844 49.433 57.876 49.497 ;
			RECT	58.845 49.433 58.877 49.497 ;
			RECT	80.657 49.433 80.689 49.497 ;
			RECT	80.993 49.433 81.025 49.497 ;
			RECT	81.329 49.433 81.361 49.497 ;
			RECT	81.665 49.433 81.697 49.497 ;
			RECT	82.001 49.433 82.033 49.497 ;
			RECT	82.337 49.433 82.369 49.497 ;
			RECT	82.673 49.433 82.705 49.497 ;
			RECT	83.009 49.433 83.041 49.497 ;
			RECT	83.345 49.433 83.377 49.497 ;
			RECT	83.681 49.433 83.713 49.497 ;
			RECT	84.017 49.433 84.049 49.497 ;
			RECT	84.353 49.433 84.385 49.497 ;
			RECT	84.689 49.433 84.721 49.497 ;
			RECT	85.025 49.433 85.057 49.497 ;
			RECT	85.361 49.433 85.393 49.497 ;
			RECT	85.697 49.433 85.729 49.497 ;
			RECT	86.033 49.433 86.065 49.497 ;
			RECT	86.369 49.433 86.401 49.497 ;
			RECT	86.705 49.433 86.737 49.497 ;
			RECT	87.041 49.433 87.073 49.497 ;
			RECT	87.377 49.433 87.409 49.497 ;
			RECT	87.713 49.433 87.745 49.497 ;
			RECT	88.049 49.433 88.081 49.497 ;
			RECT	88.385 49.433 88.417 49.497 ;
			RECT	88.721 49.433 88.753 49.497 ;
			RECT	89.057 49.433 89.089 49.497 ;
			RECT	89.393 49.433 89.425 49.497 ;
			RECT	89.729 49.433 89.761 49.497 ;
			RECT	90.065 49.433 90.097 49.497 ;
			RECT	90.401 49.433 90.433 49.497 ;
			RECT	90.737 49.433 90.769 49.497 ;
			RECT	91.073 49.433 91.105 49.497 ;
			RECT	91.409 49.433 91.441 49.497 ;
			RECT	91.745 49.433 91.777 49.497 ;
			RECT	92.081 49.433 92.113 49.497 ;
			RECT	92.417 49.433 92.449 49.497 ;
			RECT	92.753 49.433 92.785 49.497 ;
			RECT	93.089 49.433 93.121 49.497 ;
			RECT	93.425 49.433 93.457 49.497 ;
			RECT	93.761 49.433 93.793 49.497 ;
			RECT	94.097 49.433 94.129 49.497 ;
			RECT	94.433 49.433 94.465 49.497 ;
			RECT	94.769 49.433 94.801 49.497 ;
			RECT	95.105 49.433 95.137 49.497 ;
			RECT	95.441 49.433 95.473 49.497 ;
			RECT	95.777 49.433 95.809 49.497 ;
			RECT	96.113 49.433 96.145 49.497 ;
			RECT	96.449 49.433 96.481 49.497 ;
			RECT	96.785 49.433 96.817 49.497 ;
			RECT	97.121 49.433 97.153 49.497 ;
			RECT	97.457 49.433 97.489 49.497 ;
			RECT	97.793 49.433 97.825 49.497 ;
			RECT	98.129 49.433 98.161 49.497 ;
			RECT	98.465 49.433 98.497 49.497 ;
			RECT	98.801 49.433 98.833 49.497 ;
			RECT	99.137 49.433 99.169 49.497 ;
			RECT	99.473 49.433 99.505 49.497 ;
			RECT	99.809 49.433 99.841 49.497 ;
			RECT	100.145 49.433 100.177 49.497 ;
			RECT	100.481 49.433 100.513 49.497 ;
			RECT	100.817 49.433 100.849 49.497 ;
			RECT	101.153 49.433 101.185 49.497 ;
			RECT	101.489 49.433 101.521 49.497 ;
			RECT	101.825 49.433 101.857 49.497 ;
			RECT	104.345 49.433 104.377 49.497 ;
			RECT	104.681 49.433 104.713 49.497 ;
			RECT	105.017 49.433 105.049 49.497 ;
			RECT	105.353 49.433 105.385 49.497 ;
			RECT	105.689 49.433 105.721 49.497 ;
			RECT	106.025 49.433 106.057 49.497 ;
			RECT	106.361 49.433 106.393 49.497 ;
			RECT	106.697 49.433 106.729 49.497 ;
			RECT	107.033 49.433 107.065 49.497 ;
			RECT	107.369 49.433 107.401 49.497 ;
			RECT	107.705 49.433 107.737 49.497 ;
			RECT	108.041 49.433 108.073 49.497 ;
			RECT	108.377 49.433 108.409 49.497 ;
			RECT	108.713 49.433 108.745 49.497 ;
			RECT	109.049 49.433 109.081 49.497 ;
			RECT	109.385 49.433 109.417 49.497 ;
			RECT	109.721 49.433 109.753 49.497 ;
			RECT	110.057 49.433 110.089 49.497 ;
			RECT	110.393 49.433 110.425 49.497 ;
			RECT	110.729 49.433 110.761 49.497 ;
			RECT	111.065 49.433 111.097 49.497 ;
			RECT	111.401 49.433 111.433 49.497 ;
			RECT	111.737 49.433 111.769 49.497 ;
			RECT	112.073 49.433 112.105 49.497 ;
			RECT	112.409 49.433 112.441 49.497 ;
			RECT	112.745 49.433 112.777 49.497 ;
			RECT	113.081 49.433 113.113 49.497 ;
			RECT	113.417 49.433 113.449 49.497 ;
			RECT	113.753 49.433 113.785 49.497 ;
			RECT	114.089 49.433 114.121 49.497 ;
			RECT	114.425 49.433 114.457 49.497 ;
			RECT	114.761 49.433 114.793 49.497 ;
			RECT	115.097 49.433 115.129 49.497 ;
			RECT	115.433 49.433 115.465 49.497 ;
			RECT	115.769 49.433 115.801 49.497 ;
			RECT	116.105 49.433 116.137 49.497 ;
			RECT	116.441 49.433 116.473 49.497 ;
			RECT	116.777 49.433 116.809 49.497 ;
			RECT	117.113 49.433 117.145 49.497 ;
			RECT	117.449 49.433 117.481 49.497 ;
			RECT	117.785 49.433 117.817 49.497 ;
			RECT	118.121 49.433 118.153 49.497 ;
			RECT	118.457 49.433 118.489 49.497 ;
			RECT	118.793 49.433 118.825 49.497 ;
			RECT	119.129 49.433 119.161 49.497 ;
			RECT	119.465 49.433 119.497 49.497 ;
			RECT	119.801 49.433 119.833 49.497 ;
			RECT	120.137 49.433 120.169 49.497 ;
			RECT	120.473 49.433 120.505 49.497 ;
			RECT	120.809 49.433 120.841 49.497 ;
			RECT	121.145 49.433 121.177 49.497 ;
			RECT	121.481 49.433 121.513 49.497 ;
			RECT	121.817 49.433 121.849 49.497 ;
			RECT	122.153 49.433 122.185 49.497 ;
			RECT	122.489 49.433 122.521 49.497 ;
			RECT	122.825 49.433 122.857 49.497 ;
			RECT	123.161 49.433 123.193 49.497 ;
			RECT	123.497 49.433 123.529 49.497 ;
			RECT	123.833 49.433 123.865 49.497 ;
			RECT	124.169 49.433 124.201 49.497 ;
			RECT	124.505 49.433 124.537 49.497 ;
			RECT	124.841 49.433 124.873 49.497 ;
			RECT	125.177 49.433 125.209 49.497 ;
			RECT	125.513 49.433 125.545 49.497 ;
			RECT	147.325 49.433 147.357 49.497 ;
			RECT	150.122 49.433 150.154 49.497 ;
			RECT	150.576 49.433 150.608 49.497 ;
			RECT	151.146 49.433 151.178 49.497 ;
			RECT	152.249 49.433 152.281 49.497 ;
			RECT	153.576 49.433 153.608 49.497 ;
			RECT	153.801 49.433 153.833 49.497 ;
			RECT	155.842 49.433 155.874 49.497 ;
			RECT	156.843 49.433 156.875 49.497 ;
			RECT	178.655 49.433 178.687 49.497 ;
			RECT	178.991 49.433 179.023 49.497 ;
			RECT	179.327 49.433 179.359 49.497 ;
			RECT	179.663 49.433 179.695 49.497 ;
			RECT	179.999 49.433 180.031 49.497 ;
			RECT	180.335 49.433 180.367 49.497 ;
			RECT	180.671 49.433 180.703 49.497 ;
			RECT	181.007 49.433 181.039 49.497 ;
			RECT	181.343 49.433 181.375 49.497 ;
			RECT	181.679 49.433 181.711 49.497 ;
			RECT	182.015 49.433 182.047 49.497 ;
			RECT	182.351 49.433 182.383 49.497 ;
			RECT	182.687 49.433 182.719 49.497 ;
			RECT	183.023 49.433 183.055 49.497 ;
			RECT	183.359 49.433 183.391 49.497 ;
			RECT	183.695 49.433 183.727 49.497 ;
			RECT	184.031 49.433 184.063 49.497 ;
			RECT	184.367 49.433 184.399 49.497 ;
			RECT	184.703 49.433 184.735 49.497 ;
			RECT	185.039 49.433 185.071 49.497 ;
			RECT	185.375 49.433 185.407 49.497 ;
			RECT	185.711 49.433 185.743 49.497 ;
			RECT	186.047 49.433 186.079 49.497 ;
			RECT	186.383 49.433 186.415 49.497 ;
			RECT	186.719 49.433 186.751 49.497 ;
			RECT	187.055 49.433 187.087 49.497 ;
			RECT	187.391 49.433 187.423 49.497 ;
			RECT	187.727 49.433 187.759 49.497 ;
			RECT	188.063 49.433 188.095 49.497 ;
			RECT	188.399 49.433 188.431 49.497 ;
			RECT	188.735 49.433 188.767 49.497 ;
			RECT	189.071 49.433 189.103 49.497 ;
			RECT	189.407 49.433 189.439 49.497 ;
			RECT	189.743 49.433 189.775 49.497 ;
			RECT	190.079 49.433 190.111 49.497 ;
			RECT	190.415 49.433 190.447 49.497 ;
			RECT	190.751 49.433 190.783 49.497 ;
			RECT	191.087 49.433 191.119 49.497 ;
			RECT	191.423 49.433 191.455 49.497 ;
			RECT	191.759 49.433 191.791 49.497 ;
			RECT	192.095 49.433 192.127 49.497 ;
			RECT	192.431 49.433 192.463 49.497 ;
			RECT	192.767 49.433 192.799 49.497 ;
			RECT	193.103 49.433 193.135 49.497 ;
			RECT	193.439 49.433 193.471 49.497 ;
			RECT	193.775 49.433 193.807 49.497 ;
			RECT	194.111 49.433 194.143 49.497 ;
			RECT	194.447 49.433 194.479 49.497 ;
			RECT	194.783 49.433 194.815 49.497 ;
			RECT	195.119 49.433 195.151 49.497 ;
			RECT	195.455 49.433 195.487 49.497 ;
			RECT	195.791 49.433 195.823 49.497 ;
			RECT	196.127 49.433 196.159 49.497 ;
			RECT	196.463 49.433 196.495 49.497 ;
			RECT	196.799 49.433 196.831 49.497 ;
			RECT	197.135 49.433 197.167 49.497 ;
			RECT	197.471 49.433 197.503 49.497 ;
			RECT	197.807 49.433 197.839 49.497 ;
			RECT	198.143 49.433 198.175 49.497 ;
			RECT	198.479 49.433 198.511 49.497 ;
			RECT	198.815 49.433 198.847 49.497 ;
			RECT	199.151 49.433 199.183 49.497 ;
			RECT	199.487 49.433 199.519 49.497 ;
			RECT	199.823 49.433 199.855 49.497 ;
			RECT	201.403 49.433 201.435 49.497 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 49.818 201.665 49.928 ;
			LAYER	J3 ;
			RECT	1.645 49.841 1.709 49.905 ;
			RECT	2.339 49.841 2.371 49.905 ;
			RECT	3.438 49.841 3.47 49.905 ;
			RECT	4.195 49.841 4.227 49.905 ;
			RECT	4.944 49.841 5.008 49.905 ;
			RECT	6.347 49.841 6.379 49.905 ;
			RECT	6.683 49.841 6.715 49.905 ;
			RECT	7.019 49.841 7.051 49.905 ;
			RECT	7.355 49.841 7.387 49.905 ;
			RECT	7.691 49.841 7.723 49.905 ;
			RECT	8.027 49.841 8.059 49.905 ;
			RECT	8.363 49.841 8.395 49.905 ;
			RECT	8.699 49.841 8.731 49.905 ;
			RECT	9.035 49.841 9.067 49.905 ;
			RECT	9.371 49.841 9.403 49.905 ;
			RECT	9.707 49.841 9.739 49.905 ;
			RECT	10.043 49.841 10.075 49.905 ;
			RECT	10.379 49.841 10.411 49.905 ;
			RECT	10.715 49.841 10.747 49.905 ;
			RECT	11.051 49.841 11.083 49.905 ;
			RECT	11.387 49.841 11.419 49.905 ;
			RECT	11.723 49.841 11.755 49.905 ;
			RECT	12.059 49.841 12.091 49.905 ;
			RECT	12.395 49.841 12.427 49.905 ;
			RECT	12.731 49.841 12.763 49.905 ;
			RECT	13.067 49.841 13.099 49.905 ;
			RECT	13.403 49.841 13.435 49.905 ;
			RECT	13.739 49.841 13.771 49.905 ;
			RECT	14.075 49.841 14.107 49.905 ;
			RECT	14.411 49.841 14.443 49.905 ;
			RECT	14.747 49.841 14.779 49.905 ;
			RECT	15.083 49.841 15.115 49.905 ;
			RECT	15.419 49.841 15.451 49.905 ;
			RECT	15.755 49.841 15.787 49.905 ;
			RECT	16.091 49.841 16.123 49.905 ;
			RECT	16.427 49.841 16.459 49.905 ;
			RECT	16.763 49.841 16.795 49.905 ;
			RECT	17.099 49.841 17.131 49.905 ;
			RECT	17.435 49.841 17.467 49.905 ;
			RECT	17.771 49.841 17.803 49.905 ;
			RECT	18.107 49.841 18.139 49.905 ;
			RECT	18.443 49.841 18.475 49.905 ;
			RECT	18.779 49.841 18.811 49.905 ;
			RECT	19.115 49.841 19.147 49.905 ;
			RECT	19.451 49.841 19.483 49.905 ;
			RECT	19.787 49.841 19.819 49.905 ;
			RECT	20.123 49.841 20.155 49.905 ;
			RECT	20.459 49.841 20.491 49.905 ;
			RECT	20.795 49.841 20.827 49.905 ;
			RECT	21.131 49.841 21.163 49.905 ;
			RECT	21.467 49.841 21.499 49.905 ;
			RECT	21.803 49.841 21.835 49.905 ;
			RECT	22.139 49.841 22.171 49.905 ;
			RECT	22.475 49.841 22.507 49.905 ;
			RECT	22.811 49.841 22.843 49.905 ;
			RECT	23.147 49.841 23.179 49.905 ;
			RECT	23.483 49.841 23.515 49.905 ;
			RECT	23.819 49.841 23.851 49.905 ;
			RECT	24.155 49.841 24.187 49.905 ;
			RECT	24.491 49.841 24.523 49.905 ;
			RECT	24.827 49.841 24.859 49.905 ;
			RECT	25.163 49.841 25.195 49.905 ;
			RECT	25.499 49.841 25.531 49.905 ;
			RECT	25.835 49.841 25.867 49.905 ;
			RECT	26.171 49.841 26.203 49.905 ;
			RECT	26.507 49.841 26.539 49.905 ;
			RECT	26.843 49.841 26.875 49.905 ;
			RECT	27.179 49.841 27.211 49.905 ;
			RECT	27.515 49.841 27.547 49.905 ;
			RECT	49.311 49.841 49.375 49.905 ;
			RECT	52.124 49.857 52.156 49.889 ;
			RECT	52.578 49.841 52.61 49.905 ;
			RECT	53.132 49.841 53.196 49.905 ;
			RECT	54.251 49.841 54.283 49.905 ;
			RECT	55.562 49.841 55.626 49.905 ;
			RECT	55.803 49.841 55.835 49.905 ;
			RECT	57.255 49.841 57.287 49.905 ;
			RECT	58.829 49.841 58.893 49.905 ;
			RECT	80.657 49.841 80.689 49.905 ;
			RECT	80.993 49.841 81.025 49.905 ;
			RECT	81.329 49.841 81.361 49.905 ;
			RECT	81.665 49.841 81.697 49.905 ;
			RECT	82.001 49.841 82.033 49.905 ;
			RECT	82.337 49.841 82.369 49.905 ;
			RECT	82.673 49.841 82.705 49.905 ;
			RECT	83.009 49.841 83.041 49.905 ;
			RECT	83.345 49.841 83.377 49.905 ;
			RECT	83.681 49.841 83.713 49.905 ;
			RECT	84.017 49.841 84.049 49.905 ;
			RECT	84.353 49.841 84.385 49.905 ;
			RECT	84.689 49.841 84.721 49.905 ;
			RECT	85.025 49.841 85.057 49.905 ;
			RECT	85.361 49.841 85.393 49.905 ;
			RECT	85.697 49.841 85.729 49.905 ;
			RECT	86.033 49.841 86.065 49.905 ;
			RECT	86.369 49.841 86.401 49.905 ;
			RECT	86.705 49.841 86.737 49.905 ;
			RECT	87.041 49.841 87.073 49.905 ;
			RECT	87.377 49.841 87.409 49.905 ;
			RECT	87.713 49.841 87.745 49.905 ;
			RECT	88.049 49.841 88.081 49.905 ;
			RECT	88.385 49.841 88.417 49.905 ;
			RECT	88.721 49.841 88.753 49.905 ;
			RECT	89.057 49.841 89.089 49.905 ;
			RECT	89.393 49.841 89.425 49.905 ;
			RECT	89.729 49.841 89.761 49.905 ;
			RECT	90.065 49.841 90.097 49.905 ;
			RECT	90.401 49.841 90.433 49.905 ;
			RECT	90.737 49.841 90.769 49.905 ;
			RECT	91.073 49.841 91.105 49.905 ;
			RECT	91.409 49.841 91.441 49.905 ;
			RECT	91.745 49.841 91.777 49.905 ;
			RECT	92.081 49.841 92.113 49.905 ;
			RECT	92.417 49.841 92.449 49.905 ;
			RECT	92.753 49.841 92.785 49.905 ;
			RECT	93.089 49.841 93.121 49.905 ;
			RECT	93.425 49.841 93.457 49.905 ;
			RECT	93.761 49.841 93.793 49.905 ;
			RECT	94.097 49.841 94.129 49.905 ;
			RECT	94.433 49.841 94.465 49.905 ;
			RECT	94.769 49.841 94.801 49.905 ;
			RECT	95.105 49.841 95.137 49.905 ;
			RECT	95.441 49.841 95.473 49.905 ;
			RECT	95.777 49.841 95.809 49.905 ;
			RECT	96.113 49.841 96.145 49.905 ;
			RECT	96.449 49.841 96.481 49.905 ;
			RECT	96.785 49.841 96.817 49.905 ;
			RECT	97.121 49.841 97.153 49.905 ;
			RECT	97.457 49.841 97.489 49.905 ;
			RECT	97.793 49.841 97.825 49.905 ;
			RECT	98.129 49.841 98.161 49.905 ;
			RECT	98.465 49.841 98.497 49.905 ;
			RECT	98.801 49.841 98.833 49.905 ;
			RECT	99.137 49.841 99.169 49.905 ;
			RECT	99.473 49.841 99.505 49.905 ;
			RECT	99.809 49.841 99.841 49.905 ;
			RECT	100.145 49.841 100.177 49.905 ;
			RECT	100.481 49.841 100.513 49.905 ;
			RECT	100.817 49.841 100.849 49.905 ;
			RECT	101.153 49.841 101.185 49.905 ;
			RECT	101.489 49.841 101.521 49.905 ;
			RECT	101.825 49.841 101.857 49.905 ;
			RECT	104.345 49.841 104.377 49.905 ;
			RECT	104.681 49.841 104.713 49.905 ;
			RECT	105.017 49.841 105.049 49.905 ;
			RECT	105.353 49.841 105.385 49.905 ;
			RECT	105.689 49.841 105.721 49.905 ;
			RECT	106.025 49.841 106.057 49.905 ;
			RECT	106.361 49.841 106.393 49.905 ;
			RECT	106.697 49.841 106.729 49.905 ;
			RECT	107.033 49.841 107.065 49.905 ;
			RECT	107.369 49.841 107.401 49.905 ;
			RECT	107.705 49.841 107.737 49.905 ;
			RECT	108.041 49.841 108.073 49.905 ;
			RECT	108.377 49.841 108.409 49.905 ;
			RECT	108.713 49.841 108.745 49.905 ;
			RECT	109.049 49.841 109.081 49.905 ;
			RECT	109.385 49.841 109.417 49.905 ;
			RECT	109.721 49.841 109.753 49.905 ;
			RECT	110.057 49.841 110.089 49.905 ;
			RECT	110.393 49.841 110.425 49.905 ;
			RECT	110.729 49.841 110.761 49.905 ;
			RECT	111.065 49.841 111.097 49.905 ;
			RECT	111.401 49.841 111.433 49.905 ;
			RECT	111.737 49.841 111.769 49.905 ;
			RECT	112.073 49.841 112.105 49.905 ;
			RECT	112.409 49.841 112.441 49.905 ;
			RECT	112.745 49.841 112.777 49.905 ;
			RECT	113.081 49.841 113.113 49.905 ;
			RECT	113.417 49.841 113.449 49.905 ;
			RECT	113.753 49.841 113.785 49.905 ;
			RECT	114.089 49.841 114.121 49.905 ;
			RECT	114.425 49.841 114.457 49.905 ;
			RECT	114.761 49.841 114.793 49.905 ;
			RECT	115.097 49.841 115.129 49.905 ;
			RECT	115.433 49.841 115.465 49.905 ;
			RECT	115.769 49.841 115.801 49.905 ;
			RECT	116.105 49.841 116.137 49.905 ;
			RECT	116.441 49.841 116.473 49.905 ;
			RECT	116.777 49.841 116.809 49.905 ;
			RECT	117.113 49.841 117.145 49.905 ;
			RECT	117.449 49.841 117.481 49.905 ;
			RECT	117.785 49.841 117.817 49.905 ;
			RECT	118.121 49.841 118.153 49.905 ;
			RECT	118.457 49.841 118.489 49.905 ;
			RECT	118.793 49.841 118.825 49.905 ;
			RECT	119.129 49.841 119.161 49.905 ;
			RECT	119.465 49.841 119.497 49.905 ;
			RECT	119.801 49.841 119.833 49.905 ;
			RECT	120.137 49.841 120.169 49.905 ;
			RECT	120.473 49.841 120.505 49.905 ;
			RECT	120.809 49.841 120.841 49.905 ;
			RECT	121.145 49.841 121.177 49.905 ;
			RECT	121.481 49.841 121.513 49.905 ;
			RECT	121.817 49.841 121.849 49.905 ;
			RECT	122.153 49.841 122.185 49.905 ;
			RECT	122.489 49.841 122.521 49.905 ;
			RECT	122.825 49.841 122.857 49.905 ;
			RECT	123.161 49.841 123.193 49.905 ;
			RECT	123.497 49.841 123.529 49.905 ;
			RECT	123.833 49.841 123.865 49.905 ;
			RECT	124.169 49.841 124.201 49.905 ;
			RECT	124.505 49.841 124.537 49.905 ;
			RECT	124.841 49.841 124.873 49.905 ;
			RECT	125.177 49.841 125.209 49.905 ;
			RECT	125.513 49.841 125.545 49.905 ;
			RECT	147.309 49.841 147.373 49.905 ;
			RECT	150.122 49.857 150.154 49.889 ;
			RECT	150.576 49.841 150.608 49.905 ;
			RECT	151.13 49.841 151.194 49.905 ;
			RECT	152.249 49.841 152.281 49.905 ;
			RECT	153.56 49.841 153.624 49.905 ;
			RECT	153.801 49.841 153.833 49.905 ;
			RECT	155.253 49.841 155.285 49.905 ;
			RECT	156.827 49.841 156.891 49.905 ;
			RECT	178.655 49.841 178.687 49.905 ;
			RECT	178.991 49.841 179.023 49.905 ;
			RECT	179.327 49.841 179.359 49.905 ;
			RECT	179.663 49.841 179.695 49.905 ;
			RECT	179.999 49.841 180.031 49.905 ;
			RECT	180.335 49.841 180.367 49.905 ;
			RECT	180.671 49.841 180.703 49.905 ;
			RECT	181.007 49.841 181.039 49.905 ;
			RECT	181.343 49.841 181.375 49.905 ;
			RECT	181.679 49.841 181.711 49.905 ;
			RECT	182.015 49.841 182.047 49.905 ;
			RECT	182.351 49.841 182.383 49.905 ;
			RECT	182.687 49.841 182.719 49.905 ;
			RECT	183.023 49.841 183.055 49.905 ;
			RECT	183.359 49.841 183.391 49.905 ;
			RECT	183.695 49.841 183.727 49.905 ;
			RECT	184.031 49.841 184.063 49.905 ;
			RECT	184.367 49.841 184.399 49.905 ;
			RECT	184.703 49.841 184.735 49.905 ;
			RECT	185.039 49.841 185.071 49.905 ;
			RECT	185.375 49.841 185.407 49.905 ;
			RECT	185.711 49.841 185.743 49.905 ;
			RECT	186.047 49.841 186.079 49.905 ;
			RECT	186.383 49.841 186.415 49.905 ;
			RECT	186.719 49.841 186.751 49.905 ;
			RECT	187.055 49.841 187.087 49.905 ;
			RECT	187.391 49.841 187.423 49.905 ;
			RECT	187.727 49.841 187.759 49.905 ;
			RECT	188.063 49.841 188.095 49.905 ;
			RECT	188.399 49.841 188.431 49.905 ;
			RECT	188.735 49.841 188.767 49.905 ;
			RECT	189.071 49.841 189.103 49.905 ;
			RECT	189.407 49.841 189.439 49.905 ;
			RECT	189.743 49.841 189.775 49.905 ;
			RECT	190.079 49.841 190.111 49.905 ;
			RECT	190.415 49.841 190.447 49.905 ;
			RECT	190.751 49.841 190.783 49.905 ;
			RECT	191.087 49.841 191.119 49.905 ;
			RECT	191.423 49.841 191.455 49.905 ;
			RECT	191.759 49.841 191.791 49.905 ;
			RECT	192.095 49.841 192.127 49.905 ;
			RECT	192.431 49.841 192.463 49.905 ;
			RECT	192.767 49.841 192.799 49.905 ;
			RECT	193.103 49.841 193.135 49.905 ;
			RECT	193.439 49.841 193.471 49.905 ;
			RECT	193.775 49.841 193.807 49.905 ;
			RECT	194.111 49.841 194.143 49.905 ;
			RECT	194.447 49.841 194.479 49.905 ;
			RECT	194.783 49.841 194.815 49.905 ;
			RECT	195.119 49.841 195.151 49.905 ;
			RECT	195.455 49.841 195.487 49.905 ;
			RECT	195.791 49.841 195.823 49.905 ;
			RECT	196.127 49.841 196.159 49.905 ;
			RECT	196.463 49.841 196.495 49.905 ;
			RECT	196.799 49.841 196.831 49.905 ;
			RECT	197.135 49.841 197.167 49.905 ;
			RECT	197.471 49.841 197.503 49.905 ;
			RECT	197.807 49.841 197.839 49.905 ;
			RECT	198.143 49.841 198.175 49.905 ;
			RECT	198.479 49.841 198.511 49.905 ;
			RECT	198.815 49.841 198.847 49.905 ;
			RECT	199.151 49.841 199.183 49.905 ;
			RECT	199.487 49.841 199.519 49.905 ;
			RECT	199.823 49.841 199.855 49.905 ;
			RECT	201.403 49.841 201.435 49.905 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 50.528 201.665 50.638 ;
			LAYER	J3 ;
			RECT	0.755 50.551 0.787 50.615 ;
			RECT	1.164 50.551 1.196 50.615 ;
			RECT	1.645 50.551 1.709 50.615 ;
			RECT	2.339 50.551 2.371 50.615 ;
			RECT	3.438 50.551 3.47 50.615 ;
			RECT	3.585 50.551 3.617 50.615 ;
			RECT	4.195 50.551 4.227 50.615 ;
			RECT	4.944 50.551 5.008 50.615 ;
			RECT	5.409 50.551 5.441 50.615 ;
			RECT	49.311 50.551 49.375 50.615 ;
			RECT	52.124 50.567 52.156 50.599 ;
			RECT	52.578 50.551 52.61 50.615 ;
			RECT	53.132 50.551 53.196 50.615 ;
			RECT	54.251 50.551 54.283 50.615 ;
			RECT	55.562 50.567 55.626 50.599 ;
			RECT	55.803 50.551 55.835 50.615 ;
			RECT	57.255 50.551 57.287 50.615 ;
			RECT	58.829 50.551 58.893 50.615 ;
			RECT	102.763 50.551 102.795 50.615 ;
			RECT	102.995 50.551 103.027 50.615 ;
			RECT	103.175 50.551 103.207 50.615 ;
			RECT	103.407 50.551 103.439 50.615 ;
			RECT	147.309 50.551 147.373 50.615 ;
			RECT	150.122 50.567 150.154 50.599 ;
			RECT	150.576 50.551 150.608 50.615 ;
			RECT	151.13 50.551 151.194 50.615 ;
			RECT	152.249 50.551 152.281 50.615 ;
			RECT	153.56 50.567 153.624 50.599 ;
			RECT	153.801 50.551 153.833 50.615 ;
			RECT	155.253 50.551 155.285 50.615 ;
			RECT	156.827 50.551 156.891 50.615 ;
			RECT	200.761 50.551 200.793 50.615 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 79.526 201.665 79.636 ;
			LAYER	J3 ;
			RECT	0.756 79.549 0.788 79.613 ;
			RECT	1.645 79.549 1.709 79.613 ;
			RECT	2.323 79.549 2.387 79.613 ;
			RECT	3.438 79.549 3.47 79.613 ;
			RECT	3.585 79.549 3.617 79.613 ;
			RECT	4.195 79.549 4.227 79.613 ;
			RECT	4.704 79.565 4.768 79.597 ;
			RECT	4.944 79.549 5.008 79.613 ;
			RECT	52.124 79.565 52.156 79.597 ;
			RECT	52.577 79.565 52.609 79.597 ;
			RECT	53.132 79.549 53.196 79.613 ;
			RECT	54.246 79.565 54.278 79.597 ;
			RECT	55.554 79.549 55.618 79.613 ;
			RECT	55.807 79.549 55.839 79.613 ;
			RECT	102.995 79.549 103.027 79.613 ;
			RECT	103.175 79.549 103.207 79.613 ;
			RECT	150.122 79.565 150.154 79.597 ;
			RECT	150.575 79.565 150.607 79.597 ;
			RECT	151.13 79.549 151.194 79.613 ;
			RECT	152.244 79.565 152.276 79.597 ;
			RECT	153.552 79.549 153.616 79.613 ;
			RECT	153.805 79.549 153.837 79.613 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 77.606 201.665 77.716 ;
			LAYER	J3 ;
			RECT	0.756 77.629 0.788 77.693 ;
			RECT	1.645 77.629 1.709 77.693 ;
			RECT	2.323 77.629 2.387 77.693 ;
			RECT	3.438 77.629 3.47 77.693 ;
			RECT	3.585 77.629 3.617 77.693 ;
			RECT	4.195 77.629 4.227 77.693 ;
			RECT	4.704 77.645 4.768 77.677 ;
			RECT	4.944 77.629 5.008 77.693 ;
			RECT	52.124 77.645 52.156 77.677 ;
			RECT	52.577 77.645 52.609 77.677 ;
			RECT	53.132 77.629 53.196 77.693 ;
			RECT	54.246 77.645 54.278 77.677 ;
			RECT	55.554 77.629 55.618 77.693 ;
			RECT	55.807 77.629 55.839 77.693 ;
			RECT	102.995 77.629 103.027 77.693 ;
			RECT	103.175 77.629 103.207 77.693 ;
			RECT	150.122 77.645 150.154 77.677 ;
			RECT	150.575 77.645 150.607 77.677 ;
			RECT	151.13 77.629 151.194 77.693 ;
			RECT	152.244 77.645 152.276 77.677 ;
			RECT	153.552 77.629 153.616 77.693 ;
			RECT	153.805 77.629 153.837 77.693 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 31.34 201.665 31.45 ;
			LAYER	J3 ;
			RECT	0.756 31.363 0.788 31.427 ;
			RECT	1.645 31.363 1.709 31.427 ;
			RECT	2.323 31.363 2.387 31.427 ;
			RECT	3.438 31.363 3.47 31.427 ;
			RECT	3.585 31.363 3.617 31.427 ;
			RECT	4.195 31.363 4.227 31.427 ;
			RECT	4.704 31.379 4.768 31.411 ;
			RECT	4.944 31.363 5.008 31.427 ;
			RECT	52.124 31.379 52.156 31.411 ;
			RECT	52.577 31.379 52.609 31.411 ;
			RECT	53.132 31.363 53.196 31.427 ;
			RECT	54.246 31.379 54.278 31.411 ;
			RECT	55.554 31.363 55.618 31.427 ;
			RECT	55.807 31.363 55.839 31.427 ;
			RECT	102.995 31.363 103.027 31.427 ;
			RECT	103.175 31.363 103.207 31.427 ;
			RECT	150.122 31.379 150.154 31.411 ;
			RECT	150.575 31.379 150.607 31.411 ;
			RECT	151.13 31.363 151.194 31.427 ;
			RECT	152.244 31.379 152.276 31.411 ;
			RECT	153.552 31.363 153.616 31.427 ;
			RECT	153.805 31.363 153.837 31.427 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 29.42 201.665 29.53 ;
			LAYER	J3 ;
			RECT	0.756 29.443 0.788 29.507 ;
			RECT	1.645 29.443 1.709 29.507 ;
			RECT	2.323 29.443 2.387 29.507 ;
			RECT	3.438 29.443 3.47 29.507 ;
			RECT	3.585 29.443 3.617 29.507 ;
			RECT	4.195 29.443 4.227 29.507 ;
			RECT	4.704 29.459 4.768 29.491 ;
			RECT	4.944 29.443 5.008 29.507 ;
			RECT	52.124 29.459 52.156 29.491 ;
			RECT	52.577 29.459 52.609 29.491 ;
			RECT	53.132 29.443 53.196 29.507 ;
			RECT	54.246 29.459 54.278 29.491 ;
			RECT	55.554 29.443 55.618 29.507 ;
			RECT	55.807 29.443 55.839 29.507 ;
			RECT	102.995 29.443 103.027 29.507 ;
			RECT	103.175 29.443 103.207 29.507 ;
			RECT	150.122 29.459 150.154 29.491 ;
			RECT	150.575 29.459 150.607 29.491 ;
			RECT	151.13 29.443 151.194 29.507 ;
			RECT	152.244 29.459 152.276 29.491 ;
			RECT	153.552 29.443 153.616 29.507 ;
			RECT	153.805 29.443 153.837 29.507 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 27.5 201.665 27.61 ;
			LAYER	J3 ;
			RECT	0.756 27.523 0.788 27.587 ;
			RECT	1.645 27.523 1.709 27.587 ;
			RECT	2.323 27.523 2.387 27.587 ;
			RECT	3.438 27.523 3.47 27.587 ;
			RECT	3.585 27.523 3.617 27.587 ;
			RECT	4.195 27.523 4.227 27.587 ;
			RECT	4.704 27.539 4.768 27.571 ;
			RECT	4.944 27.523 5.008 27.587 ;
			RECT	52.124 27.539 52.156 27.571 ;
			RECT	52.577 27.539 52.609 27.571 ;
			RECT	53.132 27.523 53.196 27.587 ;
			RECT	54.246 27.539 54.278 27.571 ;
			RECT	55.554 27.523 55.618 27.587 ;
			RECT	55.807 27.523 55.839 27.587 ;
			RECT	102.995 27.523 103.027 27.587 ;
			RECT	103.175 27.523 103.207 27.587 ;
			RECT	150.122 27.539 150.154 27.571 ;
			RECT	150.575 27.539 150.607 27.571 ;
			RECT	151.13 27.523 151.194 27.587 ;
			RECT	152.244 27.539 152.276 27.571 ;
			RECT	153.552 27.523 153.616 27.587 ;
			RECT	153.805 27.523 153.837 27.587 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 25.58 201.665 25.69 ;
			LAYER	J3 ;
			RECT	0.756 25.603 0.788 25.667 ;
			RECT	1.645 25.603 1.709 25.667 ;
			RECT	2.323 25.603 2.387 25.667 ;
			RECT	3.438 25.603 3.47 25.667 ;
			RECT	3.585 25.603 3.617 25.667 ;
			RECT	4.195 25.603 4.227 25.667 ;
			RECT	4.704 25.619 4.768 25.651 ;
			RECT	4.944 25.603 5.008 25.667 ;
			RECT	52.124 25.619 52.156 25.651 ;
			RECT	52.577 25.619 52.609 25.651 ;
			RECT	53.132 25.603 53.196 25.667 ;
			RECT	54.246 25.619 54.278 25.651 ;
			RECT	55.554 25.603 55.618 25.667 ;
			RECT	55.807 25.603 55.839 25.667 ;
			RECT	102.995 25.603 103.027 25.667 ;
			RECT	103.175 25.603 103.207 25.667 ;
			RECT	150.122 25.619 150.154 25.651 ;
			RECT	150.575 25.619 150.607 25.651 ;
			RECT	151.13 25.603 151.194 25.667 ;
			RECT	152.244 25.619 152.276 25.651 ;
			RECT	153.552 25.603 153.616 25.667 ;
			RECT	153.805 25.603 153.837 25.667 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 23.66 201.665 23.77 ;
			LAYER	J3 ;
			RECT	0.756 23.683 0.788 23.747 ;
			RECT	1.645 23.683 1.709 23.747 ;
			RECT	2.323 23.683 2.387 23.747 ;
			RECT	3.438 23.683 3.47 23.747 ;
			RECT	3.585 23.683 3.617 23.747 ;
			RECT	4.195 23.683 4.227 23.747 ;
			RECT	4.704 23.699 4.768 23.731 ;
			RECT	4.944 23.683 5.008 23.747 ;
			RECT	52.124 23.699 52.156 23.731 ;
			RECT	52.577 23.699 52.609 23.731 ;
			RECT	53.132 23.683 53.196 23.747 ;
			RECT	54.246 23.699 54.278 23.731 ;
			RECT	55.554 23.683 55.618 23.747 ;
			RECT	55.807 23.683 55.839 23.747 ;
			RECT	102.995 23.683 103.027 23.747 ;
			RECT	103.175 23.683 103.207 23.747 ;
			RECT	150.122 23.699 150.154 23.731 ;
			RECT	150.575 23.699 150.607 23.731 ;
			RECT	151.13 23.683 151.194 23.747 ;
			RECT	152.244 23.699 152.276 23.731 ;
			RECT	153.552 23.683 153.616 23.747 ;
			RECT	153.805 23.683 153.837 23.747 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 75.686 201.665 75.796 ;
			LAYER	J3 ;
			RECT	0.756 75.709 0.788 75.773 ;
			RECT	1.645 75.709 1.709 75.773 ;
			RECT	2.323 75.709 2.387 75.773 ;
			RECT	3.438 75.709 3.47 75.773 ;
			RECT	3.585 75.709 3.617 75.773 ;
			RECT	4.195 75.709 4.227 75.773 ;
			RECT	4.704 75.725 4.768 75.757 ;
			RECT	4.944 75.709 5.008 75.773 ;
			RECT	52.124 75.725 52.156 75.757 ;
			RECT	52.577 75.725 52.609 75.757 ;
			RECT	53.132 75.709 53.196 75.773 ;
			RECT	54.246 75.725 54.278 75.757 ;
			RECT	55.554 75.709 55.618 75.773 ;
			RECT	55.807 75.709 55.839 75.773 ;
			RECT	102.995 75.709 103.027 75.773 ;
			RECT	103.175 75.709 103.207 75.773 ;
			RECT	150.122 75.725 150.154 75.757 ;
			RECT	150.575 75.725 150.607 75.757 ;
			RECT	151.13 75.709 151.194 75.773 ;
			RECT	152.244 75.725 152.276 75.757 ;
			RECT	153.552 75.709 153.616 75.773 ;
			RECT	153.805 75.709 153.837 75.773 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 21.74 201.665 21.85 ;
			LAYER	J3 ;
			RECT	0.756 21.763 0.788 21.827 ;
			RECT	1.645 21.763 1.709 21.827 ;
			RECT	2.323 21.763 2.387 21.827 ;
			RECT	3.438 21.763 3.47 21.827 ;
			RECT	3.585 21.763 3.617 21.827 ;
			RECT	4.195 21.763 4.227 21.827 ;
			RECT	4.704 21.779 4.768 21.811 ;
			RECT	4.944 21.763 5.008 21.827 ;
			RECT	52.124 21.779 52.156 21.811 ;
			RECT	52.577 21.779 52.609 21.811 ;
			RECT	53.132 21.763 53.196 21.827 ;
			RECT	54.246 21.779 54.278 21.811 ;
			RECT	55.554 21.763 55.618 21.827 ;
			RECT	55.807 21.763 55.839 21.827 ;
			RECT	102.995 21.763 103.027 21.827 ;
			RECT	103.175 21.763 103.207 21.827 ;
			RECT	150.122 21.779 150.154 21.811 ;
			RECT	150.575 21.779 150.607 21.811 ;
			RECT	151.13 21.763 151.194 21.827 ;
			RECT	152.244 21.779 152.276 21.811 ;
			RECT	153.552 21.763 153.616 21.827 ;
			RECT	153.805 21.763 153.837 21.827 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 19.82 201.665 19.93 ;
			LAYER	J3 ;
			RECT	0.756 19.843 0.788 19.907 ;
			RECT	1.645 19.843 1.709 19.907 ;
			RECT	2.323 19.843 2.387 19.907 ;
			RECT	3.438 19.843 3.47 19.907 ;
			RECT	3.585 19.843 3.617 19.907 ;
			RECT	4.195 19.843 4.227 19.907 ;
			RECT	4.704 19.859 4.768 19.891 ;
			RECT	4.944 19.843 5.008 19.907 ;
			RECT	52.124 19.859 52.156 19.891 ;
			RECT	52.577 19.859 52.609 19.891 ;
			RECT	53.132 19.843 53.196 19.907 ;
			RECT	54.246 19.859 54.278 19.891 ;
			RECT	55.554 19.843 55.618 19.907 ;
			RECT	55.807 19.843 55.839 19.907 ;
			RECT	102.995 19.843 103.027 19.907 ;
			RECT	103.175 19.843 103.207 19.907 ;
			RECT	150.122 19.859 150.154 19.891 ;
			RECT	150.575 19.859 150.607 19.891 ;
			RECT	151.13 19.843 151.194 19.907 ;
			RECT	152.244 19.859 152.276 19.891 ;
			RECT	153.552 19.843 153.616 19.907 ;
			RECT	153.805 19.843 153.837 19.907 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 17.9 201.665 18.01 ;
			LAYER	J3 ;
			RECT	0.756 17.923 0.788 17.987 ;
			RECT	1.645 17.923 1.709 17.987 ;
			RECT	2.323 17.923 2.387 17.987 ;
			RECT	3.438 17.923 3.47 17.987 ;
			RECT	3.585 17.923 3.617 17.987 ;
			RECT	4.195 17.923 4.227 17.987 ;
			RECT	4.704 17.939 4.768 17.971 ;
			RECT	4.944 17.923 5.008 17.987 ;
			RECT	52.124 17.939 52.156 17.971 ;
			RECT	52.577 17.939 52.609 17.971 ;
			RECT	53.132 17.923 53.196 17.987 ;
			RECT	54.246 17.939 54.278 17.971 ;
			RECT	55.554 17.923 55.618 17.987 ;
			RECT	55.807 17.923 55.839 17.987 ;
			RECT	102.995 17.923 103.027 17.987 ;
			RECT	103.175 17.923 103.207 17.987 ;
			RECT	150.122 17.939 150.154 17.971 ;
			RECT	150.575 17.939 150.607 17.971 ;
			RECT	151.13 17.923 151.194 17.987 ;
			RECT	152.244 17.939 152.276 17.971 ;
			RECT	153.552 17.923 153.616 17.987 ;
			RECT	153.805 17.923 153.837 17.987 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 15.98 201.665 16.09 ;
			LAYER	J3 ;
			RECT	0.756 16.003 0.788 16.067 ;
			RECT	1.645 16.003 1.709 16.067 ;
			RECT	2.323 16.003 2.387 16.067 ;
			RECT	3.438 16.003 3.47 16.067 ;
			RECT	3.585 16.003 3.617 16.067 ;
			RECT	4.195 16.003 4.227 16.067 ;
			RECT	4.704 16.019 4.768 16.051 ;
			RECT	4.944 16.003 5.008 16.067 ;
			RECT	52.124 16.019 52.156 16.051 ;
			RECT	52.577 16.019 52.609 16.051 ;
			RECT	53.132 16.003 53.196 16.067 ;
			RECT	54.246 16.019 54.278 16.051 ;
			RECT	55.554 16.003 55.618 16.067 ;
			RECT	55.807 16.003 55.839 16.067 ;
			RECT	102.995 16.003 103.027 16.067 ;
			RECT	103.175 16.003 103.207 16.067 ;
			RECT	150.122 16.019 150.154 16.051 ;
			RECT	150.575 16.019 150.607 16.051 ;
			RECT	151.13 16.003 151.194 16.067 ;
			RECT	152.244 16.019 152.276 16.051 ;
			RECT	153.552 16.003 153.616 16.067 ;
			RECT	153.805 16.003 153.837 16.067 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 14.06 201.665 14.17 ;
			LAYER	J3 ;
			RECT	0.756 14.083 0.788 14.147 ;
			RECT	1.645 14.083 1.709 14.147 ;
			RECT	2.323 14.083 2.387 14.147 ;
			RECT	3.438 14.083 3.47 14.147 ;
			RECT	3.585 14.083 3.617 14.147 ;
			RECT	4.195 14.083 4.227 14.147 ;
			RECT	4.704 14.099 4.768 14.131 ;
			RECT	4.944 14.083 5.008 14.147 ;
			RECT	52.124 14.099 52.156 14.131 ;
			RECT	52.577 14.099 52.609 14.131 ;
			RECT	53.132 14.083 53.196 14.147 ;
			RECT	54.246 14.099 54.278 14.131 ;
			RECT	55.554 14.083 55.618 14.147 ;
			RECT	55.807 14.083 55.839 14.147 ;
			RECT	102.995 14.083 103.027 14.147 ;
			RECT	103.175 14.083 103.207 14.147 ;
			RECT	150.122 14.099 150.154 14.131 ;
			RECT	150.575 14.099 150.607 14.131 ;
			RECT	151.13 14.083 151.194 14.147 ;
			RECT	152.244 14.099 152.276 14.131 ;
			RECT	153.552 14.083 153.616 14.147 ;
			RECT	153.805 14.083 153.837 14.147 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 12.14 201.665 12.25 ;
			LAYER	J3 ;
			RECT	0.756 12.163 0.788 12.227 ;
			RECT	1.645 12.163 1.709 12.227 ;
			RECT	2.323 12.163 2.387 12.227 ;
			RECT	3.438 12.163 3.47 12.227 ;
			RECT	3.585 12.163 3.617 12.227 ;
			RECT	4.195 12.163 4.227 12.227 ;
			RECT	4.704 12.179 4.768 12.211 ;
			RECT	4.944 12.163 5.008 12.227 ;
			RECT	52.124 12.179 52.156 12.211 ;
			RECT	52.577 12.179 52.609 12.211 ;
			RECT	53.132 12.163 53.196 12.227 ;
			RECT	54.246 12.179 54.278 12.211 ;
			RECT	55.554 12.163 55.618 12.227 ;
			RECT	55.807 12.163 55.839 12.227 ;
			RECT	102.995 12.163 103.027 12.227 ;
			RECT	103.175 12.163 103.207 12.227 ;
			RECT	150.122 12.179 150.154 12.211 ;
			RECT	150.575 12.179 150.607 12.211 ;
			RECT	151.13 12.163 151.194 12.227 ;
			RECT	152.244 12.179 152.276 12.211 ;
			RECT	153.552 12.163 153.616 12.227 ;
			RECT	153.805 12.163 153.837 12.227 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 10.22 201.665 10.33 ;
			LAYER	J3 ;
			RECT	0.756 10.243 0.788 10.307 ;
			RECT	1.645 10.243 1.709 10.307 ;
			RECT	2.323 10.243 2.387 10.307 ;
			RECT	3.438 10.243 3.47 10.307 ;
			RECT	3.585 10.243 3.617 10.307 ;
			RECT	4.195 10.243 4.227 10.307 ;
			RECT	4.704 10.259 4.768 10.291 ;
			RECT	4.944 10.243 5.008 10.307 ;
			RECT	52.124 10.259 52.156 10.291 ;
			RECT	52.577 10.259 52.609 10.291 ;
			RECT	53.132 10.243 53.196 10.307 ;
			RECT	54.246 10.259 54.278 10.291 ;
			RECT	55.554 10.243 55.618 10.307 ;
			RECT	55.807 10.243 55.839 10.307 ;
			RECT	102.995 10.243 103.027 10.307 ;
			RECT	103.175 10.243 103.207 10.307 ;
			RECT	150.122 10.259 150.154 10.291 ;
			RECT	150.575 10.259 150.607 10.291 ;
			RECT	151.13 10.243 151.194 10.307 ;
			RECT	152.244 10.259 152.276 10.291 ;
			RECT	153.552 10.243 153.616 10.307 ;
			RECT	153.805 10.243 153.837 10.307 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 8.3 201.665 8.41 ;
			LAYER	J3 ;
			RECT	0.756 8.323 0.788 8.387 ;
			RECT	1.645 8.323 1.709 8.387 ;
			RECT	2.323 8.323 2.387 8.387 ;
			RECT	3.438 8.323 3.47 8.387 ;
			RECT	3.585 8.323 3.617 8.387 ;
			RECT	4.195 8.323 4.227 8.387 ;
			RECT	4.704 8.339 4.768 8.371 ;
			RECT	4.944 8.323 5.008 8.387 ;
			RECT	52.124 8.339 52.156 8.371 ;
			RECT	52.577 8.339 52.609 8.371 ;
			RECT	53.132 8.323 53.196 8.387 ;
			RECT	54.246 8.339 54.278 8.371 ;
			RECT	55.554 8.323 55.618 8.387 ;
			RECT	55.807 8.323 55.839 8.387 ;
			RECT	102.995 8.323 103.027 8.387 ;
			RECT	103.175 8.323 103.207 8.387 ;
			RECT	150.122 8.339 150.154 8.371 ;
			RECT	150.575 8.339 150.607 8.371 ;
			RECT	151.13 8.323 151.194 8.387 ;
			RECT	152.244 8.339 152.276 8.371 ;
			RECT	153.552 8.323 153.616 8.387 ;
			RECT	153.805 8.323 153.837 8.387 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 6.38 201.665 6.49 ;
			LAYER	J3 ;
			RECT	0.756 6.403 0.788 6.467 ;
			RECT	1.645 6.403 1.709 6.467 ;
			RECT	2.323 6.403 2.387 6.467 ;
			RECT	3.438 6.403 3.47 6.467 ;
			RECT	3.585 6.403 3.617 6.467 ;
			RECT	4.195 6.403 4.227 6.467 ;
			RECT	4.704 6.419 4.768 6.451 ;
			RECT	4.944 6.403 5.008 6.467 ;
			RECT	52.124 6.419 52.156 6.451 ;
			RECT	52.577 6.419 52.609 6.451 ;
			RECT	53.132 6.403 53.196 6.467 ;
			RECT	54.246 6.419 54.278 6.451 ;
			RECT	55.554 6.403 55.618 6.467 ;
			RECT	55.807 6.403 55.839 6.467 ;
			RECT	102.995 6.403 103.027 6.467 ;
			RECT	103.175 6.403 103.207 6.467 ;
			RECT	150.122 6.419 150.154 6.451 ;
			RECT	150.575 6.419 150.607 6.451 ;
			RECT	151.13 6.403 151.194 6.467 ;
			RECT	152.244 6.419 152.276 6.451 ;
			RECT	153.552 6.403 153.616 6.467 ;
			RECT	153.805 6.403 153.837 6.467 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 4.46 201.665 4.57 ;
			LAYER	J3 ;
			RECT	0.756 4.483 0.788 4.547 ;
			RECT	1.645 4.483 1.709 4.547 ;
			RECT	2.323 4.483 2.387 4.547 ;
			RECT	3.438 4.483 3.47 4.547 ;
			RECT	3.585 4.483 3.617 4.547 ;
			RECT	4.195 4.483 4.227 4.547 ;
			RECT	4.704 4.499 4.768 4.531 ;
			RECT	4.944 4.483 5.008 4.547 ;
			RECT	52.124 4.499 52.156 4.531 ;
			RECT	52.577 4.499 52.609 4.531 ;
			RECT	53.132 4.483 53.196 4.547 ;
			RECT	54.246 4.499 54.278 4.531 ;
			RECT	55.554 4.483 55.618 4.547 ;
			RECT	55.807 4.483 55.839 4.547 ;
			RECT	102.995 4.483 103.027 4.547 ;
			RECT	103.175 4.483 103.207 4.547 ;
			RECT	150.122 4.499 150.154 4.531 ;
			RECT	150.575 4.499 150.607 4.531 ;
			RECT	151.13 4.483 151.194 4.547 ;
			RECT	152.244 4.499 152.276 4.531 ;
			RECT	153.552 4.483 153.616 4.547 ;
			RECT	153.805 4.483 153.837 4.547 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 73.766 201.665 73.876 ;
			LAYER	J3 ;
			RECT	0.756 73.789 0.788 73.853 ;
			RECT	1.645 73.789 1.709 73.853 ;
			RECT	2.323 73.789 2.387 73.853 ;
			RECT	3.438 73.789 3.47 73.853 ;
			RECT	3.585 73.789 3.617 73.853 ;
			RECT	4.195 73.789 4.227 73.853 ;
			RECT	4.704 73.805 4.768 73.837 ;
			RECT	4.944 73.789 5.008 73.853 ;
			RECT	52.124 73.805 52.156 73.837 ;
			RECT	52.577 73.805 52.609 73.837 ;
			RECT	53.132 73.789 53.196 73.853 ;
			RECT	54.246 73.805 54.278 73.837 ;
			RECT	55.554 73.789 55.618 73.853 ;
			RECT	55.807 73.789 55.839 73.853 ;
			RECT	102.995 73.789 103.027 73.853 ;
			RECT	103.175 73.789 103.207 73.853 ;
			RECT	150.122 73.805 150.154 73.837 ;
			RECT	150.575 73.805 150.607 73.837 ;
			RECT	151.13 73.789 151.194 73.853 ;
			RECT	152.244 73.805 152.276 73.837 ;
			RECT	153.552 73.789 153.616 73.853 ;
			RECT	153.805 73.789 153.837 73.853 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 2.54 201.665 2.65 ;
			LAYER	J3 ;
			RECT	0.756 2.563 0.788 2.627 ;
			RECT	1.645 2.563 1.709 2.627 ;
			RECT	2.323 2.563 2.387 2.627 ;
			RECT	3.438 2.563 3.47 2.627 ;
			RECT	3.585 2.563 3.617 2.627 ;
			RECT	4.195 2.563 4.227 2.627 ;
			RECT	4.704 2.579 4.768 2.611 ;
			RECT	4.944 2.563 5.008 2.627 ;
			RECT	52.124 2.579 52.156 2.611 ;
			RECT	52.577 2.579 52.609 2.611 ;
			RECT	53.132 2.563 53.196 2.627 ;
			RECT	54.246 2.579 54.278 2.611 ;
			RECT	55.554 2.563 55.618 2.627 ;
			RECT	55.807 2.563 55.839 2.627 ;
			RECT	102.995 2.563 103.027 2.627 ;
			RECT	103.175 2.563 103.207 2.627 ;
			RECT	150.122 2.579 150.154 2.611 ;
			RECT	150.575 2.579 150.607 2.611 ;
			RECT	151.13 2.563 151.194 2.627 ;
			RECT	152.244 2.579 152.276 2.611 ;
			RECT	153.552 2.563 153.616 2.627 ;
			RECT	153.805 2.563 153.837 2.627 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 71.846 201.665 71.956 ;
			LAYER	J3 ;
			RECT	0.756 71.869 0.788 71.933 ;
			RECT	1.645 71.869 1.709 71.933 ;
			RECT	2.323 71.869 2.387 71.933 ;
			RECT	3.438 71.869 3.47 71.933 ;
			RECT	3.585 71.869 3.617 71.933 ;
			RECT	4.195 71.869 4.227 71.933 ;
			RECT	4.704 71.885 4.768 71.917 ;
			RECT	4.944 71.869 5.008 71.933 ;
			RECT	52.124 71.885 52.156 71.917 ;
			RECT	52.577 71.885 52.609 71.917 ;
			RECT	53.132 71.869 53.196 71.933 ;
			RECT	54.246 71.885 54.278 71.917 ;
			RECT	55.554 71.869 55.618 71.933 ;
			RECT	55.807 71.869 55.839 71.933 ;
			RECT	102.995 71.869 103.027 71.933 ;
			RECT	103.175 71.869 103.207 71.933 ;
			RECT	150.122 71.885 150.154 71.917 ;
			RECT	150.575 71.885 150.607 71.917 ;
			RECT	151.13 71.869 151.194 71.933 ;
			RECT	152.244 71.885 152.276 71.917 ;
			RECT	153.552 71.869 153.616 71.933 ;
			RECT	153.805 71.869 153.837 71.933 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 69.926 201.665 70.036 ;
			LAYER	J3 ;
			RECT	0.756 69.949 0.788 70.013 ;
			RECT	1.645 69.949 1.709 70.013 ;
			RECT	2.323 69.949 2.387 70.013 ;
			RECT	3.438 69.949 3.47 70.013 ;
			RECT	3.585 69.949 3.617 70.013 ;
			RECT	4.195 69.949 4.227 70.013 ;
			RECT	4.704 69.965 4.768 69.997 ;
			RECT	4.944 69.949 5.008 70.013 ;
			RECT	52.124 69.965 52.156 69.997 ;
			RECT	52.577 69.965 52.609 69.997 ;
			RECT	53.132 69.949 53.196 70.013 ;
			RECT	54.246 69.965 54.278 69.997 ;
			RECT	55.554 69.949 55.618 70.013 ;
			RECT	55.807 69.949 55.839 70.013 ;
			RECT	102.995 69.949 103.027 70.013 ;
			RECT	103.175 69.949 103.207 70.013 ;
			RECT	150.122 69.965 150.154 69.997 ;
			RECT	150.575 69.965 150.607 69.997 ;
			RECT	151.13 69.949 151.194 70.013 ;
			RECT	152.244 69.965 152.276 69.997 ;
			RECT	153.552 69.949 153.616 70.013 ;
			RECT	153.805 69.949 153.837 70.013 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 68.006 201.665 68.116 ;
			LAYER	J3 ;
			RECT	0.756 68.029 0.788 68.093 ;
			RECT	1.645 68.029 1.709 68.093 ;
			RECT	2.323 68.029 2.387 68.093 ;
			RECT	3.438 68.029 3.47 68.093 ;
			RECT	3.585 68.029 3.617 68.093 ;
			RECT	4.195 68.029 4.227 68.093 ;
			RECT	4.704 68.045 4.768 68.077 ;
			RECT	4.944 68.029 5.008 68.093 ;
			RECT	52.124 68.045 52.156 68.077 ;
			RECT	52.577 68.045 52.609 68.077 ;
			RECT	53.132 68.029 53.196 68.093 ;
			RECT	54.246 68.045 54.278 68.077 ;
			RECT	55.554 68.029 55.618 68.093 ;
			RECT	55.807 68.029 55.839 68.093 ;
			RECT	102.995 68.029 103.027 68.093 ;
			RECT	103.175 68.029 103.207 68.093 ;
			RECT	150.122 68.045 150.154 68.077 ;
			RECT	150.575 68.045 150.607 68.077 ;
			RECT	151.13 68.029 151.194 68.093 ;
			RECT	152.244 68.045 152.276 68.077 ;
			RECT	153.552 68.029 153.616 68.093 ;
			RECT	153.805 68.029 153.837 68.093 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 66.086 201.665 66.196 ;
			LAYER	J3 ;
			RECT	0.756 66.109 0.788 66.173 ;
			RECT	1.645 66.109 1.709 66.173 ;
			RECT	2.323 66.109 2.387 66.173 ;
			RECT	3.438 66.109 3.47 66.173 ;
			RECT	3.585 66.109 3.617 66.173 ;
			RECT	4.195 66.109 4.227 66.173 ;
			RECT	4.704 66.125 4.768 66.157 ;
			RECT	4.944 66.109 5.008 66.173 ;
			RECT	52.124 66.125 52.156 66.157 ;
			RECT	52.577 66.125 52.609 66.157 ;
			RECT	53.132 66.109 53.196 66.173 ;
			RECT	54.246 66.125 54.278 66.157 ;
			RECT	55.554 66.109 55.618 66.173 ;
			RECT	55.807 66.109 55.839 66.173 ;
			RECT	102.995 66.109 103.027 66.173 ;
			RECT	103.175 66.109 103.207 66.173 ;
			RECT	150.122 66.125 150.154 66.157 ;
			RECT	150.575 66.125 150.607 66.157 ;
			RECT	151.13 66.109 151.194 66.173 ;
			RECT	152.244 66.125 152.276 66.157 ;
			RECT	153.552 66.109 153.616 66.173 ;
			RECT	153.805 66.109 153.837 66.173 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 64.166 201.665 64.276 ;
			LAYER	J3 ;
			RECT	0.756 64.189 0.788 64.253 ;
			RECT	1.645 64.189 1.709 64.253 ;
			RECT	2.323 64.189 2.387 64.253 ;
			RECT	3.438 64.189 3.47 64.253 ;
			RECT	3.585 64.189 3.617 64.253 ;
			RECT	4.195 64.189 4.227 64.253 ;
			RECT	4.704 64.205 4.768 64.237 ;
			RECT	4.944 64.189 5.008 64.253 ;
			RECT	52.124 64.205 52.156 64.237 ;
			RECT	52.577 64.205 52.609 64.237 ;
			RECT	53.132 64.189 53.196 64.253 ;
			RECT	54.246 64.205 54.278 64.237 ;
			RECT	55.554 64.189 55.618 64.253 ;
			RECT	55.807 64.189 55.839 64.253 ;
			RECT	102.995 64.189 103.027 64.253 ;
			RECT	103.175 64.189 103.207 64.253 ;
			RECT	150.122 64.205 150.154 64.237 ;
			RECT	150.575 64.205 150.607 64.237 ;
			RECT	151.13 64.189 151.194 64.253 ;
			RECT	152.244 64.205 152.276 64.237 ;
			RECT	153.552 64.189 153.616 64.253 ;
			RECT	153.805 64.189 153.837 64.253 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 62.246 201.665 62.356 ;
			LAYER	J3 ;
			RECT	0.756 62.269 0.788 62.333 ;
			RECT	1.645 62.269 1.709 62.333 ;
			RECT	2.323 62.269 2.387 62.333 ;
			RECT	3.438 62.269 3.47 62.333 ;
			RECT	3.585 62.269 3.617 62.333 ;
			RECT	4.195 62.269 4.227 62.333 ;
			RECT	4.704 62.285 4.768 62.317 ;
			RECT	4.944 62.269 5.008 62.333 ;
			RECT	52.124 62.285 52.156 62.317 ;
			RECT	52.577 62.285 52.609 62.317 ;
			RECT	53.132 62.269 53.196 62.333 ;
			RECT	54.246 62.285 54.278 62.317 ;
			RECT	55.554 62.269 55.618 62.333 ;
			RECT	55.807 62.269 55.839 62.333 ;
			RECT	102.995 62.269 103.027 62.333 ;
			RECT	103.175 62.269 103.207 62.333 ;
			RECT	150.122 62.285 150.154 62.317 ;
			RECT	150.575 62.285 150.607 62.317 ;
			RECT	151.13 62.269 151.194 62.333 ;
			RECT	152.244 62.285 152.276 62.317 ;
			RECT	153.552 62.269 153.616 62.333 ;
			RECT	153.805 62.269 153.837 62.333 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 60.326 201.665 60.436 ;
			LAYER	J3 ;
			RECT	0.756 60.349 0.788 60.413 ;
			RECT	1.645 60.349 1.709 60.413 ;
			RECT	2.323 60.349 2.387 60.413 ;
			RECT	3.438 60.349 3.47 60.413 ;
			RECT	3.585 60.349 3.617 60.413 ;
			RECT	4.195 60.349 4.227 60.413 ;
			RECT	4.704 60.365 4.768 60.397 ;
			RECT	4.944 60.349 5.008 60.413 ;
			RECT	52.124 60.365 52.156 60.397 ;
			RECT	52.577 60.365 52.609 60.397 ;
			RECT	53.132 60.349 53.196 60.413 ;
			RECT	54.246 60.365 54.278 60.397 ;
			RECT	55.554 60.349 55.618 60.413 ;
			RECT	55.807 60.349 55.839 60.413 ;
			RECT	102.995 60.349 103.027 60.413 ;
			RECT	103.175 60.349 103.207 60.413 ;
			RECT	150.122 60.365 150.154 60.397 ;
			RECT	150.575 60.365 150.607 60.397 ;
			RECT	151.13 60.349 151.194 60.413 ;
			RECT	152.244 60.365 152.276 60.397 ;
			RECT	153.552 60.349 153.616 60.413 ;
			RECT	153.805 60.349 153.837 60.413 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 58.406 201.665 58.516 ;
			LAYER	J3 ;
			RECT	0.756 58.429 0.788 58.493 ;
			RECT	1.645 58.429 1.709 58.493 ;
			RECT	2.323 58.429 2.387 58.493 ;
			RECT	3.438 58.429 3.47 58.493 ;
			RECT	3.585 58.429 3.617 58.493 ;
			RECT	4.195 58.429 4.227 58.493 ;
			RECT	4.704 58.445 4.768 58.477 ;
			RECT	4.944 58.429 5.008 58.493 ;
			RECT	52.124 58.445 52.156 58.477 ;
			RECT	52.577 58.445 52.609 58.477 ;
			RECT	53.132 58.429 53.196 58.493 ;
			RECT	54.246 58.445 54.278 58.477 ;
			RECT	55.554 58.429 55.618 58.493 ;
			RECT	55.807 58.429 55.839 58.493 ;
			RECT	102.995 58.429 103.027 58.493 ;
			RECT	103.175 58.429 103.207 58.493 ;
			RECT	150.122 58.445 150.154 58.477 ;
			RECT	150.575 58.445 150.607 58.477 ;
			RECT	151.13 58.429 151.194 58.493 ;
			RECT	152.244 58.445 152.276 58.477 ;
			RECT	153.552 58.429 153.616 58.493 ;
			RECT	153.805 58.429 153.837 58.493 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 56.486 201.665 56.596 ;
			LAYER	J3 ;
			RECT	0.756 56.509 0.788 56.573 ;
			RECT	1.645 56.509 1.709 56.573 ;
			RECT	2.323 56.509 2.387 56.573 ;
			RECT	3.438 56.509 3.47 56.573 ;
			RECT	3.585 56.509 3.617 56.573 ;
			RECT	4.195 56.509 4.227 56.573 ;
			RECT	4.704 56.525 4.768 56.557 ;
			RECT	4.944 56.509 5.008 56.573 ;
			RECT	52.124 56.525 52.156 56.557 ;
			RECT	52.577 56.525 52.609 56.557 ;
			RECT	53.132 56.509 53.196 56.573 ;
			RECT	54.246 56.525 54.278 56.557 ;
			RECT	55.554 56.509 55.618 56.573 ;
			RECT	55.807 56.509 55.839 56.573 ;
			RECT	102.995 56.509 103.027 56.573 ;
			RECT	103.175 56.509 103.207 56.573 ;
			RECT	150.122 56.525 150.154 56.557 ;
			RECT	150.575 56.525 150.607 56.557 ;
			RECT	151.13 56.509 151.194 56.573 ;
			RECT	152.244 56.525 152.276 56.557 ;
			RECT	153.552 56.509 153.616 56.573 ;
			RECT	153.805 56.509 153.837 56.573 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 54.566 201.665 54.676 ;
			LAYER	J3 ;
			RECT	0.756 54.589 0.788 54.653 ;
			RECT	1.645 54.589 1.709 54.653 ;
			RECT	2.323 54.589 2.387 54.653 ;
			RECT	3.438 54.589 3.47 54.653 ;
			RECT	3.585 54.589 3.617 54.653 ;
			RECT	4.195 54.589 4.227 54.653 ;
			RECT	4.704 54.605 4.768 54.637 ;
			RECT	4.944 54.589 5.008 54.653 ;
			RECT	52.124 54.605 52.156 54.637 ;
			RECT	52.577 54.605 52.609 54.637 ;
			RECT	53.132 54.589 53.196 54.653 ;
			RECT	54.246 54.605 54.278 54.637 ;
			RECT	55.554 54.589 55.618 54.653 ;
			RECT	55.807 54.589 55.839 54.653 ;
			RECT	102.995 54.589 103.027 54.653 ;
			RECT	103.175 54.589 103.207 54.653 ;
			RECT	150.122 54.605 150.154 54.637 ;
			RECT	150.575 54.605 150.607 54.637 ;
			RECT	151.13 54.589 151.194 54.653 ;
			RECT	152.244 54.605 152.276 54.637 ;
			RECT	153.552 54.589 153.616 54.653 ;
			RECT	153.805 54.589 153.837 54.653 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 52.646 201.665 52.756 ;
			LAYER	J3 ;
			RECT	0.756 52.669 0.788 52.733 ;
			RECT	1.645 52.669 1.709 52.733 ;
			RECT	2.323 52.669 2.387 52.733 ;
			RECT	3.438 52.669 3.47 52.733 ;
			RECT	3.585 52.669 3.617 52.733 ;
			RECT	4.195 52.669 4.227 52.733 ;
			RECT	4.704 52.685 4.768 52.717 ;
			RECT	4.944 52.669 5.008 52.733 ;
			RECT	52.124 52.685 52.156 52.717 ;
			RECT	52.577 52.685 52.609 52.717 ;
			RECT	53.132 52.669 53.196 52.733 ;
			RECT	54.246 52.685 54.278 52.717 ;
			RECT	55.554 52.669 55.618 52.733 ;
			RECT	55.807 52.669 55.839 52.733 ;
			RECT	102.995 52.669 103.027 52.733 ;
			RECT	103.175 52.669 103.207 52.733 ;
			RECT	150.122 52.685 150.154 52.717 ;
			RECT	150.575 52.685 150.607 52.717 ;
			RECT	151.13 52.669 151.194 52.733 ;
			RECT	152.244 52.685 152.276 52.717 ;
			RECT	153.552 52.669 153.616 52.733 ;
			RECT	153.805 52.669 153.837 52.733 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 50.726 201.665 50.836 ;
			LAYER	J3 ;
			RECT	0.756 50.749 0.788 50.813 ;
			RECT	1.645 50.749 1.709 50.813 ;
			RECT	2.323 50.749 2.387 50.813 ;
			RECT	3.438 50.749 3.47 50.813 ;
			RECT	3.585 50.749 3.617 50.813 ;
			RECT	4.195 50.749 4.227 50.813 ;
			RECT	4.704 50.765 4.768 50.797 ;
			RECT	4.944 50.749 5.008 50.813 ;
			RECT	52.124 50.765 52.156 50.797 ;
			RECT	52.577 50.765 52.609 50.797 ;
			RECT	53.132 50.749 53.196 50.813 ;
			RECT	54.246 50.765 54.278 50.797 ;
			RECT	55.554 50.749 55.618 50.813 ;
			RECT	55.807 50.749 55.839 50.813 ;
			RECT	102.995 50.749 103.027 50.813 ;
			RECT	103.175 50.749 103.207 50.813 ;
			RECT	150.122 50.765 150.154 50.797 ;
			RECT	150.575 50.765 150.607 50.797 ;
			RECT	151.13 50.749 151.194 50.813 ;
			RECT	152.244 50.765 152.276 50.797 ;
			RECT	153.552 50.749 153.616 50.813 ;
			RECT	153.805 50.749 153.837 50.813 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 81.458 201.665 81.578 ;
			LAYER	J3 ;
			RECT	0.755 81.486 0.787 81.55 ;
			RECT	1.645 81.486 1.709 81.55 ;
			RECT	2.323 81.486 2.387 81.55 ;
			RECT	3.438 81.486 3.47 81.55 ;
			RECT	3.585 81.486 3.617 81.55 ;
			RECT	4.195 81.486 4.227 81.55 ;
			RECT	4.944 81.486 5.008 81.55 ;
			RECT	5.927 81.486 5.959 81.55 ;
			RECT	6.179 81.486 6.211 81.55 ;
			RECT	6.347 81.486 6.379 81.55 ;
			RECT	6.515 81.486 6.547 81.55 ;
			RECT	6.683 81.486 6.715 81.55 ;
			RECT	6.851 81.486 6.883 81.55 ;
			RECT	7.019 81.486 7.051 81.55 ;
			RECT	7.187 81.486 7.219 81.55 ;
			RECT	7.355 81.486 7.387 81.55 ;
			RECT	7.523 81.486 7.555 81.55 ;
			RECT	7.691 81.486 7.723 81.55 ;
			RECT	7.859 81.486 7.891 81.55 ;
			RECT	8.027 81.486 8.059 81.55 ;
			RECT	8.195 81.486 8.227 81.55 ;
			RECT	8.363 81.486 8.395 81.55 ;
			RECT	8.531 81.486 8.563 81.55 ;
			RECT	8.699 81.486 8.731 81.55 ;
			RECT	8.867 81.486 8.899 81.55 ;
			RECT	9.035 81.486 9.067 81.55 ;
			RECT	9.203 81.486 9.235 81.55 ;
			RECT	9.371 81.486 9.403 81.55 ;
			RECT	9.539 81.486 9.571 81.55 ;
			RECT	9.707 81.486 9.739 81.55 ;
			RECT	9.875 81.486 9.907 81.55 ;
			RECT	10.043 81.486 10.075 81.55 ;
			RECT	10.211 81.486 10.243 81.55 ;
			RECT	10.379 81.486 10.411 81.55 ;
			RECT	10.547 81.486 10.579 81.55 ;
			RECT	10.715 81.486 10.747 81.55 ;
			RECT	10.883 81.486 10.915 81.55 ;
			RECT	11.051 81.486 11.083 81.55 ;
			RECT	11.219 81.486 11.251 81.55 ;
			RECT	11.387 81.486 11.419 81.55 ;
			RECT	11.555 81.486 11.587 81.55 ;
			RECT	11.723 81.486 11.755 81.55 ;
			RECT	11.891 81.486 11.923 81.55 ;
			RECT	12.059 81.486 12.091 81.55 ;
			RECT	12.227 81.486 12.259 81.55 ;
			RECT	12.395 81.486 12.427 81.55 ;
			RECT	12.563 81.486 12.595 81.55 ;
			RECT	12.731 81.486 12.763 81.55 ;
			RECT	12.899 81.486 12.931 81.55 ;
			RECT	13.067 81.486 13.099 81.55 ;
			RECT	13.235 81.486 13.267 81.55 ;
			RECT	13.403 81.486 13.435 81.55 ;
			RECT	13.571 81.486 13.603 81.55 ;
			RECT	13.739 81.486 13.771 81.55 ;
			RECT	13.907 81.486 13.939 81.55 ;
			RECT	14.075 81.486 14.107 81.55 ;
			RECT	14.243 81.486 14.275 81.55 ;
			RECT	14.411 81.486 14.443 81.55 ;
			RECT	14.579 81.486 14.611 81.55 ;
			RECT	14.747 81.486 14.779 81.55 ;
			RECT	14.915 81.486 14.947 81.55 ;
			RECT	15.083 81.486 15.115 81.55 ;
			RECT	15.251 81.486 15.283 81.55 ;
			RECT	15.419 81.486 15.451 81.55 ;
			RECT	15.587 81.486 15.619 81.55 ;
			RECT	15.755 81.486 15.787 81.55 ;
			RECT	15.923 81.486 15.955 81.55 ;
			RECT	16.091 81.486 16.123 81.55 ;
			RECT	16.259 81.486 16.291 81.55 ;
			RECT	16.427 81.486 16.459 81.55 ;
			RECT	16.595 81.486 16.627 81.55 ;
			RECT	16.763 81.486 16.795 81.55 ;
			RECT	16.931 81.486 16.963 81.55 ;
			RECT	17.099 81.486 17.131 81.55 ;
			RECT	17.267 81.486 17.299 81.55 ;
			RECT	17.435 81.486 17.467 81.55 ;
			RECT	17.603 81.486 17.635 81.55 ;
			RECT	17.771 81.486 17.803 81.55 ;
			RECT	17.939 81.486 17.971 81.55 ;
			RECT	18.107 81.486 18.139 81.55 ;
			RECT	18.275 81.486 18.307 81.55 ;
			RECT	18.443 81.486 18.475 81.55 ;
			RECT	18.611 81.486 18.643 81.55 ;
			RECT	18.779 81.486 18.811 81.55 ;
			RECT	18.947 81.486 18.979 81.55 ;
			RECT	19.115 81.486 19.147 81.55 ;
			RECT	19.283 81.486 19.315 81.55 ;
			RECT	19.451 81.486 19.483 81.55 ;
			RECT	19.619 81.486 19.651 81.55 ;
			RECT	19.787 81.486 19.819 81.55 ;
			RECT	19.955 81.486 19.987 81.55 ;
			RECT	20.123 81.486 20.155 81.55 ;
			RECT	20.291 81.486 20.323 81.55 ;
			RECT	20.459 81.486 20.491 81.55 ;
			RECT	20.627 81.486 20.659 81.55 ;
			RECT	20.795 81.486 20.827 81.55 ;
			RECT	20.963 81.486 20.995 81.55 ;
			RECT	21.131 81.486 21.163 81.55 ;
			RECT	21.299 81.486 21.331 81.55 ;
			RECT	21.467 81.486 21.499 81.55 ;
			RECT	21.635 81.486 21.667 81.55 ;
			RECT	21.803 81.486 21.835 81.55 ;
			RECT	21.971 81.486 22.003 81.55 ;
			RECT	22.139 81.486 22.171 81.55 ;
			RECT	22.307 81.486 22.339 81.55 ;
			RECT	22.475 81.486 22.507 81.55 ;
			RECT	22.643 81.486 22.675 81.55 ;
			RECT	22.811 81.486 22.843 81.55 ;
			RECT	22.979 81.486 23.011 81.55 ;
			RECT	23.147 81.486 23.179 81.55 ;
			RECT	23.315 81.486 23.347 81.55 ;
			RECT	23.483 81.486 23.515 81.55 ;
			RECT	23.651 81.486 23.683 81.55 ;
			RECT	23.819 81.486 23.851 81.55 ;
			RECT	23.987 81.486 24.019 81.55 ;
			RECT	24.155 81.486 24.187 81.55 ;
			RECT	24.323 81.486 24.355 81.55 ;
			RECT	24.491 81.486 24.523 81.55 ;
			RECT	24.659 81.486 24.691 81.55 ;
			RECT	24.827 81.486 24.859 81.55 ;
			RECT	24.995 81.486 25.027 81.55 ;
			RECT	25.163 81.486 25.195 81.55 ;
			RECT	25.331 81.486 25.363 81.55 ;
			RECT	25.499 81.486 25.531 81.55 ;
			RECT	25.667 81.486 25.699 81.55 ;
			RECT	25.835 81.486 25.867 81.55 ;
			RECT	26.003 81.486 26.035 81.55 ;
			RECT	26.171 81.486 26.203 81.55 ;
			RECT	26.339 81.486 26.371 81.55 ;
			RECT	26.507 81.486 26.539 81.55 ;
			RECT	26.675 81.486 26.707 81.55 ;
			RECT	26.843 81.486 26.875 81.55 ;
			RECT	27.011 81.486 27.043 81.55 ;
			RECT	27.179 81.486 27.211 81.55 ;
			RECT	27.347 81.486 27.379 81.55 ;
			RECT	27.515 81.486 27.547 81.55 ;
			RECT	27.683 81.486 27.715 81.55 ;
			RECT	27.851 81.486 27.883 81.55 ;
			RECT	28.019 81.486 28.051 81.55 ;
			RECT	28.187 81.486 28.219 81.55 ;
			RECT	28.355 81.486 28.387 81.55 ;
			RECT	28.523 81.486 28.555 81.55 ;
			RECT	28.691 81.486 28.723 81.55 ;
			RECT	28.859 81.486 28.891 81.55 ;
			RECT	29.027 81.486 29.059 81.55 ;
			RECT	29.195 81.486 29.227 81.55 ;
			RECT	29.363 81.486 29.395 81.55 ;
			RECT	29.531 81.486 29.563 81.55 ;
			RECT	29.699 81.486 29.731 81.55 ;
			RECT	29.867 81.486 29.899 81.55 ;
			RECT	30.035 81.486 30.067 81.55 ;
			RECT	30.203 81.486 30.235 81.55 ;
			RECT	30.371 81.486 30.403 81.55 ;
			RECT	30.539 81.486 30.571 81.55 ;
			RECT	30.707 81.486 30.739 81.55 ;
			RECT	30.875 81.486 30.907 81.55 ;
			RECT	31.043 81.486 31.075 81.55 ;
			RECT	31.211 81.486 31.243 81.55 ;
			RECT	31.379 81.486 31.411 81.55 ;
			RECT	31.547 81.486 31.579 81.55 ;
			RECT	31.715 81.486 31.747 81.55 ;
			RECT	31.883 81.486 31.915 81.55 ;
			RECT	32.051 81.486 32.083 81.55 ;
			RECT	32.219 81.486 32.251 81.55 ;
			RECT	32.387 81.486 32.419 81.55 ;
			RECT	32.555 81.486 32.587 81.55 ;
			RECT	32.723 81.486 32.755 81.55 ;
			RECT	32.891 81.486 32.923 81.55 ;
			RECT	33.059 81.486 33.091 81.55 ;
			RECT	33.227 81.486 33.259 81.55 ;
			RECT	33.395 81.486 33.427 81.55 ;
			RECT	33.563 81.486 33.595 81.55 ;
			RECT	33.731 81.486 33.763 81.55 ;
			RECT	33.899 81.486 33.931 81.55 ;
			RECT	34.067 81.486 34.099 81.55 ;
			RECT	34.235 81.486 34.267 81.55 ;
			RECT	34.403 81.486 34.435 81.55 ;
			RECT	34.571 81.486 34.603 81.55 ;
			RECT	34.739 81.486 34.771 81.55 ;
			RECT	34.907 81.486 34.939 81.55 ;
			RECT	35.075 81.486 35.107 81.55 ;
			RECT	35.243 81.486 35.275 81.55 ;
			RECT	35.411 81.486 35.443 81.55 ;
			RECT	35.579 81.486 35.611 81.55 ;
			RECT	35.747 81.486 35.779 81.55 ;
			RECT	35.915 81.486 35.947 81.55 ;
			RECT	36.083 81.486 36.115 81.55 ;
			RECT	36.251 81.486 36.283 81.55 ;
			RECT	36.419 81.486 36.451 81.55 ;
			RECT	36.587 81.486 36.619 81.55 ;
			RECT	36.755 81.486 36.787 81.55 ;
			RECT	36.923 81.486 36.955 81.55 ;
			RECT	37.091 81.486 37.123 81.55 ;
			RECT	37.259 81.486 37.291 81.55 ;
			RECT	37.427 81.486 37.459 81.55 ;
			RECT	37.595 81.486 37.627 81.55 ;
			RECT	37.763 81.486 37.795 81.55 ;
			RECT	37.931 81.486 37.963 81.55 ;
			RECT	38.099 81.486 38.131 81.55 ;
			RECT	38.267 81.486 38.299 81.55 ;
			RECT	38.435 81.486 38.467 81.55 ;
			RECT	38.603 81.486 38.635 81.55 ;
			RECT	38.771 81.486 38.803 81.55 ;
			RECT	38.939 81.486 38.971 81.55 ;
			RECT	39.107 81.486 39.139 81.55 ;
			RECT	39.275 81.486 39.307 81.55 ;
			RECT	39.443 81.486 39.475 81.55 ;
			RECT	39.611 81.486 39.643 81.55 ;
			RECT	39.779 81.486 39.811 81.55 ;
			RECT	39.947 81.486 39.979 81.55 ;
			RECT	40.115 81.486 40.147 81.55 ;
			RECT	40.283 81.486 40.315 81.55 ;
			RECT	40.451 81.486 40.483 81.55 ;
			RECT	40.619 81.486 40.651 81.55 ;
			RECT	40.787 81.486 40.819 81.55 ;
			RECT	40.955 81.486 40.987 81.55 ;
			RECT	41.123 81.486 41.155 81.55 ;
			RECT	41.291 81.486 41.323 81.55 ;
			RECT	41.459 81.486 41.491 81.55 ;
			RECT	41.627 81.486 41.659 81.55 ;
			RECT	41.795 81.486 41.827 81.55 ;
			RECT	41.963 81.486 41.995 81.55 ;
			RECT	42.131 81.486 42.163 81.55 ;
			RECT	42.299 81.486 42.331 81.55 ;
			RECT	42.467 81.486 42.499 81.55 ;
			RECT	42.635 81.486 42.667 81.55 ;
			RECT	42.803 81.486 42.835 81.55 ;
			RECT	42.971 81.486 43.003 81.55 ;
			RECT	43.139 81.486 43.171 81.55 ;
			RECT	43.307 81.486 43.339 81.55 ;
			RECT	43.475 81.486 43.507 81.55 ;
			RECT	43.643 81.486 43.675 81.55 ;
			RECT	43.811 81.486 43.843 81.55 ;
			RECT	43.979 81.486 44.011 81.55 ;
			RECT	44.147 81.486 44.179 81.55 ;
			RECT	44.315 81.486 44.347 81.55 ;
			RECT	44.483 81.486 44.515 81.55 ;
			RECT	44.651 81.486 44.683 81.55 ;
			RECT	44.819 81.486 44.851 81.55 ;
			RECT	44.987 81.486 45.019 81.55 ;
			RECT	45.155 81.486 45.187 81.55 ;
			RECT	45.323 81.486 45.355 81.55 ;
			RECT	45.491 81.486 45.523 81.55 ;
			RECT	45.659 81.486 45.691 81.55 ;
			RECT	45.827 81.486 45.859 81.55 ;
			RECT	45.995 81.486 46.027 81.55 ;
			RECT	46.163 81.486 46.195 81.55 ;
			RECT	46.331 81.486 46.363 81.55 ;
			RECT	46.499 81.486 46.531 81.55 ;
			RECT	46.667 81.486 46.699 81.55 ;
			RECT	46.835 81.486 46.867 81.55 ;
			RECT	47.003 81.486 47.035 81.55 ;
			RECT	47.171 81.486 47.203 81.55 ;
			RECT	47.339 81.486 47.371 81.55 ;
			RECT	47.507 81.486 47.539 81.55 ;
			RECT	47.675 81.486 47.707 81.55 ;
			RECT	47.843 81.486 47.875 81.55 ;
			RECT	48.011 81.486 48.043 81.55 ;
			RECT	48.179 81.486 48.211 81.55 ;
			RECT	48.347 81.486 48.379 81.55 ;
			RECT	48.515 81.486 48.547 81.55 ;
			RECT	48.683 81.486 48.715 81.55 ;
			RECT	48.851 81.486 48.883 81.55 ;
			RECT	49.019 81.486 49.051 81.55 ;
			RECT	49.187 81.486 49.219 81.55 ;
			RECT	49.541 81.486 49.605 81.55 ;
			RECT	52.124 81.486 52.156 81.55 ;
			RECT	52.578 81.486 52.61 81.55 ;
			RECT	53.132 81.486 53.196 81.55 ;
			RECT	53.911 81.486 53.943 81.55 ;
			RECT	54.251 81.486 54.283 81.55 ;
			RECT	55.562 81.486 55.626 81.55 ;
			RECT	58.599 81.486 58.663 81.55 ;
			RECT	58.985 81.486 59.017 81.55 ;
			RECT	59.153 81.486 59.185 81.55 ;
			RECT	59.321 81.486 59.353 81.55 ;
			RECT	59.489 81.486 59.521 81.55 ;
			RECT	59.657 81.486 59.689 81.55 ;
			RECT	59.825 81.486 59.857 81.55 ;
			RECT	59.993 81.486 60.025 81.55 ;
			RECT	60.161 81.486 60.193 81.55 ;
			RECT	60.329 81.486 60.361 81.55 ;
			RECT	60.497 81.486 60.529 81.55 ;
			RECT	60.665 81.486 60.697 81.55 ;
			RECT	60.833 81.486 60.865 81.55 ;
			RECT	61.001 81.486 61.033 81.55 ;
			RECT	61.169 81.486 61.201 81.55 ;
			RECT	61.337 81.486 61.369 81.55 ;
			RECT	61.505 81.486 61.537 81.55 ;
			RECT	61.673 81.486 61.705 81.55 ;
			RECT	61.841 81.486 61.873 81.55 ;
			RECT	62.009 81.486 62.041 81.55 ;
			RECT	62.177 81.486 62.209 81.55 ;
			RECT	62.345 81.486 62.377 81.55 ;
			RECT	62.513 81.486 62.545 81.55 ;
			RECT	62.681 81.486 62.713 81.55 ;
			RECT	62.849 81.486 62.881 81.55 ;
			RECT	63.017 81.486 63.049 81.55 ;
			RECT	63.185 81.486 63.217 81.55 ;
			RECT	63.353 81.486 63.385 81.55 ;
			RECT	63.521 81.486 63.553 81.55 ;
			RECT	63.689 81.486 63.721 81.55 ;
			RECT	63.857 81.486 63.889 81.55 ;
			RECT	64.025 81.486 64.057 81.55 ;
			RECT	64.193 81.486 64.225 81.55 ;
			RECT	64.361 81.486 64.393 81.55 ;
			RECT	64.529 81.486 64.561 81.55 ;
			RECT	64.697 81.486 64.729 81.55 ;
			RECT	64.865 81.486 64.897 81.55 ;
			RECT	65.033 81.486 65.065 81.55 ;
			RECT	65.201 81.486 65.233 81.55 ;
			RECT	65.369 81.486 65.401 81.55 ;
			RECT	65.537 81.486 65.569 81.55 ;
			RECT	65.705 81.486 65.737 81.55 ;
			RECT	65.873 81.486 65.905 81.55 ;
			RECT	66.041 81.486 66.073 81.55 ;
			RECT	66.209 81.486 66.241 81.55 ;
			RECT	66.377 81.486 66.409 81.55 ;
			RECT	66.545 81.486 66.577 81.55 ;
			RECT	66.713 81.486 66.745 81.55 ;
			RECT	66.881 81.486 66.913 81.55 ;
			RECT	67.049 81.486 67.081 81.55 ;
			RECT	67.217 81.486 67.249 81.55 ;
			RECT	67.385 81.486 67.417 81.55 ;
			RECT	67.553 81.486 67.585 81.55 ;
			RECT	67.721 81.486 67.753 81.55 ;
			RECT	67.889 81.486 67.921 81.55 ;
			RECT	68.057 81.486 68.089 81.55 ;
			RECT	68.225 81.486 68.257 81.55 ;
			RECT	68.393 81.486 68.425 81.55 ;
			RECT	68.561 81.486 68.593 81.55 ;
			RECT	68.729 81.486 68.761 81.55 ;
			RECT	68.897 81.486 68.929 81.55 ;
			RECT	69.065 81.486 69.097 81.55 ;
			RECT	69.233 81.486 69.265 81.55 ;
			RECT	69.401 81.486 69.433 81.55 ;
			RECT	69.569 81.486 69.601 81.55 ;
			RECT	69.737 81.486 69.769 81.55 ;
			RECT	69.905 81.486 69.937 81.55 ;
			RECT	70.073 81.486 70.105 81.55 ;
			RECT	70.241 81.486 70.273 81.55 ;
			RECT	70.409 81.486 70.441 81.55 ;
			RECT	70.577 81.486 70.609 81.55 ;
			RECT	70.745 81.486 70.777 81.55 ;
			RECT	70.913 81.486 70.945 81.55 ;
			RECT	71.081 81.486 71.113 81.55 ;
			RECT	71.249 81.486 71.281 81.55 ;
			RECT	71.417 81.486 71.449 81.55 ;
			RECT	71.585 81.486 71.617 81.55 ;
			RECT	71.753 81.486 71.785 81.55 ;
			RECT	71.921 81.486 71.953 81.55 ;
			RECT	72.089 81.486 72.121 81.55 ;
			RECT	72.257 81.486 72.289 81.55 ;
			RECT	72.425 81.486 72.457 81.55 ;
			RECT	72.593 81.486 72.625 81.55 ;
			RECT	72.761 81.486 72.793 81.55 ;
			RECT	72.929 81.486 72.961 81.55 ;
			RECT	73.097 81.486 73.129 81.55 ;
			RECT	73.265 81.486 73.297 81.55 ;
			RECT	73.433 81.486 73.465 81.55 ;
			RECT	73.601 81.486 73.633 81.55 ;
			RECT	73.769 81.486 73.801 81.55 ;
			RECT	73.937 81.486 73.969 81.55 ;
			RECT	74.105 81.486 74.137 81.55 ;
			RECT	74.273 81.486 74.305 81.55 ;
			RECT	74.441 81.486 74.473 81.55 ;
			RECT	74.609 81.486 74.641 81.55 ;
			RECT	74.777 81.486 74.809 81.55 ;
			RECT	74.945 81.486 74.977 81.55 ;
			RECT	75.113 81.486 75.145 81.55 ;
			RECT	75.281 81.486 75.313 81.55 ;
			RECT	75.449 81.486 75.481 81.55 ;
			RECT	75.617 81.486 75.649 81.55 ;
			RECT	75.785 81.486 75.817 81.55 ;
			RECT	75.953 81.486 75.985 81.55 ;
			RECT	76.121 81.486 76.153 81.55 ;
			RECT	76.289 81.486 76.321 81.55 ;
			RECT	76.457 81.486 76.489 81.55 ;
			RECT	76.625 81.486 76.657 81.55 ;
			RECT	76.793 81.486 76.825 81.55 ;
			RECT	76.961 81.486 76.993 81.55 ;
			RECT	77.129 81.486 77.161 81.55 ;
			RECT	77.297 81.486 77.329 81.55 ;
			RECT	77.465 81.486 77.497 81.55 ;
			RECT	77.633 81.486 77.665 81.55 ;
			RECT	77.801 81.486 77.833 81.55 ;
			RECT	77.969 81.486 78.001 81.55 ;
			RECT	78.137 81.486 78.169 81.55 ;
			RECT	78.305 81.486 78.337 81.55 ;
			RECT	78.473 81.486 78.505 81.55 ;
			RECT	78.641 81.486 78.673 81.55 ;
			RECT	78.809 81.486 78.841 81.55 ;
			RECT	78.977 81.486 79.009 81.55 ;
			RECT	79.145 81.486 79.177 81.55 ;
			RECT	79.313 81.486 79.345 81.55 ;
			RECT	79.481 81.486 79.513 81.55 ;
			RECT	79.649 81.486 79.681 81.55 ;
			RECT	79.817 81.486 79.849 81.55 ;
			RECT	79.985 81.486 80.017 81.55 ;
			RECT	80.153 81.486 80.185 81.55 ;
			RECT	80.321 81.486 80.353 81.55 ;
			RECT	80.489 81.486 80.521 81.55 ;
			RECT	80.657 81.486 80.689 81.55 ;
			RECT	80.825 81.486 80.857 81.55 ;
			RECT	80.993 81.486 81.025 81.55 ;
			RECT	81.161 81.486 81.193 81.55 ;
			RECT	81.329 81.486 81.361 81.55 ;
			RECT	81.497 81.486 81.529 81.55 ;
			RECT	81.665 81.486 81.697 81.55 ;
			RECT	81.833 81.486 81.865 81.55 ;
			RECT	82.001 81.486 82.033 81.55 ;
			RECT	82.169 81.486 82.201 81.55 ;
			RECT	82.337 81.486 82.369 81.55 ;
			RECT	82.505 81.486 82.537 81.55 ;
			RECT	82.673 81.486 82.705 81.55 ;
			RECT	82.841 81.486 82.873 81.55 ;
			RECT	83.009 81.486 83.041 81.55 ;
			RECT	83.177 81.486 83.209 81.55 ;
			RECT	83.345 81.486 83.377 81.55 ;
			RECT	83.513 81.486 83.545 81.55 ;
			RECT	83.681 81.486 83.713 81.55 ;
			RECT	83.849 81.486 83.881 81.55 ;
			RECT	84.017 81.486 84.049 81.55 ;
			RECT	84.185 81.486 84.217 81.55 ;
			RECT	84.353 81.486 84.385 81.55 ;
			RECT	84.521 81.486 84.553 81.55 ;
			RECT	84.689 81.486 84.721 81.55 ;
			RECT	84.857 81.486 84.889 81.55 ;
			RECT	85.025 81.486 85.057 81.55 ;
			RECT	85.193 81.486 85.225 81.55 ;
			RECT	85.361 81.486 85.393 81.55 ;
			RECT	85.529 81.486 85.561 81.55 ;
			RECT	85.697 81.486 85.729 81.55 ;
			RECT	85.865 81.486 85.897 81.55 ;
			RECT	86.033 81.486 86.065 81.55 ;
			RECT	86.201 81.486 86.233 81.55 ;
			RECT	86.369 81.486 86.401 81.55 ;
			RECT	86.537 81.486 86.569 81.55 ;
			RECT	86.705 81.486 86.737 81.55 ;
			RECT	86.873 81.486 86.905 81.55 ;
			RECT	87.041 81.486 87.073 81.55 ;
			RECT	87.209 81.486 87.241 81.55 ;
			RECT	87.377 81.486 87.409 81.55 ;
			RECT	87.545 81.486 87.577 81.55 ;
			RECT	87.713 81.486 87.745 81.55 ;
			RECT	87.881 81.486 87.913 81.55 ;
			RECT	88.049 81.486 88.081 81.55 ;
			RECT	88.217 81.486 88.249 81.55 ;
			RECT	88.385 81.486 88.417 81.55 ;
			RECT	88.553 81.486 88.585 81.55 ;
			RECT	88.721 81.486 88.753 81.55 ;
			RECT	88.889 81.486 88.921 81.55 ;
			RECT	89.057 81.486 89.089 81.55 ;
			RECT	89.225 81.486 89.257 81.55 ;
			RECT	89.393 81.486 89.425 81.55 ;
			RECT	89.561 81.486 89.593 81.55 ;
			RECT	89.729 81.486 89.761 81.55 ;
			RECT	89.897 81.486 89.929 81.55 ;
			RECT	90.065 81.486 90.097 81.55 ;
			RECT	90.233 81.486 90.265 81.55 ;
			RECT	90.401 81.486 90.433 81.55 ;
			RECT	90.569 81.486 90.601 81.55 ;
			RECT	90.737 81.486 90.769 81.55 ;
			RECT	90.905 81.486 90.937 81.55 ;
			RECT	91.073 81.486 91.105 81.55 ;
			RECT	91.241 81.486 91.273 81.55 ;
			RECT	91.409 81.486 91.441 81.55 ;
			RECT	91.577 81.486 91.609 81.55 ;
			RECT	91.745 81.486 91.777 81.55 ;
			RECT	91.913 81.486 91.945 81.55 ;
			RECT	92.081 81.486 92.113 81.55 ;
			RECT	92.249 81.486 92.281 81.55 ;
			RECT	92.417 81.486 92.449 81.55 ;
			RECT	92.585 81.486 92.617 81.55 ;
			RECT	92.753 81.486 92.785 81.55 ;
			RECT	92.921 81.486 92.953 81.55 ;
			RECT	93.089 81.486 93.121 81.55 ;
			RECT	93.257 81.486 93.289 81.55 ;
			RECT	93.425 81.486 93.457 81.55 ;
			RECT	93.593 81.486 93.625 81.55 ;
			RECT	93.761 81.486 93.793 81.55 ;
			RECT	93.929 81.486 93.961 81.55 ;
			RECT	94.097 81.486 94.129 81.55 ;
			RECT	94.265 81.486 94.297 81.55 ;
			RECT	94.433 81.486 94.465 81.55 ;
			RECT	94.601 81.486 94.633 81.55 ;
			RECT	94.769 81.486 94.801 81.55 ;
			RECT	94.937 81.486 94.969 81.55 ;
			RECT	95.105 81.486 95.137 81.55 ;
			RECT	95.273 81.486 95.305 81.55 ;
			RECT	95.441 81.486 95.473 81.55 ;
			RECT	95.609 81.486 95.641 81.55 ;
			RECT	95.777 81.486 95.809 81.55 ;
			RECT	95.945 81.486 95.977 81.55 ;
			RECT	96.113 81.486 96.145 81.55 ;
			RECT	96.281 81.486 96.313 81.55 ;
			RECT	96.449 81.486 96.481 81.55 ;
			RECT	96.617 81.486 96.649 81.55 ;
			RECT	96.785 81.486 96.817 81.55 ;
			RECT	96.953 81.486 96.985 81.55 ;
			RECT	97.121 81.486 97.153 81.55 ;
			RECT	97.289 81.486 97.321 81.55 ;
			RECT	97.457 81.486 97.489 81.55 ;
			RECT	97.625 81.486 97.657 81.55 ;
			RECT	97.793 81.486 97.825 81.55 ;
			RECT	97.961 81.486 97.993 81.55 ;
			RECT	98.129 81.486 98.161 81.55 ;
			RECT	98.297 81.486 98.329 81.55 ;
			RECT	98.465 81.486 98.497 81.55 ;
			RECT	98.633 81.486 98.665 81.55 ;
			RECT	98.801 81.486 98.833 81.55 ;
			RECT	98.969 81.486 99.001 81.55 ;
			RECT	99.137 81.486 99.169 81.55 ;
			RECT	99.305 81.486 99.337 81.55 ;
			RECT	99.473 81.486 99.505 81.55 ;
			RECT	99.641 81.486 99.673 81.55 ;
			RECT	99.809 81.486 99.841 81.55 ;
			RECT	99.977 81.486 100.009 81.55 ;
			RECT	100.145 81.486 100.177 81.55 ;
			RECT	100.313 81.486 100.345 81.55 ;
			RECT	100.481 81.486 100.513 81.55 ;
			RECT	100.649 81.486 100.681 81.55 ;
			RECT	100.817 81.486 100.849 81.55 ;
			RECT	100.985 81.486 101.017 81.55 ;
			RECT	101.153 81.486 101.185 81.55 ;
			RECT	101.321 81.486 101.353 81.55 ;
			RECT	101.489 81.486 101.521 81.55 ;
			RECT	101.657 81.486 101.689 81.55 ;
			RECT	101.825 81.486 101.857 81.55 ;
			RECT	101.993 81.486 102.025 81.55 ;
			RECT	102.245 81.486 102.277 81.55 ;
			RECT	103.085 81.486 103.117 81.55 ;
			RECT	103.925 81.486 103.957 81.55 ;
			RECT	104.177 81.486 104.209 81.55 ;
			RECT	104.345 81.486 104.377 81.55 ;
			RECT	104.513 81.486 104.545 81.55 ;
			RECT	104.681 81.486 104.713 81.55 ;
			RECT	104.849 81.486 104.881 81.55 ;
			RECT	105.017 81.486 105.049 81.55 ;
			RECT	105.185 81.486 105.217 81.55 ;
			RECT	105.353 81.486 105.385 81.55 ;
			RECT	105.521 81.486 105.553 81.55 ;
			RECT	105.689 81.486 105.721 81.55 ;
			RECT	105.857 81.486 105.889 81.55 ;
			RECT	106.025 81.486 106.057 81.55 ;
			RECT	106.193 81.486 106.225 81.55 ;
			RECT	106.361 81.486 106.393 81.55 ;
			RECT	106.529 81.486 106.561 81.55 ;
			RECT	106.697 81.486 106.729 81.55 ;
			RECT	106.865 81.486 106.897 81.55 ;
			RECT	107.033 81.486 107.065 81.55 ;
			RECT	107.201 81.486 107.233 81.55 ;
			RECT	107.369 81.486 107.401 81.55 ;
			RECT	107.537 81.486 107.569 81.55 ;
			RECT	107.705 81.486 107.737 81.55 ;
			RECT	107.873 81.486 107.905 81.55 ;
			RECT	108.041 81.486 108.073 81.55 ;
			RECT	108.209 81.486 108.241 81.55 ;
			RECT	108.377 81.486 108.409 81.55 ;
			RECT	108.545 81.486 108.577 81.55 ;
			RECT	108.713 81.486 108.745 81.55 ;
			RECT	108.881 81.486 108.913 81.55 ;
			RECT	109.049 81.486 109.081 81.55 ;
			RECT	109.217 81.486 109.249 81.55 ;
			RECT	109.385 81.486 109.417 81.55 ;
			RECT	109.553 81.486 109.585 81.55 ;
			RECT	109.721 81.486 109.753 81.55 ;
			RECT	109.889 81.486 109.921 81.55 ;
			RECT	110.057 81.486 110.089 81.55 ;
			RECT	110.225 81.486 110.257 81.55 ;
			RECT	110.393 81.486 110.425 81.55 ;
			RECT	110.561 81.486 110.593 81.55 ;
			RECT	110.729 81.486 110.761 81.55 ;
			RECT	110.897 81.486 110.929 81.55 ;
			RECT	111.065 81.486 111.097 81.55 ;
			RECT	111.233 81.486 111.265 81.55 ;
			RECT	111.401 81.486 111.433 81.55 ;
			RECT	111.569 81.486 111.601 81.55 ;
			RECT	111.737 81.486 111.769 81.55 ;
			RECT	111.905 81.486 111.937 81.55 ;
			RECT	112.073 81.486 112.105 81.55 ;
			RECT	112.241 81.486 112.273 81.55 ;
			RECT	112.409 81.486 112.441 81.55 ;
			RECT	112.577 81.486 112.609 81.55 ;
			RECT	112.745 81.486 112.777 81.55 ;
			RECT	112.913 81.486 112.945 81.55 ;
			RECT	113.081 81.486 113.113 81.55 ;
			RECT	113.249 81.486 113.281 81.55 ;
			RECT	113.417 81.486 113.449 81.55 ;
			RECT	113.585 81.486 113.617 81.55 ;
			RECT	113.753 81.486 113.785 81.55 ;
			RECT	113.921 81.486 113.953 81.55 ;
			RECT	114.089 81.486 114.121 81.55 ;
			RECT	114.257 81.486 114.289 81.55 ;
			RECT	114.425 81.486 114.457 81.55 ;
			RECT	114.593 81.486 114.625 81.55 ;
			RECT	114.761 81.486 114.793 81.55 ;
			RECT	114.929 81.486 114.961 81.55 ;
			RECT	115.097 81.486 115.129 81.55 ;
			RECT	115.265 81.486 115.297 81.55 ;
			RECT	115.433 81.486 115.465 81.55 ;
			RECT	115.601 81.486 115.633 81.55 ;
			RECT	115.769 81.486 115.801 81.55 ;
			RECT	115.937 81.486 115.969 81.55 ;
			RECT	116.105 81.486 116.137 81.55 ;
			RECT	116.273 81.486 116.305 81.55 ;
			RECT	116.441 81.486 116.473 81.55 ;
			RECT	116.609 81.486 116.641 81.55 ;
			RECT	116.777 81.486 116.809 81.55 ;
			RECT	116.945 81.486 116.977 81.55 ;
			RECT	117.113 81.486 117.145 81.55 ;
			RECT	117.281 81.486 117.313 81.55 ;
			RECT	117.449 81.486 117.481 81.55 ;
			RECT	117.617 81.486 117.649 81.55 ;
			RECT	117.785 81.486 117.817 81.55 ;
			RECT	117.953 81.486 117.985 81.55 ;
			RECT	118.121 81.486 118.153 81.55 ;
			RECT	118.289 81.486 118.321 81.55 ;
			RECT	118.457 81.486 118.489 81.55 ;
			RECT	118.625 81.486 118.657 81.55 ;
			RECT	118.793 81.486 118.825 81.55 ;
			RECT	118.961 81.486 118.993 81.55 ;
			RECT	119.129 81.486 119.161 81.55 ;
			RECT	119.297 81.486 119.329 81.55 ;
			RECT	119.465 81.486 119.497 81.55 ;
			RECT	119.633 81.486 119.665 81.55 ;
			RECT	119.801 81.486 119.833 81.55 ;
			RECT	119.969 81.486 120.001 81.55 ;
			RECT	120.137 81.486 120.169 81.55 ;
			RECT	120.305 81.486 120.337 81.55 ;
			RECT	120.473 81.486 120.505 81.55 ;
			RECT	120.641 81.486 120.673 81.55 ;
			RECT	120.809 81.486 120.841 81.55 ;
			RECT	120.977 81.486 121.009 81.55 ;
			RECT	121.145 81.486 121.177 81.55 ;
			RECT	121.313 81.486 121.345 81.55 ;
			RECT	121.481 81.486 121.513 81.55 ;
			RECT	121.649 81.486 121.681 81.55 ;
			RECT	121.817 81.486 121.849 81.55 ;
			RECT	121.985 81.486 122.017 81.55 ;
			RECT	122.153 81.486 122.185 81.55 ;
			RECT	122.321 81.486 122.353 81.55 ;
			RECT	122.489 81.486 122.521 81.55 ;
			RECT	122.657 81.486 122.689 81.55 ;
			RECT	122.825 81.486 122.857 81.55 ;
			RECT	122.993 81.486 123.025 81.55 ;
			RECT	123.161 81.486 123.193 81.55 ;
			RECT	123.329 81.486 123.361 81.55 ;
			RECT	123.497 81.486 123.529 81.55 ;
			RECT	123.665 81.486 123.697 81.55 ;
			RECT	123.833 81.486 123.865 81.55 ;
			RECT	124.001 81.486 124.033 81.55 ;
			RECT	124.169 81.486 124.201 81.55 ;
			RECT	124.337 81.486 124.369 81.55 ;
			RECT	124.505 81.486 124.537 81.55 ;
			RECT	124.673 81.486 124.705 81.55 ;
			RECT	124.841 81.486 124.873 81.55 ;
			RECT	125.009 81.486 125.041 81.55 ;
			RECT	125.177 81.486 125.209 81.55 ;
			RECT	125.345 81.486 125.377 81.55 ;
			RECT	125.513 81.486 125.545 81.55 ;
			RECT	125.681 81.486 125.713 81.55 ;
			RECT	125.849 81.486 125.881 81.55 ;
			RECT	126.017 81.486 126.049 81.55 ;
			RECT	126.185 81.486 126.217 81.55 ;
			RECT	126.353 81.486 126.385 81.55 ;
			RECT	126.521 81.486 126.553 81.55 ;
			RECT	126.689 81.486 126.721 81.55 ;
			RECT	126.857 81.486 126.889 81.55 ;
			RECT	127.025 81.486 127.057 81.55 ;
			RECT	127.193 81.486 127.225 81.55 ;
			RECT	127.361 81.486 127.393 81.55 ;
			RECT	127.529 81.486 127.561 81.55 ;
			RECT	127.697 81.486 127.729 81.55 ;
			RECT	127.865 81.486 127.897 81.55 ;
			RECT	128.033 81.486 128.065 81.55 ;
			RECT	128.201 81.486 128.233 81.55 ;
			RECT	128.369 81.486 128.401 81.55 ;
			RECT	128.537 81.486 128.569 81.55 ;
			RECT	128.705 81.486 128.737 81.55 ;
			RECT	128.873 81.486 128.905 81.55 ;
			RECT	129.041 81.486 129.073 81.55 ;
			RECT	129.209 81.486 129.241 81.55 ;
			RECT	129.377 81.486 129.409 81.55 ;
			RECT	129.545 81.486 129.577 81.55 ;
			RECT	129.713 81.486 129.745 81.55 ;
			RECT	129.881 81.486 129.913 81.55 ;
			RECT	130.049 81.486 130.081 81.55 ;
			RECT	130.217 81.486 130.249 81.55 ;
			RECT	130.385 81.486 130.417 81.55 ;
			RECT	130.553 81.486 130.585 81.55 ;
			RECT	130.721 81.486 130.753 81.55 ;
			RECT	130.889 81.486 130.921 81.55 ;
			RECT	131.057 81.486 131.089 81.55 ;
			RECT	131.225 81.486 131.257 81.55 ;
			RECT	131.393 81.486 131.425 81.55 ;
			RECT	131.561 81.486 131.593 81.55 ;
			RECT	131.729 81.486 131.761 81.55 ;
			RECT	131.897 81.486 131.929 81.55 ;
			RECT	132.065 81.486 132.097 81.55 ;
			RECT	132.233 81.486 132.265 81.55 ;
			RECT	132.401 81.486 132.433 81.55 ;
			RECT	132.569 81.486 132.601 81.55 ;
			RECT	132.737 81.486 132.769 81.55 ;
			RECT	132.905 81.486 132.937 81.55 ;
			RECT	133.073 81.486 133.105 81.55 ;
			RECT	133.241 81.486 133.273 81.55 ;
			RECT	133.409 81.486 133.441 81.55 ;
			RECT	133.577 81.486 133.609 81.55 ;
			RECT	133.745 81.486 133.777 81.55 ;
			RECT	133.913 81.486 133.945 81.55 ;
			RECT	134.081 81.486 134.113 81.55 ;
			RECT	134.249 81.486 134.281 81.55 ;
			RECT	134.417 81.486 134.449 81.55 ;
			RECT	134.585 81.486 134.617 81.55 ;
			RECT	134.753 81.486 134.785 81.55 ;
			RECT	134.921 81.486 134.953 81.55 ;
			RECT	135.089 81.486 135.121 81.55 ;
			RECT	135.257 81.486 135.289 81.55 ;
			RECT	135.425 81.486 135.457 81.55 ;
			RECT	135.593 81.486 135.625 81.55 ;
			RECT	135.761 81.486 135.793 81.55 ;
			RECT	135.929 81.486 135.961 81.55 ;
			RECT	136.097 81.486 136.129 81.55 ;
			RECT	136.265 81.486 136.297 81.55 ;
			RECT	136.433 81.486 136.465 81.55 ;
			RECT	136.601 81.486 136.633 81.55 ;
			RECT	136.769 81.486 136.801 81.55 ;
			RECT	136.937 81.486 136.969 81.55 ;
			RECT	137.105 81.486 137.137 81.55 ;
			RECT	137.273 81.486 137.305 81.55 ;
			RECT	137.441 81.486 137.473 81.55 ;
			RECT	137.609 81.486 137.641 81.55 ;
			RECT	137.777 81.486 137.809 81.55 ;
			RECT	137.945 81.486 137.977 81.55 ;
			RECT	138.113 81.486 138.145 81.55 ;
			RECT	138.281 81.486 138.313 81.55 ;
			RECT	138.449 81.486 138.481 81.55 ;
			RECT	138.617 81.486 138.649 81.55 ;
			RECT	138.785 81.486 138.817 81.55 ;
			RECT	138.953 81.486 138.985 81.55 ;
			RECT	139.121 81.486 139.153 81.55 ;
			RECT	139.289 81.486 139.321 81.55 ;
			RECT	139.457 81.486 139.489 81.55 ;
			RECT	139.625 81.486 139.657 81.55 ;
			RECT	139.793 81.486 139.825 81.55 ;
			RECT	139.961 81.486 139.993 81.55 ;
			RECT	140.129 81.486 140.161 81.55 ;
			RECT	140.297 81.486 140.329 81.55 ;
			RECT	140.465 81.486 140.497 81.55 ;
			RECT	140.633 81.486 140.665 81.55 ;
			RECT	140.801 81.486 140.833 81.55 ;
			RECT	140.969 81.486 141.001 81.55 ;
			RECT	141.137 81.486 141.169 81.55 ;
			RECT	141.305 81.486 141.337 81.55 ;
			RECT	141.473 81.486 141.505 81.55 ;
			RECT	141.641 81.486 141.673 81.55 ;
			RECT	141.809 81.486 141.841 81.55 ;
			RECT	141.977 81.486 142.009 81.55 ;
			RECT	142.145 81.486 142.177 81.55 ;
			RECT	142.313 81.486 142.345 81.55 ;
			RECT	142.481 81.486 142.513 81.55 ;
			RECT	142.649 81.486 142.681 81.55 ;
			RECT	142.817 81.486 142.849 81.55 ;
			RECT	142.985 81.486 143.017 81.55 ;
			RECT	143.153 81.486 143.185 81.55 ;
			RECT	143.321 81.486 143.353 81.55 ;
			RECT	143.489 81.486 143.521 81.55 ;
			RECT	143.657 81.486 143.689 81.55 ;
			RECT	143.825 81.486 143.857 81.55 ;
			RECT	143.993 81.486 144.025 81.55 ;
			RECT	144.161 81.486 144.193 81.55 ;
			RECT	144.329 81.486 144.361 81.55 ;
			RECT	144.497 81.486 144.529 81.55 ;
			RECT	144.665 81.486 144.697 81.55 ;
			RECT	144.833 81.486 144.865 81.55 ;
			RECT	145.001 81.486 145.033 81.55 ;
			RECT	145.169 81.486 145.201 81.55 ;
			RECT	145.337 81.486 145.369 81.55 ;
			RECT	145.505 81.486 145.537 81.55 ;
			RECT	145.673 81.486 145.705 81.55 ;
			RECT	145.841 81.486 145.873 81.55 ;
			RECT	146.009 81.486 146.041 81.55 ;
			RECT	146.177 81.486 146.209 81.55 ;
			RECT	146.345 81.486 146.377 81.55 ;
			RECT	146.513 81.486 146.545 81.55 ;
			RECT	146.681 81.486 146.713 81.55 ;
			RECT	146.849 81.486 146.881 81.55 ;
			RECT	147.017 81.486 147.049 81.55 ;
			RECT	147.185 81.486 147.217 81.55 ;
			RECT	147.539 81.486 147.603 81.55 ;
			RECT	150.122 81.486 150.154 81.55 ;
			RECT	150.576 81.486 150.608 81.55 ;
			RECT	151.13 81.486 151.194 81.55 ;
			RECT	151.909 81.486 151.941 81.55 ;
			RECT	152.249 81.486 152.281 81.55 ;
			RECT	153.56 81.486 153.624 81.55 ;
			RECT	156.597 81.486 156.661 81.55 ;
			RECT	156.983 81.486 157.015 81.55 ;
			RECT	157.151 81.486 157.183 81.55 ;
			RECT	157.319 81.486 157.351 81.55 ;
			RECT	157.487 81.486 157.519 81.55 ;
			RECT	157.655 81.486 157.687 81.55 ;
			RECT	157.823 81.486 157.855 81.55 ;
			RECT	157.991 81.486 158.023 81.55 ;
			RECT	158.159 81.486 158.191 81.55 ;
			RECT	158.327 81.486 158.359 81.55 ;
			RECT	158.495 81.486 158.527 81.55 ;
			RECT	158.663 81.486 158.695 81.55 ;
			RECT	158.831 81.486 158.863 81.55 ;
			RECT	158.999 81.486 159.031 81.55 ;
			RECT	159.167 81.486 159.199 81.55 ;
			RECT	159.335 81.486 159.367 81.55 ;
			RECT	159.503 81.486 159.535 81.55 ;
			RECT	159.671 81.486 159.703 81.55 ;
			RECT	159.839 81.486 159.871 81.55 ;
			RECT	160.007 81.486 160.039 81.55 ;
			RECT	160.175 81.486 160.207 81.55 ;
			RECT	160.343 81.486 160.375 81.55 ;
			RECT	160.511 81.486 160.543 81.55 ;
			RECT	160.679 81.486 160.711 81.55 ;
			RECT	160.847 81.486 160.879 81.55 ;
			RECT	161.015 81.486 161.047 81.55 ;
			RECT	161.183 81.486 161.215 81.55 ;
			RECT	161.351 81.486 161.383 81.55 ;
			RECT	161.519 81.486 161.551 81.55 ;
			RECT	161.687 81.486 161.719 81.55 ;
			RECT	161.855 81.486 161.887 81.55 ;
			RECT	162.023 81.486 162.055 81.55 ;
			RECT	162.191 81.486 162.223 81.55 ;
			RECT	162.359 81.486 162.391 81.55 ;
			RECT	162.527 81.486 162.559 81.55 ;
			RECT	162.695 81.486 162.727 81.55 ;
			RECT	162.863 81.486 162.895 81.55 ;
			RECT	163.031 81.486 163.063 81.55 ;
			RECT	163.199 81.486 163.231 81.55 ;
			RECT	163.367 81.486 163.399 81.55 ;
			RECT	163.535 81.486 163.567 81.55 ;
			RECT	163.703 81.486 163.735 81.55 ;
			RECT	163.871 81.486 163.903 81.55 ;
			RECT	164.039 81.486 164.071 81.55 ;
			RECT	164.207 81.486 164.239 81.55 ;
			RECT	164.375 81.486 164.407 81.55 ;
			RECT	164.543 81.486 164.575 81.55 ;
			RECT	164.711 81.486 164.743 81.55 ;
			RECT	164.879 81.486 164.911 81.55 ;
			RECT	165.047 81.486 165.079 81.55 ;
			RECT	165.215 81.486 165.247 81.55 ;
			RECT	165.383 81.486 165.415 81.55 ;
			RECT	165.551 81.486 165.583 81.55 ;
			RECT	165.719 81.486 165.751 81.55 ;
			RECT	165.887 81.486 165.919 81.55 ;
			RECT	166.055 81.486 166.087 81.55 ;
			RECT	166.223 81.486 166.255 81.55 ;
			RECT	166.391 81.486 166.423 81.55 ;
			RECT	166.559 81.486 166.591 81.55 ;
			RECT	166.727 81.486 166.759 81.55 ;
			RECT	166.895 81.486 166.927 81.55 ;
			RECT	167.063 81.486 167.095 81.55 ;
			RECT	167.231 81.486 167.263 81.55 ;
			RECT	167.399 81.486 167.431 81.55 ;
			RECT	167.567 81.486 167.599 81.55 ;
			RECT	167.735 81.486 167.767 81.55 ;
			RECT	167.903 81.486 167.935 81.55 ;
			RECT	168.071 81.486 168.103 81.55 ;
			RECT	168.239 81.486 168.271 81.55 ;
			RECT	168.407 81.486 168.439 81.55 ;
			RECT	168.575 81.486 168.607 81.55 ;
			RECT	168.743 81.486 168.775 81.55 ;
			RECT	168.911 81.486 168.943 81.55 ;
			RECT	169.079 81.486 169.111 81.55 ;
			RECT	169.247 81.486 169.279 81.55 ;
			RECT	169.415 81.486 169.447 81.55 ;
			RECT	169.583 81.486 169.615 81.55 ;
			RECT	169.751 81.486 169.783 81.55 ;
			RECT	169.919 81.486 169.951 81.55 ;
			RECT	170.087 81.486 170.119 81.55 ;
			RECT	170.255 81.486 170.287 81.55 ;
			RECT	170.423 81.486 170.455 81.55 ;
			RECT	170.591 81.486 170.623 81.55 ;
			RECT	170.759 81.486 170.791 81.55 ;
			RECT	170.927 81.486 170.959 81.55 ;
			RECT	171.095 81.486 171.127 81.55 ;
			RECT	171.263 81.486 171.295 81.55 ;
			RECT	171.431 81.486 171.463 81.55 ;
			RECT	171.599 81.486 171.631 81.55 ;
			RECT	171.767 81.486 171.799 81.55 ;
			RECT	171.935 81.486 171.967 81.55 ;
			RECT	172.103 81.486 172.135 81.55 ;
			RECT	172.271 81.486 172.303 81.55 ;
			RECT	172.439 81.486 172.471 81.55 ;
			RECT	172.607 81.486 172.639 81.55 ;
			RECT	172.775 81.486 172.807 81.55 ;
			RECT	172.943 81.486 172.975 81.55 ;
			RECT	173.111 81.486 173.143 81.55 ;
			RECT	173.279 81.486 173.311 81.55 ;
			RECT	173.447 81.486 173.479 81.55 ;
			RECT	173.615 81.486 173.647 81.55 ;
			RECT	173.783 81.486 173.815 81.55 ;
			RECT	173.951 81.486 173.983 81.55 ;
			RECT	174.119 81.486 174.151 81.55 ;
			RECT	174.287 81.486 174.319 81.55 ;
			RECT	174.455 81.486 174.487 81.55 ;
			RECT	174.623 81.486 174.655 81.55 ;
			RECT	174.791 81.486 174.823 81.55 ;
			RECT	174.959 81.486 174.991 81.55 ;
			RECT	175.127 81.486 175.159 81.55 ;
			RECT	175.295 81.486 175.327 81.55 ;
			RECT	175.463 81.486 175.495 81.55 ;
			RECT	175.631 81.486 175.663 81.55 ;
			RECT	175.799 81.486 175.831 81.55 ;
			RECT	175.967 81.486 175.999 81.55 ;
			RECT	176.135 81.486 176.167 81.55 ;
			RECT	176.303 81.486 176.335 81.55 ;
			RECT	176.471 81.486 176.503 81.55 ;
			RECT	176.639 81.486 176.671 81.55 ;
			RECT	176.807 81.486 176.839 81.55 ;
			RECT	176.975 81.486 177.007 81.55 ;
			RECT	177.143 81.486 177.175 81.55 ;
			RECT	177.311 81.486 177.343 81.55 ;
			RECT	177.479 81.486 177.511 81.55 ;
			RECT	177.647 81.486 177.679 81.55 ;
			RECT	177.815 81.486 177.847 81.55 ;
			RECT	177.983 81.486 178.015 81.55 ;
			RECT	178.151 81.486 178.183 81.55 ;
			RECT	178.319 81.486 178.351 81.55 ;
			RECT	178.487 81.486 178.519 81.55 ;
			RECT	178.655 81.486 178.687 81.55 ;
			RECT	178.823 81.486 178.855 81.55 ;
			RECT	178.991 81.486 179.023 81.55 ;
			RECT	179.159 81.486 179.191 81.55 ;
			RECT	179.327 81.486 179.359 81.55 ;
			RECT	179.495 81.486 179.527 81.55 ;
			RECT	179.663 81.486 179.695 81.55 ;
			RECT	179.831 81.486 179.863 81.55 ;
			RECT	179.999 81.486 180.031 81.55 ;
			RECT	180.167 81.486 180.199 81.55 ;
			RECT	180.335 81.486 180.367 81.55 ;
			RECT	180.503 81.486 180.535 81.55 ;
			RECT	180.671 81.486 180.703 81.55 ;
			RECT	180.839 81.486 180.871 81.55 ;
			RECT	181.007 81.486 181.039 81.55 ;
			RECT	181.175 81.486 181.207 81.55 ;
			RECT	181.343 81.486 181.375 81.55 ;
			RECT	181.511 81.486 181.543 81.55 ;
			RECT	181.679 81.486 181.711 81.55 ;
			RECT	181.847 81.486 181.879 81.55 ;
			RECT	182.015 81.486 182.047 81.55 ;
			RECT	182.183 81.486 182.215 81.55 ;
			RECT	182.351 81.486 182.383 81.55 ;
			RECT	182.519 81.486 182.551 81.55 ;
			RECT	182.687 81.486 182.719 81.55 ;
			RECT	182.855 81.486 182.887 81.55 ;
			RECT	183.023 81.486 183.055 81.55 ;
			RECT	183.191 81.486 183.223 81.55 ;
			RECT	183.359 81.486 183.391 81.55 ;
			RECT	183.527 81.486 183.559 81.55 ;
			RECT	183.695 81.486 183.727 81.55 ;
			RECT	183.863 81.486 183.895 81.55 ;
			RECT	184.031 81.486 184.063 81.55 ;
			RECT	184.199 81.486 184.231 81.55 ;
			RECT	184.367 81.486 184.399 81.55 ;
			RECT	184.535 81.486 184.567 81.55 ;
			RECT	184.703 81.486 184.735 81.55 ;
			RECT	184.871 81.486 184.903 81.55 ;
			RECT	185.039 81.486 185.071 81.55 ;
			RECT	185.207 81.486 185.239 81.55 ;
			RECT	185.375 81.486 185.407 81.55 ;
			RECT	185.543 81.486 185.575 81.55 ;
			RECT	185.711 81.486 185.743 81.55 ;
			RECT	185.879 81.486 185.911 81.55 ;
			RECT	186.047 81.486 186.079 81.55 ;
			RECT	186.215 81.486 186.247 81.55 ;
			RECT	186.383 81.486 186.415 81.55 ;
			RECT	186.551 81.486 186.583 81.55 ;
			RECT	186.719 81.486 186.751 81.55 ;
			RECT	186.887 81.486 186.919 81.55 ;
			RECT	187.055 81.486 187.087 81.55 ;
			RECT	187.223 81.486 187.255 81.55 ;
			RECT	187.391 81.486 187.423 81.55 ;
			RECT	187.559 81.486 187.591 81.55 ;
			RECT	187.727 81.486 187.759 81.55 ;
			RECT	187.895 81.486 187.927 81.55 ;
			RECT	188.063 81.486 188.095 81.55 ;
			RECT	188.231 81.486 188.263 81.55 ;
			RECT	188.399 81.486 188.431 81.55 ;
			RECT	188.567 81.486 188.599 81.55 ;
			RECT	188.735 81.486 188.767 81.55 ;
			RECT	188.903 81.486 188.935 81.55 ;
			RECT	189.071 81.486 189.103 81.55 ;
			RECT	189.239 81.486 189.271 81.55 ;
			RECT	189.407 81.486 189.439 81.55 ;
			RECT	189.575 81.486 189.607 81.55 ;
			RECT	189.743 81.486 189.775 81.55 ;
			RECT	189.911 81.486 189.943 81.55 ;
			RECT	190.079 81.486 190.111 81.55 ;
			RECT	190.247 81.486 190.279 81.55 ;
			RECT	190.415 81.486 190.447 81.55 ;
			RECT	190.583 81.486 190.615 81.55 ;
			RECT	190.751 81.486 190.783 81.55 ;
			RECT	190.919 81.486 190.951 81.55 ;
			RECT	191.087 81.486 191.119 81.55 ;
			RECT	191.255 81.486 191.287 81.55 ;
			RECT	191.423 81.486 191.455 81.55 ;
			RECT	191.591 81.486 191.623 81.55 ;
			RECT	191.759 81.486 191.791 81.55 ;
			RECT	191.927 81.486 191.959 81.55 ;
			RECT	192.095 81.486 192.127 81.55 ;
			RECT	192.263 81.486 192.295 81.55 ;
			RECT	192.431 81.486 192.463 81.55 ;
			RECT	192.599 81.486 192.631 81.55 ;
			RECT	192.767 81.486 192.799 81.55 ;
			RECT	192.935 81.486 192.967 81.55 ;
			RECT	193.103 81.486 193.135 81.55 ;
			RECT	193.271 81.486 193.303 81.55 ;
			RECT	193.439 81.486 193.471 81.55 ;
			RECT	193.607 81.486 193.639 81.55 ;
			RECT	193.775 81.486 193.807 81.55 ;
			RECT	193.943 81.486 193.975 81.55 ;
			RECT	194.111 81.486 194.143 81.55 ;
			RECT	194.279 81.486 194.311 81.55 ;
			RECT	194.447 81.486 194.479 81.55 ;
			RECT	194.615 81.486 194.647 81.55 ;
			RECT	194.783 81.486 194.815 81.55 ;
			RECT	194.951 81.486 194.983 81.55 ;
			RECT	195.119 81.486 195.151 81.55 ;
			RECT	195.287 81.486 195.319 81.55 ;
			RECT	195.455 81.486 195.487 81.55 ;
			RECT	195.623 81.486 195.655 81.55 ;
			RECT	195.791 81.486 195.823 81.55 ;
			RECT	195.959 81.486 195.991 81.55 ;
			RECT	196.127 81.486 196.159 81.55 ;
			RECT	196.295 81.486 196.327 81.55 ;
			RECT	196.463 81.486 196.495 81.55 ;
			RECT	196.631 81.486 196.663 81.55 ;
			RECT	196.799 81.486 196.831 81.55 ;
			RECT	196.967 81.486 196.999 81.55 ;
			RECT	197.135 81.486 197.167 81.55 ;
			RECT	197.303 81.486 197.335 81.55 ;
			RECT	197.471 81.486 197.503 81.55 ;
			RECT	197.639 81.486 197.671 81.55 ;
			RECT	197.807 81.486 197.839 81.55 ;
			RECT	197.975 81.486 198.007 81.55 ;
			RECT	198.143 81.486 198.175 81.55 ;
			RECT	198.311 81.486 198.343 81.55 ;
			RECT	198.479 81.486 198.511 81.55 ;
			RECT	198.647 81.486 198.679 81.55 ;
			RECT	198.815 81.486 198.847 81.55 ;
			RECT	198.983 81.486 199.015 81.55 ;
			RECT	199.151 81.486 199.183 81.55 ;
			RECT	199.319 81.486 199.351 81.55 ;
			RECT	199.487 81.486 199.519 81.55 ;
			RECT	199.655 81.486 199.687 81.55 ;
			RECT	199.823 81.486 199.855 81.55 ;
			RECT	199.991 81.486 200.023 81.55 ;
			RECT	200.243 81.486 200.275 81.55 ;
			RECT	200.9 81.486 200.932 81.55 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 0.598 201.665 0.718 ;
			LAYER	J3 ;
			RECT	0.755 0.626 0.787 0.69 ;
			RECT	1.645 0.626 1.709 0.69 ;
			RECT	2.323 0.626 2.387 0.69 ;
			RECT	3.438 0.626 3.47 0.69 ;
			RECT	3.585 0.626 3.617 0.69 ;
			RECT	4.195 0.626 4.227 0.69 ;
			RECT	4.944 0.626 5.008 0.69 ;
			RECT	5.927 0.626 5.959 0.69 ;
			RECT	6.179 0.626 6.211 0.69 ;
			RECT	6.347 0.626 6.379 0.69 ;
			RECT	6.515 0.626 6.547 0.69 ;
			RECT	6.683 0.626 6.715 0.69 ;
			RECT	6.851 0.626 6.883 0.69 ;
			RECT	7.019 0.626 7.051 0.69 ;
			RECT	7.187 0.626 7.219 0.69 ;
			RECT	7.355 0.626 7.387 0.69 ;
			RECT	7.523 0.626 7.555 0.69 ;
			RECT	7.691 0.626 7.723 0.69 ;
			RECT	7.859 0.626 7.891 0.69 ;
			RECT	8.027 0.626 8.059 0.69 ;
			RECT	8.195 0.626 8.227 0.69 ;
			RECT	8.363 0.626 8.395 0.69 ;
			RECT	8.531 0.626 8.563 0.69 ;
			RECT	8.699 0.626 8.731 0.69 ;
			RECT	8.867 0.626 8.899 0.69 ;
			RECT	9.035 0.626 9.067 0.69 ;
			RECT	9.203 0.626 9.235 0.69 ;
			RECT	9.371 0.626 9.403 0.69 ;
			RECT	9.539 0.626 9.571 0.69 ;
			RECT	9.707 0.626 9.739 0.69 ;
			RECT	9.875 0.626 9.907 0.69 ;
			RECT	10.043 0.626 10.075 0.69 ;
			RECT	10.211 0.626 10.243 0.69 ;
			RECT	10.379 0.626 10.411 0.69 ;
			RECT	10.547 0.626 10.579 0.69 ;
			RECT	10.715 0.626 10.747 0.69 ;
			RECT	10.883 0.626 10.915 0.69 ;
			RECT	11.051 0.626 11.083 0.69 ;
			RECT	11.219 0.626 11.251 0.69 ;
			RECT	11.387 0.626 11.419 0.69 ;
			RECT	11.555 0.626 11.587 0.69 ;
			RECT	11.723 0.626 11.755 0.69 ;
			RECT	11.891 0.626 11.923 0.69 ;
			RECT	12.059 0.626 12.091 0.69 ;
			RECT	12.227 0.626 12.259 0.69 ;
			RECT	12.395 0.626 12.427 0.69 ;
			RECT	12.563 0.626 12.595 0.69 ;
			RECT	12.731 0.626 12.763 0.69 ;
			RECT	12.899 0.626 12.931 0.69 ;
			RECT	13.067 0.626 13.099 0.69 ;
			RECT	13.235 0.626 13.267 0.69 ;
			RECT	13.403 0.626 13.435 0.69 ;
			RECT	13.571 0.626 13.603 0.69 ;
			RECT	13.739 0.626 13.771 0.69 ;
			RECT	13.907 0.626 13.939 0.69 ;
			RECT	14.075 0.626 14.107 0.69 ;
			RECT	14.243 0.626 14.275 0.69 ;
			RECT	14.411 0.626 14.443 0.69 ;
			RECT	14.579 0.626 14.611 0.69 ;
			RECT	14.747 0.626 14.779 0.69 ;
			RECT	14.915 0.626 14.947 0.69 ;
			RECT	15.083 0.626 15.115 0.69 ;
			RECT	15.251 0.626 15.283 0.69 ;
			RECT	15.419 0.626 15.451 0.69 ;
			RECT	15.587 0.626 15.619 0.69 ;
			RECT	15.755 0.626 15.787 0.69 ;
			RECT	15.923 0.626 15.955 0.69 ;
			RECT	16.091 0.626 16.123 0.69 ;
			RECT	16.259 0.626 16.291 0.69 ;
			RECT	16.427 0.626 16.459 0.69 ;
			RECT	16.595 0.626 16.627 0.69 ;
			RECT	16.763 0.626 16.795 0.69 ;
			RECT	16.931 0.626 16.963 0.69 ;
			RECT	17.099 0.626 17.131 0.69 ;
			RECT	17.267 0.626 17.299 0.69 ;
			RECT	17.435 0.626 17.467 0.69 ;
			RECT	17.603 0.626 17.635 0.69 ;
			RECT	17.771 0.626 17.803 0.69 ;
			RECT	17.939 0.626 17.971 0.69 ;
			RECT	18.107 0.626 18.139 0.69 ;
			RECT	18.275 0.626 18.307 0.69 ;
			RECT	18.443 0.626 18.475 0.69 ;
			RECT	18.611 0.626 18.643 0.69 ;
			RECT	18.779 0.626 18.811 0.69 ;
			RECT	18.947 0.626 18.979 0.69 ;
			RECT	19.115 0.626 19.147 0.69 ;
			RECT	19.283 0.626 19.315 0.69 ;
			RECT	19.451 0.626 19.483 0.69 ;
			RECT	19.619 0.626 19.651 0.69 ;
			RECT	19.787 0.626 19.819 0.69 ;
			RECT	19.955 0.626 19.987 0.69 ;
			RECT	20.123 0.626 20.155 0.69 ;
			RECT	20.291 0.626 20.323 0.69 ;
			RECT	20.459 0.626 20.491 0.69 ;
			RECT	20.627 0.626 20.659 0.69 ;
			RECT	20.795 0.626 20.827 0.69 ;
			RECT	20.963 0.626 20.995 0.69 ;
			RECT	21.131 0.626 21.163 0.69 ;
			RECT	21.299 0.626 21.331 0.69 ;
			RECT	21.467 0.626 21.499 0.69 ;
			RECT	21.635 0.626 21.667 0.69 ;
			RECT	21.803 0.626 21.835 0.69 ;
			RECT	21.971 0.626 22.003 0.69 ;
			RECT	22.139 0.626 22.171 0.69 ;
			RECT	22.307 0.626 22.339 0.69 ;
			RECT	22.475 0.626 22.507 0.69 ;
			RECT	22.643 0.626 22.675 0.69 ;
			RECT	22.811 0.626 22.843 0.69 ;
			RECT	22.979 0.626 23.011 0.69 ;
			RECT	23.147 0.626 23.179 0.69 ;
			RECT	23.315 0.626 23.347 0.69 ;
			RECT	23.483 0.626 23.515 0.69 ;
			RECT	23.651 0.626 23.683 0.69 ;
			RECT	23.819 0.626 23.851 0.69 ;
			RECT	23.987 0.626 24.019 0.69 ;
			RECT	24.155 0.626 24.187 0.69 ;
			RECT	24.323 0.626 24.355 0.69 ;
			RECT	24.491 0.626 24.523 0.69 ;
			RECT	24.659 0.626 24.691 0.69 ;
			RECT	24.827 0.626 24.859 0.69 ;
			RECT	24.995 0.626 25.027 0.69 ;
			RECT	25.163 0.626 25.195 0.69 ;
			RECT	25.331 0.626 25.363 0.69 ;
			RECT	25.499 0.626 25.531 0.69 ;
			RECT	25.667 0.626 25.699 0.69 ;
			RECT	25.835 0.626 25.867 0.69 ;
			RECT	26.003 0.626 26.035 0.69 ;
			RECT	26.171 0.626 26.203 0.69 ;
			RECT	26.339 0.626 26.371 0.69 ;
			RECT	26.507 0.626 26.539 0.69 ;
			RECT	26.675 0.626 26.707 0.69 ;
			RECT	26.843 0.626 26.875 0.69 ;
			RECT	27.011 0.626 27.043 0.69 ;
			RECT	27.179 0.626 27.211 0.69 ;
			RECT	27.347 0.626 27.379 0.69 ;
			RECT	27.515 0.626 27.547 0.69 ;
			RECT	27.683 0.626 27.715 0.69 ;
			RECT	27.851 0.626 27.883 0.69 ;
			RECT	28.019 0.626 28.051 0.69 ;
			RECT	28.187 0.626 28.219 0.69 ;
			RECT	28.355 0.626 28.387 0.69 ;
			RECT	28.523 0.626 28.555 0.69 ;
			RECT	28.691 0.626 28.723 0.69 ;
			RECT	28.859 0.626 28.891 0.69 ;
			RECT	29.027 0.626 29.059 0.69 ;
			RECT	29.195 0.626 29.227 0.69 ;
			RECT	29.363 0.626 29.395 0.69 ;
			RECT	29.531 0.626 29.563 0.69 ;
			RECT	29.699 0.626 29.731 0.69 ;
			RECT	29.867 0.626 29.899 0.69 ;
			RECT	30.035 0.626 30.067 0.69 ;
			RECT	30.203 0.626 30.235 0.69 ;
			RECT	30.371 0.626 30.403 0.69 ;
			RECT	30.539 0.626 30.571 0.69 ;
			RECT	30.707 0.626 30.739 0.69 ;
			RECT	30.875 0.626 30.907 0.69 ;
			RECT	31.043 0.626 31.075 0.69 ;
			RECT	31.211 0.626 31.243 0.69 ;
			RECT	31.379 0.626 31.411 0.69 ;
			RECT	31.547 0.626 31.579 0.69 ;
			RECT	31.715 0.626 31.747 0.69 ;
			RECT	31.883 0.626 31.915 0.69 ;
			RECT	32.051 0.626 32.083 0.69 ;
			RECT	32.219 0.626 32.251 0.69 ;
			RECT	32.387 0.626 32.419 0.69 ;
			RECT	32.555 0.626 32.587 0.69 ;
			RECT	32.723 0.626 32.755 0.69 ;
			RECT	32.891 0.626 32.923 0.69 ;
			RECT	33.059 0.626 33.091 0.69 ;
			RECT	33.227 0.626 33.259 0.69 ;
			RECT	33.395 0.626 33.427 0.69 ;
			RECT	33.563 0.626 33.595 0.69 ;
			RECT	33.731 0.626 33.763 0.69 ;
			RECT	33.899 0.626 33.931 0.69 ;
			RECT	34.067 0.626 34.099 0.69 ;
			RECT	34.235 0.626 34.267 0.69 ;
			RECT	34.403 0.626 34.435 0.69 ;
			RECT	34.571 0.626 34.603 0.69 ;
			RECT	34.739 0.626 34.771 0.69 ;
			RECT	34.907 0.626 34.939 0.69 ;
			RECT	35.075 0.626 35.107 0.69 ;
			RECT	35.243 0.626 35.275 0.69 ;
			RECT	35.411 0.626 35.443 0.69 ;
			RECT	35.579 0.626 35.611 0.69 ;
			RECT	35.747 0.626 35.779 0.69 ;
			RECT	35.915 0.626 35.947 0.69 ;
			RECT	36.083 0.626 36.115 0.69 ;
			RECT	36.251 0.626 36.283 0.69 ;
			RECT	36.419 0.626 36.451 0.69 ;
			RECT	36.587 0.626 36.619 0.69 ;
			RECT	36.755 0.626 36.787 0.69 ;
			RECT	36.923 0.626 36.955 0.69 ;
			RECT	37.091 0.626 37.123 0.69 ;
			RECT	37.259 0.626 37.291 0.69 ;
			RECT	37.427 0.626 37.459 0.69 ;
			RECT	37.595 0.626 37.627 0.69 ;
			RECT	37.763 0.626 37.795 0.69 ;
			RECT	37.931 0.626 37.963 0.69 ;
			RECT	38.099 0.626 38.131 0.69 ;
			RECT	38.267 0.626 38.299 0.69 ;
			RECT	38.435 0.626 38.467 0.69 ;
			RECT	38.603 0.626 38.635 0.69 ;
			RECT	38.771 0.626 38.803 0.69 ;
			RECT	38.939 0.626 38.971 0.69 ;
			RECT	39.107 0.626 39.139 0.69 ;
			RECT	39.275 0.626 39.307 0.69 ;
			RECT	39.443 0.626 39.475 0.69 ;
			RECT	39.611 0.626 39.643 0.69 ;
			RECT	39.779 0.626 39.811 0.69 ;
			RECT	39.947 0.626 39.979 0.69 ;
			RECT	40.115 0.626 40.147 0.69 ;
			RECT	40.283 0.626 40.315 0.69 ;
			RECT	40.451 0.626 40.483 0.69 ;
			RECT	40.619 0.626 40.651 0.69 ;
			RECT	40.787 0.626 40.819 0.69 ;
			RECT	40.955 0.626 40.987 0.69 ;
			RECT	41.123 0.626 41.155 0.69 ;
			RECT	41.291 0.626 41.323 0.69 ;
			RECT	41.459 0.626 41.491 0.69 ;
			RECT	41.627 0.626 41.659 0.69 ;
			RECT	41.795 0.626 41.827 0.69 ;
			RECT	41.963 0.626 41.995 0.69 ;
			RECT	42.131 0.626 42.163 0.69 ;
			RECT	42.299 0.626 42.331 0.69 ;
			RECT	42.467 0.626 42.499 0.69 ;
			RECT	42.635 0.626 42.667 0.69 ;
			RECT	42.803 0.626 42.835 0.69 ;
			RECT	42.971 0.626 43.003 0.69 ;
			RECT	43.139 0.626 43.171 0.69 ;
			RECT	43.307 0.626 43.339 0.69 ;
			RECT	43.475 0.626 43.507 0.69 ;
			RECT	43.643 0.626 43.675 0.69 ;
			RECT	43.811 0.626 43.843 0.69 ;
			RECT	43.979 0.626 44.011 0.69 ;
			RECT	44.147 0.626 44.179 0.69 ;
			RECT	44.315 0.626 44.347 0.69 ;
			RECT	44.483 0.626 44.515 0.69 ;
			RECT	44.651 0.626 44.683 0.69 ;
			RECT	44.819 0.626 44.851 0.69 ;
			RECT	44.987 0.626 45.019 0.69 ;
			RECT	45.155 0.626 45.187 0.69 ;
			RECT	45.323 0.626 45.355 0.69 ;
			RECT	45.491 0.626 45.523 0.69 ;
			RECT	45.659 0.626 45.691 0.69 ;
			RECT	45.827 0.626 45.859 0.69 ;
			RECT	45.995 0.626 46.027 0.69 ;
			RECT	46.163 0.626 46.195 0.69 ;
			RECT	46.331 0.626 46.363 0.69 ;
			RECT	46.499 0.626 46.531 0.69 ;
			RECT	46.667 0.626 46.699 0.69 ;
			RECT	46.835 0.626 46.867 0.69 ;
			RECT	47.003 0.626 47.035 0.69 ;
			RECT	47.171 0.626 47.203 0.69 ;
			RECT	47.339 0.626 47.371 0.69 ;
			RECT	47.507 0.626 47.539 0.69 ;
			RECT	47.675 0.626 47.707 0.69 ;
			RECT	47.843 0.626 47.875 0.69 ;
			RECT	48.011 0.626 48.043 0.69 ;
			RECT	48.179 0.626 48.211 0.69 ;
			RECT	48.347 0.626 48.379 0.69 ;
			RECT	48.515 0.626 48.547 0.69 ;
			RECT	48.683 0.626 48.715 0.69 ;
			RECT	48.851 0.626 48.883 0.69 ;
			RECT	49.019 0.626 49.051 0.69 ;
			RECT	49.187 0.626 49.219 0.69 ;
			RECT	49.541 0.626 49.605 0.69 ;
			RECT	52.124 0.626 52.156 0.69 ;
			RECT	52.578 0.626 52.61 0.69 ;
			RECT	53.132 0.626 53.196 0.69 ;
			RECT	53.911 0.626 53.943 0.69 ;
			RECT	54.251 0.626 54.283 0.69 ;
			RECT	55.562 0.626 55.626 0.69 ;
			RECT	58.599 0.626 58.663 0.69 ;
			RECT	58.985 0.626 59.017 0.69 ;
			RECT	59.153 0.626 59.185 0.69 ;
			RECT	59.321 0.626 59.353 0.69 ;
			RECT	59.489 0.626 59.521 0.69 ;
			RECT	59.657 0.626 59.689 0.69 ;
			RECT	59.825 0.626 59.857 0.69 ;
			RECT	59.993 0.626 60.025 0.69 ;
			RECT	60.161 0.626 60.193 0.69 ;
			RECT	60.329 0.626 60.361 0.69 ;
			RECT	60.497 0.626 60.529 0.69 ;
			RECT	60.665 0.626 60.697 0.69 ;
			RECT	60.833 0.626 60.865 0.69 ;
			RECT	61.001 0.626 61.033 0.69 ;
			RECT	61.169 0.626 61.201 0.69 ;
			RECT	61.337 0.626 61.369 0.69 ;
			RECT	61.505 0.626 61.537 0.69 ;
			RECT	61.673 0.626 61.705 0.69 ;
			RECT	61.841 0.626 61.873 0.69 ;
			RECT	62.009 0.626 62.041 0.69 ;
			RECT	62.177 0.626 62.209 0.69 ;
			RECT	62.345 0.626 62.377 0.69 ;
			RECT	62.513 0.626 62.545 0.69 ;
			RECT	62.681 0.626 62.713 0.69 ;
			RECT	62.849 0.626 62.881 0.69 ;
			RECT	63.017 0.626 63.049 0.69 ;
			RECT	63.185 0.626 63.217 0.69 ;
			RECT	63.353 0.626 63.385 0.69 ;
			RECT	63.521 0.626 63.553 0.69 ;
			RECT	63.689 0.626 63.721 0.69 ;
			RECT	63.857 0.626 63.889 0.69 ;
			RECT	64.025 0.626 64.057 0.69 ;
			RECT	64.193 0.626 64.225 0.69 ;
			RECT	64.361 0.626 64.393 0.69 ;
			RECT	64.529 0.626 64.561 0.69 ;
			RECT	64.697 0.626 64.729 0.69 ;
			RECT	64.865 0.626 64.897 0.69 ;
			RECT	65.033 0.626 65.065 0.69 ;
			RECT	65.201 0.626 65.233 0.69 ;
			RECT	65.369 0.626 65.401 0.69 ;
			RECT	65.537 0.626 65.569 0.69 ;
			RECT	65.705 0.626 65.737 0.69 ;
			RECT	65.873 0.626 65.905 0.69 ;
			RECT	66.041 0.626 66.073 0.69 ;
			RECT	66.209 0.626 66.241 0.69 ;
			RECT	66.377 0.626 66.409 0.69 ;
			RECT	66.545 0.626 66.577 0.69 ;
			RECT	66.713 0.626 66.745 0.69 ;
			RECT	66.881 0.626 66.913 0.69 ;
			RECT	67.049 0.626 67.081 0.69 ;
			RECT	67.217 0.626 67.249 0.69 ;
			RECT	67.385 0.626 67.417 0.69 ;
			RECT	67.553 0.626 67.585 0.69 ;
			RECT	67.721 0.626 67.753 0.69 ;
			RECT	67.889 0.626 67.921 0.69 ;
			RECT	68.057 0.626 68.089 0.69 ;
			RECT	68.225 0.626 68.257 0.69 ;
			RECT	68.393 0.626 68.425 0.69 ;
			RECT	68.561 0.626 68.593 0.69 ;
			RECT	68.729 0.626 68.761 0.69 ;
			RECT	68.897 0.626 68.929 0.69 ;
			RECT	69.065 0.626 69.097 0.69 ;
			RECT	69.233 0.626 69.265 0.69 ;
			RECT	69.401 0.626 69.433 0.69 ;
			RECT	69.569 0.626 69.601 0.69 ;
			RECT	69.737 0.626 69.769 0.69 ;
			RECT	69.905 0.626 69.937 0.69 ;
			RECT	70.073 0.626 70.105 0.69 ;
			RECT	70.241 0.626 70.273 0.69 ;
			RECT	70.409 0.626 70.441 0.69 ;
			RECT	70.577 0.626 70.609 0.69 ;
			RECT	70.745 0.626 70.777 0.69 ;
			RECT	70.913 0.626 70.945 0.69 ;
			RECT	71.081 0.626 71.113 0.69 ;
			RECT	71.249 0.626 71.281 0.69 ;
			RECT	71.417 0.626 71.449 0.69 ;
			RECT	71.585 0.626 71.617 0.69 ;
			RECT	71.753 0.626 71.785 0.69 ;
			RECT	71.921 0.626 71.953 0.69 ;
			RECT	72.089 0.626 72.121 0.69 ;
			RECT	72.257 0.626 72.289 0.69 ;
			RECT	72.425 0.626 72.457 0.69 ;
			RECT	72.593 0.626 72.625 0.69 ;
			RECT	72.761 0.626 72.793 0.69 ;
			RECT	72.929 0.626 72.961 0.69 ;
			RECT	73.097 0.626 73.129 0.69 ;
			RECT	73.265 0.626 73.297 0.69 ;
			RECT	73.433 0.626 73.465 0.69 ;
			RECT	73.601 0.626 73.633 0.69 ;
			RECT	73.769 0.626 73.801 0.69 ;
			RECT	73.937 0.626 73.969 0.69 ;
			RECT	74.105 0.626 74.137 0.69 ;
			RECT	74.273 0.626 74.305 0.69 ;
			RECT	74.441 0.626 74.473 0.69 ;
			RECT	74.609 0.626 74.641 0.69 ;
			RECT	74.777 0.626 74.809 0.69 ;
			RECT	74.945 0.626 74.977 0.69 ;
			RECT	75.113 0.626 75.145 0.69 ;
			RECT	75.281 0.626 75.313 0.69 ;
			RECT	75.449 0.626 75.481 0.69 ;
			RECT	75.617 0.626 75.649 0.69 ;
			RECT	75.785 0.626 75.817 0.69 ;
			RECT	75.953 0.626 75.985 0.69 ;
			RECT	76.121 0.626 76.153 0.69 ;
			RECT	76.289 0.626 76.321 0.69 ;
			RECT	76.457 0.626 76.489 0.69 ;
			RECT	76.625 0.626 76.657 0.69 ;
			RECT	76.793 0.626 76.825 0.69 ;
			RECT	76.961 0.626 76.993 0.69 ;
			RECT	77.129 0.626 77.161 0.69 ;
			RECT	77.297 0.626 77.329 0.69 ;
			RECT	77.465 0.626 77.497 0.69 ;
			RECT	77.633 0.626 77.665 0.69 ;
			RECT	77.801 0.626 77.833 0.69 ;
			RECT	77.969 0.626 78.001 0.69 ;
			RECT	78.137 0.626 78.169 0.69 ;
			RECT	78.305 0.626 78.337 0.69 ;
			RECT	78.473 0.626 78.505 0.69 ;
			RECT	78.641 0.626 78.673 0.69 ;
			RECT	78.809 0.626 78.841 0.69 ;
			RECT	78.977 0.626 79.009 0.69 ;
			RECT	79.145 0.626 79.177 0.69 ;
			RECT	79.313 0.626 79.345 0.69 ;
			RECT	79.481 0.626 79.513 0.69 ;
			RECT	79.649 0.626 79.681 0.69 ;
			RECT	79.817 0.626 79.849 0.69 ;
			RECT	79.985 0.626 80.017 0.69 ;
			RECT	80.153 0.626 80.185 0.69 ;
			RECT	80.321 0.626 80.353 0.69 ;
			RECT	80.489 0.626 80.521 0.69 ;
			RECT	80.657 0.626 80.689 0.69 ;
			RECT	80.825 0.626 80.857 0.69 ;
			RECT	80.993 0.626 81.025 0.69 ;
			RECT	81.161 0.626 81.193 0.69 ;
			RECT	81.329 0.626 81.361 0.69 ;
			RECT	81.497 0.626 81.529 0.69 ;
			RECT	81.665 0.626 81.697 0.69 ;
			RECT	81.833 0.626 81.865 0.69 ;
			RECT	82.001 0.626 82.033 0.69 ;
			RECT	82.169 0.626 82.201 0.69 ;
			RECT	82.337 0.626 82.369 0.69 ;
			RECT	82.505 0.626 82.537 0.69 ;
			RECT	82.673 0.626 82.705 0.69 ;
			RECT	82.841 0.626 82.873 0.69 ;
			RECT	83.009 0.626 83.041 0.69 ;
			RECT	83.177 0.626 83.209 0.69 ;
			RECT	83.345 0.626 83.377 0.69 ;
			RECT	83.513 0.626 83.545 0.69 ;
			RECT	83.681 0.626 83.713 0.69 ;
			RECT	83.849 0.626 83.881 0.69 ;
			RECT	84.017 0.626 84.049 0.69 ;
			RECT	84.185 0.626 84.217 0.69 ;
			RECT	84.353 0.626 84.385 0.69 ;
			RECT	84.521 0.626 84.553 0.69 ;
			RECT	84.689 0.626 84.721 0.69 ;
			RECT	84.857 0.626 84.889 0.69 ;
			RECT	85.025 0.626 85.057 0.69 ;
			RECT	85.193 0.626 85.225 0.69 ;
			RECT	85.361 0.626 85.393 0.69 ;
			RECT	85.529 0.626 85.561 0.69 ;
			RECT	85.697 0.626 85.729 0.69 ;
			RECT	85.865 0.626 85.897 0.69 ;
			RECT	86.033 0.626 86.065 0.69 ;
			RECT	86.201 0.626 86.233 0.69 ;
			RECT	86.369 0.626 86.401 0.69 ;
			RECT	86.537 0.626 86.569 0.69 ;
			RECT	86.705 0.626 86.737 0.69 ;
			RECT	86.873 0.626 86.905 0.69 ;
			RECT	87.041 0.626 87.073 0.69 ;
			RECT	87.209 0.626 87.241 0.69 ;
			RECT	87.377 0.626 87.409 0.69 ;
			RECT	87.545 0.626 87.577 0.69 ;
			RECT	87.713 0.626 87.745 0.69 ;
			RECT	87.881 0.626 87.913 0.69 ;
			RECT	88.049 0.626 88.081 0.69 ;
			RECT	88.217 0.626 88.249 0.69 ;
			RECT	88.385 0.626 88.417 0.69 ;
			RECT	88.553 0.626 88.585 0.69 ;
			RECT	88.721 0.626 88.753 0.69 ;
			RECT	88.889 0.626 88.921 0.69 ;
			RECT	89.057 0.626 89.089 0.69 ;
			RECT	89.225 0.626 89.257 0.69 ;
			RECT	89.393 0.626 89.425 0.69 ;
			RECT	89.561 0.626 89.593 0.69 ;
			RECT	89.729 0.626 89.761 0.69 ;
			RECT	89.897 0.626 89.929 0.69 ;
			RECT	90.065 0.626 90.097 0.69 ;
			RECT	90.233 0.626 90.265 0.69 ;
			RECT	90.401 0.626 90.433 0.69 ;
			RECT	90.569 0.626 90.601 0.69 ;
			RECT	90.737 0.626 90.769 0.69 ;
			RECT	90.905 0.626 90.937 0.69 ;
			RECT	91.073 0.626 91.105 0.69 ;
			RECT	91.241 0.626 91.273 0.69 ;
			RECT	91.409 0.626 91.441 0.69 ;
			RECT	91.577 0.626 91.609 0.69 ;
			RECT	91.745 0.626 91.777 0.69 ;
			RECT	91.913 0.626 91.945 0.69 ;
			RECT	92.081 0.626 92.113 0.69 ;
			RECT	92.249 0.626 92.281 0.69 ;
			RECT	92.417 0.626 92.449 0.69 ;
			RECT	92.585 0.626 92.617 0.69 ;
			RECT	92.753 0.626 92.785 0.69 ;
			RECT	92.921 0.626 92.953 0.69 ;
			RECT	93.089 0.626 93.121 0.69 ;
			RECT	93.257 0.626 93.289 0.69 ;
			RECT	93.425 0.626 93.457 0.69 ;
			RECT	93.593 0.626 93.625 0.69 ;
			RECT	93.761 0.626 93.793 0.69 ;
			RECT	93.929 0.626 93.961 0.69 ;
			RECT	94.097 0.626 94.129 0.69 ;
			RECT	94.265 0.626 94.297 0.69 ;
			RECT	94.433 0.626 94.465 0.69 ;
			RECT	94.601 0.626 94.633 0.69 ;
			RECT	94.769 0.626 94.801 0.69 ;
			RECT	94.937 0.626 94.969 0.69 ;
			RECT	95.105 0.626 95.137 0.69 ;
			RECT	95.273 0.626 95.305 0.69 ;
			RECT	95.441 0.626 95.473 0.69 ;
			RECT	95.609 0.626 95.641 0.69 ;
			RECT	95.777 0.626 95.809 0.69 ;
			RECT	95.945 0.626 95.977 0.69 ;
			RECT	96.113 0.626 96.145 0.69 ;
			RECT	96.281 0.626 96.313 0.69 ;
			RECT	96.449 0.626 96.481 0.69 ;
			RECT	96.617 0.626 96.649 0.69 ;
			RECT	96.785 0.626 96.817 0.69 ;
			RECT	96.953 0.626 96.985 0.69 ;
			RECT	97.121 0.626 97.153 0.69 ;
			RECT	97.289 0.626 97.321 0.69 ;
			RECT	97.457 0.626 97.489 0.69 ;
			RECT	97.625 0.626 97.657 0.69 ;
			RECT	97.793 0.626 97.825 0.69 ;
			RECT	97.961 0.626 97.993 0.69 ;
			RECT	98.129 0.626 98.161 0.69 ;
			RECT	98.297 0.626 98.329 0.69 ;
			RECT	98.465 0.626 98.497 0.69 ;
			RECT	98.633 0.626 98.665 0.69 ;
			RECT	98.801 0.626 98.833 0.69 ;
			RECT	98.969 0.626 99.001 0.69 ;
			RECT	99.137 0.626 99.169 0.69 ;
			RECT	99.305 0.626 99.337 0.69 ;
			RECT	99.473 0.626 99.505 0.69 ;
			RECT	99.641 0.626 99.673 0.69 ;
			RECT	99.809 0.626 99.841 0.69 ;
			RECT	99.977 0.626 100.009 0.69 ;
			RECT	100.145 0.626 100.177 0.69 ;
			RECT	100.313 0.626 100.345 0.69 ;
			RECT	100.481 0.626 100.513 0.69 ;
			RECT	100.649 0.626 100.681 0.69 ;
			RECT	100.817 0.626 100.849 0.69 ;
			RECT	100.985 0.626 101.017 0.69 ;
			RECT	101.153 0.626 101.185 0.69 ;
			RECT	101.321 0.626 101.353 0.69 ;
			RECT	101.489 0.626 101.521 0.69 ;
			RECT	101.657 0.626 101.689 0.69 ;
			RECT	101.825 0.626 101.857 0.69 ;
			RECT	101.993 0.626 102.025 0.69 ;
			RECT	102.245 0.626 102.277 0.69 ;
			RECT	103.085 0.626 103.117 0.69 ;
			RECT	103.925 0.626 103.957 0.69 ;
			RECT	104.177 0.626 104.209 0.69 ;
			RECT	104.345 0.626 104.377 0.69 ;
			RECT	104.513 0.626 104.545 0.69 ;
			RECT	104.681 0.626 104.713 0.69 ;
			RECT	104.849 0.626 104.881 0.69 ;
			RECT	105.017 0.626 105.049 0.69 ;
			RECT	105.185 0.626 105.217 0.69 ;
			RECT	105.353 0.626 105.385 0.69 ;
			RECT	105.521 0.626 105.553 0.69 ;
			RECT	105.689 0.626 105.721 0.69 ;
			RECT	105.857 0.626 105.889 0.69 ;
			RECT	106.025 0.626 106.057 0.69 ;
			RECT	106.193 0.626 106.225 0.69 ;
			RECT	106.361 0.626 106.393 0.69 ;
			RECT	106.529 0.626 106.561 0.69 ;
			RECT	106.697 0.626 106.729 0.69 ;
			RECT	106.865 0.626 106.897 0.69 ;
			RECT	107.033 0.626 107.065 0.69 ;
			RECT	107.201 0.626 107.233 0.69 ;
			RECT	107.369 0.626 107.401 0.69 ;
			RECT	107.537 0.626 107.569 0.69 ;
			RECT	107.705 0.626 107.737 0.69 ;
			RECT	107.873 0.626 107.905 0.69 ;
			RECT	108.041 0.626 108.073 0.69 ;
			RECT	108.209 0.626 108.241 0.69 ;
			RECT	108.377 0.626 108.409 0.69 ;
			RECT	108.545 0.626 108.577 0.69 ;
			RECT	108.713 0.626 108.745 0.69 ;
			RECT	108.881 0.626 108.913 0.69 ;
			RECT	109.049 0.626 109.081 0.69 ;
			RECT	109.217 0.626 109.249 0.69 ;
			RECT	109.385 0.626 109.417 0.69 ;
			RECT	109.553 0.626 109.585 0.69 ;
			RECT	109.721 0.626 109.753 0.69 ;
			RECT	109.889 0.626 109.921 0.69 ;
			RECT	110.057 0.626 110.089 0.69 ;
			RECT	110.225 0.626 110.257 0.69 ;
			RECT	110.393 0.626 110.425 0.69 ;
			RECT	110.561 0.626 110.593 0.69 ;
			RECT	110.729 0.626 110.761 0.69 ;
			RECT	110.897 0.626 110.929 0.69 ;
			RECT	111.065 0.626 111.097 0.69 ;
			RECT	111.233 0.626 111.265 0.69 ;
			RECT	111.401 0.626 111.433 0.69 ;
			RECT	111.569 0.626 111.601 0.69 ;
			RECT	111.737 0.626 111.769 0.69 ;
			RECT	111.905 0.626 111.937 0.69 ;
			RECT	112.073 0.626 112.105 0.69 ;
			RECT	112.241 0.626 112.273 0.69 ;
			RECT	112.409 0.626 112.441 0.69 ;
			RECT	112.577 0.626 112.609 0.69 ;
			RECT	112.745 0.626 112.777 0.69 ;
			RECT	112.913 0.626 112.945 0.69 ;
			RECT	113.081 0.626 113.113 0.69 ;
			RECT	113.249 0.626 113.281 0.69 ;
			RECT	113.417 0.626 113.449 0.69 ;
			RECT	113.585 0.626 113.617 0.69 ;
			RECT	113.753 0.626 113.785 0.69 ;
			RECT	113.921 0.626 113.953 0.69 ;
			RECT	114.089 0.626 114.121 0.69 ;
			RECT	114.257 0.626 114.289 0.69 ;
			RECT	114.425 0.626 114.457 0.69 ;
			RECT	114.593 0.626 114.625 0.69 ;
			RECT	114.761 0.626 114.793 0.69 ;
			RECT	114.929 0.626 114.961 0.69 ;
			RECT	115.097 0.626 115.129 0.69 ;
			RECT	115.265 0.626 115.297 0.69 ;
			RECT	115.433 0.626 115.465 0.69 ;
			RECT	115.601 0.626 115.633 0.69 ;
			RECT	115.769 0.626 115.801 0.69 ;
			RECT	115.937 0.626 115.969 0.69 ;
			RECT	116.105 0.626 116.137 0.69 ;
			RECT	116.273 0.626 116.305 0.69 ;
			RECT	116.441 0.626 116.473 0.69 ;
			RECT	116.609 0.626 116.641 0.69 ;
			RECT	116.777 0.626 116.809 0.69 ;
			RECT	116.945 0.626 116.977 0.69 ;
			RECT	117.113 0.626 117.145 0.69 ;
			RECT	117.281 0.626 117.313 0.69 ;
			RECT	117.449 0.626 117.481 0.69 ;
			RECT	117.617 0.626 117.649 0.69 ;
			RECT	117.785 0.626 117.817 0.69 ;
			RECT	117.953 0.626 117.985 0.69 ;
			RECT	118.121 0.626 118.153 0.69 ;
			RECT	118.289 0.626 118.321 0.69 ;
			RECT	118.457 0.626 118.489 0.69 ;
			RECT	118.625 0.626 118.657 0.69 ;
			RECT	118.793 0.626 118.825 0.69 ;
			RECT	118.961 0.626 118.993 0.69 ;
			RECT	119.129 0.626 119.161 0.69 ;
			RECT	119.297 0.626 119.329 0.69 ;
			RECT	119.465 0.626 119.497 0.69 ;
			RECT	119.633 0.626 119.665 0.69 ;
			RECT	119.801 0.626 119.833 0.69 ;
			RECT	119.969 0.626 120.001 0.69 ;
			RECT	120.137 0.626 120.169 0.69 ;
			RECT	120.305 0.626 120.337 0.69 ;
			RECT	120.473 0.626 120.505 0.69 ;
			RECT	120.641 0.626 120.673 0.69 ;
			RECT	120.809 0.626 120.841 0.69 ;
			RECT	120.977 0.626 121.009 0.69 ;
			RECT	121.145 0.626 121.177 0.69 ;
			RECT	121.313 0.626 121.345 0.69 ;
			RECT	121.481 0.626 121.513 0.69 ;
			RECT	121.649 0.626 121.681 0.69 ;
			RECT	121.817 0.626 121.849 0.69 ;
			RECT	121.985 0.626 122.017 0.69 ;
			RECT	122.153 0.626 122.185 0.69 ;
			RECT	122.321 0.626 122.353 0.69 ;
			RECT	122.489 0.626 122.521 0.69 ;
			RECT	122.657 0.626 122.689 0.69 ;
			RECT	122.825 0.626 122.857 0.69 ;
			RECT	122.993 0.626 123.025 0.69 ;
			RECT	123.161 0.626 123.193 0.69 ;
			RECT	123.329 0.626 123.361 0.69 ;
			RECT	123.497 0.626 123.529 0.69 ;
			RECT	123.665 0.626 123.697 0.69 ;
			RECT	123.833 0.626 123.865 0.69 ;
			RECT	124.001 0.626 124.033 0.69 ;
			RECT	124.169 0.626 124.201 0.69 ;
			RECT	124.337 0.626 124.369 0.69 ;
			RECT	124.505 0.626 124.537 0.69 ;
			RECT	124.673 0.626 124.705 0.69 ;
			RECT	124.841 0.626 124.873 0.69 ;
			RECT	125.009 0.626 125.041 0.69 ;
			RECT	125.177 0.626 125.209 0.69 ;
			RECT	125.345 0.626 125.377 0.69 ;
			RECT	125.513 0.626 125.545 0.69 ;
			RECT	125.681 0.626 125.713 0.69 ;
			RECT	125.849 0.626 125.881 0.69 ;
			RECT	126.017 0.626 126.049 0.69 ;
			RECT	126.185 0.626 126.217 0.69 ;
			RECT	126.353 0.626 126.385 0.69 ;
			RECT	126.521 0.626 126.553 0.69 ;
			RECT	126.689 0.626 126.721 0.69 ;
			RECT	126.857 0.626 126.889 0.69 ;
			RECT	127.025 0.626 127.057 0.69 ;
			RECT	127.193 0.626 127.225 0.69 ;
			RECT	127.361 0.626 127.393 0.69 ;
			RECT	127.529 0.626 127.561 0.69 ;
			RECT	127.697 0.626 127.729 0.69 ;
			RECT	127.865 0.626 127.897 0.69 ;
			RECT	128.033 0.626 128.065 0.69 ;
			RECT	128.201 0.626 128.233 0.69 ;
			RECT	128.369 0.626 128.401 0.69 ;
			RECT	128.537 0.626 128.569 0.69 ;
			RECT	128.705 0.626 128.737 0.69 ;
			RECT	128.873 0.626 128.905 0.69 ;
			RECT	129.041 0.626 129.073 0.69 ;
			RECT	129.209 0.626 129.241 0.69 ;
			RECT	129.377 0.626 129.409 0.69 ;
			RECT	129.545 0.626 129.577 0.69 ;
			RECT	129.713 0.626 129.745 0.69 ;
			RECT	129.881 0.626 129.913 0.69 ;
			RECT	130.049 0.626 130.081 0.69 ;
			RECT	130.217 0.626 130.249 0.69 ;
			RECT	130.385 0.626 130.417 0.69 ;
			RECT	130.553 0.626 130.585 0.69 ;
			RECT	130.721 0.626 130.753 0.69 ;
			RECT	130.889 0.626 130.921 0.69 ;
			RECT	131.057 0.626 131.089 0.69 ;
			RECT	131.225 0.626 131.257 0.69 ;
			RECT	131.393 0.626 131.425 0.69 ;
			RECT	131.561 0.626 131.593 0.69 ;
			RECT	131.729 0.626 131.761 0.69 ;
			RECT	131.897 0.626 131.929 0.69 ;
			RECT	132.065 0.626 132.097 0.69 ;
			RECT	132.233 0.626 132.265 0.69 ;
			RECT	132.401 0.626 132.433 0.69 ;
			RECT	132.569 0.626 132.601 0.69 ;
			RECT	132.737 0.626 132.769 0.69 ;
			RECT	132.905 0.626 132.937 0.69 ;
			RECT	133.073 0.626 133.105 0.69 ;
			RECT	133.241 0.626 133.273 0.69 ;
			RECT	133.409 0.626 133.441 0.69 ;
			RECT	133.577 0.626 133.609 0.69 ;
			RECT	133.745 0.626 133.777 0.69 ;
			RECT	133.913 0.626 133.945 0.69 ;
			RECT	134.081 0.626 134.113 0.69 ;
			RECT	134.249 0.626 134.281 0.69 ;
			RECT	134.417 0.626 134.449 0.69 ;
			RECT	134.585 0.626 134.617 0.69 ;
			RECT	134.753 0.626 134.785 0.69 ;
			RECT	134.921 0.626 134.953 0.69 ;
			RECT	135.089 0.626 135.121 0.69 ;
			RECT	135.257 0.626 135.289 0.69 ;
			RECT	135.425 0.626 135.457 0.69 ;
			RECT	135.593 0.626 135.625 0.69 ;
			RECT	135.761 0.626 135.793 0.69 ;
			RECT	135.929 0.626 135.961 0.69 ;
			RECT	136.097 0.626 136.129 0.69 ;
			RECT	136.265 0.626 136.297 0.69 ;
			RECT	136.433 0.626 136.465 0.69 ;
			RECT	136.601 0.626 136.633 0.69 ;
			RECT	136.769 0.626 136.801 0.69 ;
			RECT	136.937 0.626 136.969 0.69 ;
			RECT	137.105 0.626 137.137 0.69 ;
			RECT	137.273 0.626 137.305 0.69 ;
			RECT	137.441 0.626 137.473 0.69 ;
			RECT	137.609 0.626 137.641 0.69 ;
			RECT	137.777 0.626 137.809 0.69 ;
			RECT	137.945 0.626 137.977 0.69 ;
			RECT	138.113 0.626 138.145 0.69 ;
			RECT	138.281 0.626 138.313 0.69 ;
			RECT	138.449 0.626 138.481 0.69 ;
			RECT	138.617 0.626 138.649 0.69 ;
			RECT	138.785 0.626 138.817 0.69 ;
			RECT	138.953 0.626 138.985 0.69 ;
			RECT	139.121 0.626 139.153 0.69 ;
			RECT	139.289 0.626 139.321 0.69 ;
			RECT	139.457 0.626 139.489 0.69 ;
			RECT	139.625 0.626 139.657 0.69 ;
			RECT	139.793 0.626 139.825 0.69 ;
			RECT	139.961 0.626 139.993 0.69 ;
			RECT	140.129 0.626 140.161 0.69 ;
			RECT	140.297 0.626 140.329 0.69 ;
			RECT	140.465 0.626 140.497 0.69 ;
			RECT	140.633 0.626 140.665 0.69 ;
			RECT	140.801 0.626 140.833 0.69 ;
			RECT	140.969 0.626 141.001 0.69 ;
			RECT	141.137 0.626 141.169 0.69 ;
			RECT	141.305 0.626 141.337 0.69 ;
			RECT	141.473 0.626 141.505 0.69 ;
			RECT	141.641 0.626 141.673 0.69 ;
			RECT	141.809 0.626 141.841 0.69 ;
			RECT	141.977 0.626 142.009 0.69 ;
			RECT	142.145 0.626 142.177 0.69 ;
			RECT	142.313 0.626 142.345 0.69 ;
			RECT	142.481 0.626 142.513 0.69 ;
			RECT	142.649 0.626 142.681 0.69 ;
			RECT	142.817 0.626 142.849 0.69 ;
			RECT	142.985 0.626 143.017 0.69 ;
			RECT	143.153 0.626 143.185 0.69 ;
			RECT	143.321 0.626 143.353 0.69 ;
			RECT	143.489 0.626 143.521 0.69 ;
			RECT	143.657 0.626 143.689 0.69 ;
			RECT	143.825 0.626 143.857 0.69 ;
			RECT	143.993 0.626 144.025 0.69 ;
			RECT	144.161 0.626 144.193 0.69 ;
			RECT	144.329 0.626 144.361 0.69 ;
			RECT	144.497 0.626 144.529 0.69 ;
			RECT	144.665 0.626 144.697 0.69 ;
			RECT	144.833 0.626 144.865 0.69 ;
			RECT	145.001 0.626 145.033 0.69 ;
			RECT	145.169 0.626 145.201 0.69 ;
			RECT	145.337 0.626 145.369 0.69 ;
			RECT	145.505 0.626 145.537 0.69 ;
			RECT	145.673 0.626 145.705 0.69 ;
			RECT	145.841 0.626 145.873 0.69 ;
			RECT	146.009 0.626 146.041 0.69 ;
			RECT	146.177 0.626 146.209 0.69 ;
			RECT	146.345 0.626 146.377 0.69 ;
			RECT	146.513 0.626 146.545 0.69 ;
			RECT	146.681 0.626 146.713 0.69 ;
			RECT	146.849 0.626 146.881 0.69 ;
			RECT	147.017 0.626 147.049 0.69 ;
			RECT	147.185 0.626 147.217 0.69 ;
			RECT	147.539 0.626 147.603 0.69 ;
			RECT	150.122 0.626 150.154 0.69 ;
			RECT	150.576 0.626 150.608 0.69 ;
			RECT	151.13 0.626 151.194 0.69 ;
			RECT	151.909 0.626 151.941 0.69 ;
			RECT	152.249 0.626 152.281 0.69 ;
			RECT	153.56 0.626 153.624 0.69 ;
			RECT	156.597 0.626 156.661 0.69 ;
			RECT	156.983 0.626 157.015 0.69 ;
			RECT	157.151 0.626 157.183 0.69 ;
			RECT	157.319 0.626 157.351 0.69 ;
			RECT	157.487 0.626 157.519 0.69 ;
			RECT	157.655 0.626 157.687 0.69 ;
			RECT	157.823 0.626 157.855 0.69 ;
			RECT	157.991 0.626 158.023 0.69 ;
			RECT	158.159 0.626 158.191 0.69 ;
			RECT	158.327 0.626 158.359 0.69 ;
			RECT	158.495 0.626 158.527 0.69 ;
			RECT	158.663 0.626 158.695 0.69 ;
			RECT	158.831 0.626 158.863 0.69 ;
			RECT	158.999 0.626 159.031 0.69 ;
			RECT	159.167 0.626 159.199 0.69 ;
			RECT	159.335 0.626 159.367 0.69 ;
			RECT	159.503 0.626 159.535 0.69 ;
			RECT	159.671 0.626 159.703 0.69 ;
			RECT	159.839 0.626 159.871 0.69 ;
			RECT	160.007 0.626 160.039 0.69 ;
			RECT	160.175 0.626 160.207 0.69 ;
			RECT	160.343 0.626 160.375 0.69 ;
			RECT	160.511 0.626 160.543 0.69 ;
			RECT	160.679 0.626 160.711 0.69 ;
			RECT	160.847 0.626 160.879 0.69 ;
			RECT	161.015 0.626 161.047 0.69 ;
			RECT	161.183 0.626 161.215 0.69 ;
			RECT	161.351 0.626 161.383 0.69 ;
			RECT	161.519 0.626 161.551 0.69 ;
			RECT	161.687 0.626 161.719 0.69 ;
			RECT	161.855 0.626 161.887 0.69 ;
			RECT	162.023 0.626 162.055 0.69 ;
			RECT	162.191 0.626 162.223 0.69 ;
			RECT	162.359 0.626 162.391 0.69 ;
			RECT	162.527 0.626 162.559 0.69 ;
			RECT	162.695 0.626 162.727 0.69 ;
			RECT	162.863 0.626 162.895 0.69 ;
			RECT	163.031 0.626 163.063 0.69 ;
			RECT	163.199 0.626 163.231 0.69 ;
			RECT	163.367 0.626 163.399 0.69 ;
			RECT	163.535 0.626 163.567 0.69 ;
			RECT	163.703 0.626 163.735 0.69 ;
			RECT	163.871 0.626 163.903 0.69 ;
			RECT	164.039 0.626 164.071 0.69 ;
			RECT	164.207 0.626 164.239 0.69 ;
			RECT	164.375 0.626 164.407 0.69 ;
			RECT	164.543 0.626 164.575 0.69 ;
			RECT	164.711 0.626 164.743 0.69 ;
			RECT	164.879 0.626 164.911 0.69 ;
			RECT	165.047 0.626 165.079 0.69 ;
			RECT	165.215 0.626 165.247 0.69 ;
			RECT	165.383 0.626 165.415 0.69 ;
			RECT	165.551 0.626 165.583 0.69 ;
			RECT	165.719 0.626 165.751 0.69 ;
			RECT	165.887 0.626 165.919 0.69 ;
			RECT	166.055 0.626 166.087 0.69 ;
			RECT	166.223 0.626 166.255 0.69 ;
			RECT	166.391 0.626 166.423 0.69 ;
			RECT	166.559 0.626 166.591 0.69 ;
			RECT	166.727 0.626 166.759 0.69 ;
			RECT	166.895 0.626 166.927 0.69 ;
			RECT	167.063 0.626 167.095 0.69 ;
			RECT	167.231 0.626 167.263 0.69 ;
			RECT	167.399 0.626 167.431 0.69 ;
			RECT	167.567 0.626 167.599 0.69 ;
			RECT	167.735 0.626 167.767 0.69 ;
			RECT	167.903 0.626 167.935 0.69 ;
			RECT	168.071 0.626 168.103 0.69 ;
			RECT	168.239 0.626 168.271 0.69 ;
			RECT	168.407 0.626 168.439 0.69 ;
			RECT	168.575 0.626 168.607 0.69 ;
			RECT	168.743 0.626 168.775 0.69 ;
			RECT	168.911 0.626 168.943 0.69 ;
			RECT	169.079 0.626 169.111 0.69 ;
			RECT	169.247 0.626 169.279 0.69 ;
			RECT	169.415 0.626 169.447 0.69 ;
			RECT	169.583 0.626 169.615 0.69 ;
			RECT	169.751 0.626 169.783 0.69 ;
			RECT	169.919 0.626 169.951 0.69 ;
			RECT	170.087 0.626 170.119 0.69 ;
			RECT	170.255 0.626 170.287 0.69 ;
			RECT	170.423 0.626 170.455 0.69 ;
			RECT	170.591 0.626 170.623 0.69 ;
			RECT	170.759 0.626 170.791 0.69 ;
			RECT	170.927 0.626 170.959 0.69 ;
			RECT	171.095 0.626 171.127 0.69 ;
			RECT	171.263 0.626 171.295 0.69 ;
			RECT	171.431 0.626 171.463 0.69 ;
			RECT	171.599 0.626 171.631 0.69 ;
			RECT	171.767 0.626 171.799 0.69 ;
			RECT	171.935 0.626 171.967 0.69 ;
			RECT	172.103 0.626 172.135 0.69 ;
			RECT	172.271 0.626 172.303 0.69 ;
			RECT	172.439 0.626 172.471 0.69 ;
			RECT	172.607 0.626 172.639 0.69 ;
			RECT	172.775 0.626 172.807 0.69 ;
			RECT	172.943 0.626 172.975 0.69 ;
			RECT	173.111 0.626 173.143 0.69 ;
			RECT	173.279 0.626 173.311 0.69 ;
			RECT	173.447 0.626 173.479 0.69 ;
			RECT	173.615 0.626 173.647 0.69 ;
			RECT	173.783 0.626 173.815 0.69 ;
			RECT	173.951 0.626 173.983 0.69 ;
			RECT	174.119 0.626 174.151 0.69 ;
			RECT	174.287 0.626 174.319 0.69 ;
			RECT	174.455 0.626 174.487 0.69 ;
			RECT	174.623 0.626 174.655 0.69 ;
			RECT	174.791 0.626 174.823 0.69 ;
			RECT	174.959 0.626 174.991 0.69 ;
			RECT	175.127 0.626 175.159 0.69 ;
			RECT	175.295 0.626 175.327 0.69 ;
			RECT	175.463 0.626 175.495 0.69 ;
			RECT	175.631 0.626 175.663 0.69 ;
			RECT	175.799 0.626 175.831 0.69 ;
			RECT	175.967 0.626 175.999 0.69 ;
			RECT	176.135 0.626 176.167 0.69 ;
			RECT	176.303 0.626 176.335 0.69 ;
			RECT	176.471 0.626 176.503 0.69 ;
			RECT	176.639 0.626 176.671 0.69 ;
			RECT	176.807 0.626 176.839 0.69 ;
			RECT	176.975 0.626 177.007 0.69 ;
			RECT	177.143 0.626 177.175 0.69 ;
			RECT	177.311 0.626 177.343 0.69 ;
			RECT	177.479 0.626 177.511 0.69 ;
			RECT	177.647 0.626 177.679 0.69 ;
			RECT	177.815 0.626 177.847 0.69 ;
			RECT	177.983 0.626 178.015 0.69 ;
			RECT	178.151 0.626 178.183 0.69 ;
			RECT	178.319 0.626 178.351 0.69 ;
			RECT	178.487 0.626 178.519 0.69 ;
			RECT	178.655 0.626 178.687 0.69 ;
			RECT	178.823 0.626 178.855 0.69 ;
			RECT	178.991 0.626 179.023 0.69 ;
			RECT	179.159 0.626 179.191 0.69 ;
			RECT	179.327 0.626 179.359 0.69 ;
			RECT	179.495 0.626 179.527 0.69 ;
			RECT	179.663 0.626 179.695 0.69 ;
			RECT	179.831 0.626 179.863 0.69 ;
			RECT	179.999 0.626 180.031 0.69 ;
			RECT	180.167 0.626 180.199 0.69 ;
			RECT	180.335 0.626 180.367 0.69 ;
			RECT	180.503 0.626 180.535 0.69 ;
			RECT	180.671 0.626 180.703 0.69 ;
			RECT	180.839 0.626 180.871 0.69 ;
			RECT	181.007 0.626 181.039 0.69 ;
			RECT	181.175 0.626 181.207 0.69 ;
			RECT	181.343 0.626 181.375 0.69 ;
			RECT	181.511 0.626 181.543 0.69 ;
			RECT	181.679 0.626 181.711 0.69 ;
			RECT	181.847 0.626 181.879 0.69 ;
			RECT	182.015 0.626 182.047 0.69 ;
			RECT	182.183 0.626 182.215 0.69 ;
			RECT	182.351 0.626 182.383 0.69 ;
			RECT	182.519 0.626 182.551 0.69 ;
			RECT	182.687 0.626 182.719 0.69 ;
			RECT	182.855 0.626 182.887 0.69 ;
			RECT	183.023 0.626 183.055 0.69 ;
			RECT	183.191 0.626 183.223 0.69 ;
			RECT	183.359 0.626 183.391 0.69 ;
			RECT	183.527 0.626 183.559 0.69 ;
			RECT	183.695 0.626 183.727 0.69 ;
			RECT	183.863 0.626 183.895 0.69 ;
			RECT	184.031 0.626 184.063 0.69 ;
			RECT	184.199 0.626 184.231 0.69 ;
			RECT	184.367 0.626 184.399 0.69 ;
			RECT	184.535 0.626 184.567 0.69 ;
			RECT	184.703 0.626 184.735 0.69 ;
			RECT	184.871 0.626 184.903 0.69 ;
			RECT	185.039 0.626 185.071 0.69 ;
			RECT	185.207 0.626 185.239 0.69 ;
			RECT	185.375 0.626 185.407 0.69 ;
			RECT	185.543 0.626 185.575 0.69 ;
			RECT	185.711 0.626 185.743 0.69 ;
			RECT	185.879 0.626 185.911 0.69 ;
			RECT	186.047 0.626 186.079 0.69 ;
			RECT	186.215 0.626 186.247 0.69 ;
			RECT	186.383 0.626 186.415 0.69 ;
			RECT	186.551 0.626 186.583 0.69 ;
			RECT	186.719 0.626 186.751 0.69 ;
			RECT	186.887 0.626 186.919 0.69 ;
			RECT	187.055 0.626 187.087 0.69 ;
			RECT	187.223 0.626 187.255 0.69 ;
			RECT	187.391 0.626 187.423 0.69 ;
			RECT	187.559 0.626 187.591 0.69 ;
			RECT	187.727 0.626 187.759 0.69 ;
			RECT	187.895 0.626 187.927 0.69 ;
			RECT	188.063 0.626 188.095 0.69 ;
			RECT	188.231 0.626 188.263 0.69 ;
			RECT	188.399 0.626 188.431 0.69 ;
			RECT	188.567 0.626 188.599 0.69 ;
			RECT	188.735 0.626 188.767 0.69 ;
			RECT	188.903 0.626 188.935 0.69 ;
			RECT	189.071 0.626 189.103 0.69 ;
			RECT	189.239 0.626 189.271 0.69 ;
			RECT	189.407 0.626 189.439 0.69 ;
			RECT	189.575 0.626 189.607 0.69 ;
			RECT	189.743 0.626 189.775 0.69 ;
			RECT	189.911 0.626 189.943 0.69 ;
			RECT	190.079 0.626 190.111 0.69 ;
			RECT	190.247 0.626 190.279 0.69 ;
			RECT	190.415 0.626 190.447 0.69 ;
			RECT	190.583 0.626 190.615 0.69 ;
			RECT	190.751 0.626 190.783 0.69 ;
			RECT	190.919 0.626 190.951 0.69 ;
			RECT	191.087 0.626 191.119 0.69 ;
			RECT	191.255 0.626 191.287 0.69 ;
			RECT	191.423 0.626 191.455 0.69 ;
			RECT	191.591 0.626 191.623 0.69 ;
			RECT	191.759 0.626 191.791 0.69 ;
			RECT	191.927 0.626 191.959 0.69 ;
			RECT	192.095 0.626 192.127 0.69 ;
			RECT	192.263 0.626 192.295 0.69 ;
			RECT	192.431 0.626 192.463 0.69 ;
			RECT	192.599 0.626 192.631 0.69 ;
			RECT	192.767 0.626 192.799 0.69 ;
			RECT	192.935 0.626 192.967 0.69 ;
			RECT	193.103 0.626 193.135 0.69 ;
			RECT	193.271 0.626 193.303 0.69 ;
			RECT	193.439 0.626 193.471 0.69 ;
			RECT	193.607 0.626 193.639 0.69 ;
			RECT	193.775 0.626 193.807 0.69 ;
			RECT	193.943 0.626 193.975 0.69 ;
			RECT	194.111 0.626 194.143 0.69 ;
			RECT	194.279 0.626 194.311 0.69 ;
			RECT	194.447 0.626 194.479 0.69 ;
			RECT	194.615 0.626 194.647 0.69 ;
			RECT	194.783 0.626 194.815 0.69 ;
			RECT	194.951 0.626 194.983 0.69 ;
			RECT	195.119 0.626 195.151 0.69 ;
			RECT	195.287 0.626 195.319 0.69 ;
			RECT	195.455 0.626 195.487 0.69 ;
			RECT	195.623 0.626 195.655 0.69 ;
			RECT	195.791 0.626 195.823 0.69 ;
			RECT	195.959 0.626 195.991 0.69 ;
			RECT	196.127 0.626 196.159 0.69 ;
			RECT	196.295 0.626 196.327 0.69 ;
			RECT	196.463 0.626 196.495 0.69 ;
			RECT	196.631 0.626 196.663 0.69 ;
			RECT	196.799 0.626 196.831 0.69 ;
			RECT	196.967 0.626 196.999 0.69 ;
			RECT	197.135 0.626 197.167 0.69 ;
			RECT	197.303 0.626 197.335 0.69 ;
			RECT	197.471 0.626 197.503 0.69 ;
			RECT	197.639 0.626 197.671 0.69 ;
			RECT	197.807 0.626 197.839 0.69 ;
			RECT	197.975 0.626 198.007 0.69 ;
			RECT	198.143 0.626 198.175 0.69 ;
			RECT	198.311 0.626 198.343 0.69 ;
			RECT	198.479 0.626 198.511 0.69 ;
			RECT	198.647 0.626 198.679 0.69 ;
			RECT	198.815 0.626 198.847 0.69 ;
			RECT	198.983 0.626 199.015 0.69 ;
			RECT	199.151 0.626 199.183 0.69 ;
			RECT	199.319 0.626 199.351 0.69 ;
			RECT	199.487 0.626 199.519 0.69 ;
			RECT	199.655 0.626 199.687 0.69 ;
			RECT	199.823 0.626 199.855 0.69 ;
			RECT	199.991 0.626 200.023 0.69 ;
			RECT	200.243 0.626 200.275 0.69 ;
			RECT	200.9 0.626 200.932 0.69 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 31.908 201.665 32.018 ;
			LAYER	J3 ;
			RECT	1.645 31.931 1.709 31.995 ;
			RECT	2.129 31.931 2.161 31.995 ;
			RECT	2.323 31.931 2.387 31.995 ;
			RECT	3.438 31.931 3.47 31.995 ;
			RECT	4.195 31.931 4.227 31.995 ;
			RECT	4.96 31.931 4.992 31.995 ;
			RECT	5.252 31.931 5.284 31.995 ;
			RECT	5.927 31.931 5.959 31.995 ;
			RECT	6.179 31.931 6.211 31.995 ;
			RECT	6.347 31.931 6.379 31.995 ;
			RECT	6.515 31.931 6.547 31.995 ;
			RECT	6.683 31.931 6.715 31.995 ;
			RECT	6.851 31.931 6.883 31.995 ;
			RECT	7.019 31.931 7.051 31.995 ;
			RECT	7.187 31.931 7.219 31.995 ;
			RECT	7.355 31.931 7.387 31.995 ;
			RECT	7.523 31.931 7.555 31.995 ;
			RECT	7.691 31.931 7.723 31.995 ;
			RECT	7.859 31.931 7.891 31.995 ;
			RECT	8.027 31.931 8.059 31.995 ;
			RECT	8.195 31.931 8.227 31.995 ;
			RECT	8.363 31.931 8.395 31.995 ;
			RECT	8.531 31.931 8.563 31.995 ;
			RECT	8.699 31.931 8.731 31.995 ;
			RECT	8.867 31.931 8.899 31.995 ;
			RECT	9.035 31.931 9.067 31.995 ;
			RECT	9.203 31.931 9.235 31.995 ;
			RECT	9.371 31.931 9.403 31.995 ;
			RECT	9.539 31.931 9.571 31.995 ;
			RECT	9.707 31.931 9.739 31.995 ;
			RECT	9.875 31.931 9.907 31.995 ;
			RECT	10.043 31.931 10.075 31.995 ;
			RECT	10.211 31.931 10.243 31.995 ;
			RECT	10.379 31.931 10.411 31.995 ;
			RECT	10.547 31.931 10.579 31.995 ;
			RECT	10.715 31.931 10.747 31.995 ;
			RECT	10.883 31.931 10.915 31.995 ;
			RECT	11.051 31.931 11.083 31.995 ;
			RECT	11.219 31.931 11.251 31.995 ;
			RECT	11.387 31.931 11.419 31.995 ;
			RECT	11.555 31.931 11.587 31.995 ;
			RECT	11.723 31.931 11.755 31.995 ;
			RECT	11.891 31.931 11.923 31.995 ;
			RECT	12.059 31.931 12.091 31.995 ;
			RECT	12.227 31.931 12.259 31.995 ;
			RECT	12.395 31.931 12.427 31.995 ;
			RECT	12.563 31.931 12.595 31.995 ;
			RECT	12.731 31.931 12.763 31.995 ;
			RECT	12.899 31.931 12.931 31.995 ;
			RECT	13.067 31.931 13.099 31.995 ;
			RECT	13.235 31.931 13.267 31.995 ;
			RECT	13.403 31.931 13.435 31.995 ;
			RECT	13.571 31.931 13.603 31.995 ;
			RECT	13.739 31.931 13.771 31.995 ;
			RECT	13.907 31.931 13.939 31.995 ;
			RECT	14.075 31.931 14.107 31.995 ;
			RECT	14.243 31.931 14.275 31.995 ;
			RECT	14.411 31.931 14.443 31.995 ;
			RECT	14.579 31.931 14.611 31.995 ;
			RECT	14.747 31.931 14.779 31.995 ;
			RECT	14.915 31.931 14.947 31.995 ;
			RECT	15.083 31.931 15.115 31.995 ;
			RECT	15.251 31.931 15.283 31.995 ;
			RECT	15.419 31.931 15.451 31.995 ;
			RECT	15.587 31.931 15.619 31.995 ;
			RECT	15.755 31.931 15.787 31.995 ;
			RECT	15.923 31.931 15.955 31.995 ;
			RECT	16.091 31.931 16.123 31.995 ;
			RECT	16.259 31.931 16.291 31.995 ;
			RECT	16.427 31.931 16.459 31.995 ;
			RECT	16.595 31.931 16.627 31.995 ;
			RECT	16.763 31.931 16.795 31.995 ;
			RECT	16.931 31.931 16.963 31.995 ;
			RECT	17.099 31.931 17.131 31.995 ;
			RECT	17.267 31.931 17.299 31.995 ;
			RECT	17.435 31.931 17.467 31.995 ;
			RECT	17.603 31.931 17.635 31.995 ;
			RECT	17.771 31.931 17.803 31.995 ;
			RECT	17.939 31.931 17.971 31.995 ;
			RECT	18.107 31.931 18.139 31.995 ;
			RECT	18.275 31.931 18.307 31.995 ;
			RECT	18.443 31.931 18.475 31.995 ;
			RECT	18.611 31.931 18.643 31.995 ;
			RECT	18.779 31.931 18.811 31.995 ;
			RECT	18.947 31.931 18.979 31.995 ;
			RECT	19.115 31.931 19.147 31.995 ;
			RECT	19.283 31.931 19.315 31.995 ;
			RECT	19.451 31.931 19.483 31.995 ;
			RECT	19.619 31.931 19.651 31.995 ;
			RECT	19.787 31.931 19.819 31.995 ;
			RECT	19.955 31.931 19.987 31.995 ;
			RECT	20.123 31.931 20.155 31.995 ;
			RECT	20.291 31.931 20.323 31.995 ;
			RECT	20.459 31.931 20.491 31.995 ;
			RECT	20.627 31.931 20.659 31.995 ;
			RECT	20.795 31.931 20.827 31.995 ;
			RECT	20.963 31.931 20.995 31.995 ;
			RECT	21.131 31.931 21.163 31.995 ;
			RECT	21.299 31.931 21.331 31.995 ;
			RECT	21.467 31.931 21.499 31.995 ;
			RECT	21.635 31.931 21.667 31.995 ;
			RECT	21.803 31.931 21.835 31.995 ;
			RECT	21.971 31.931 22.003 31.995 ;
			RECT	22.139 31.931 22.171 31.995 ;
			RECT	22.307 31.931 22.339 31.995 ;
			RECT	22.475 31.931 22.507 31.995 ;
			RECT	22.643 31.931 22.675 31.995 ;
			RECT	22.811 31.931 22.843 31.995 ;
			RECT	22.979 31.931 23.011 31.995 ;
			RECT	23.147 31.931 23.179 31.995 ;
			RECT	23.315 31.931 23.347 31.995 ;
			RECT	23.483 31.931 23.515 31.995 ;
			RECT	23.651 31.931 23.683 31.995 ;
			RECT	23.819 31.931 23.851 31.995 ;
			RECT	23.987 31.931 24.019 31.995 ;
			RECT	24.155 31.931 24.187 31.995 ;
			RECT	24.323 31.931 24.355 31.995 ;
			RECT	24.491 31.931 24.523 31.995 ;
			RECT	24.659 31.931 24.691 31.995 ;
			RECT	24.827 31.931 24.859 31.995 ;
			RECT	24.995 31.931 25.027 31.995 ;
			RECT	25.163 31.931 25.195 31.995 ;
			RECT	25.331 31.931 25.363 31.995 ;
			RECT	25.499 31.931 25.531 31.995 ;
			RECT	25.667 31.931 25.699 31.995 ;
			RECT	25.835 31.931 25.867 31.995 ;
			RECT	26.003 31.931 26.035 31.995 ;
			RECT	26.171 31.931 26.203 31.995 ;
			RECT	26.339 31.931 26.371 31.995 ;
			RECT	26.507 31.931 26.539 31.995 ;
			RECT	26.675 31.931 26.707 31.995 ;
			RECT	26.843 31.931 26.875 31.995 ;
			RECT	27.011 31.931 27.043 31.995 ;
			RECT	27.179 31.931 27.211 31.995 ;
			RECT	27.347 31.931 27.379 31.995 ;
			RECT	27.515 31.931 27.547 31.995 ;
			RECT	27.683 31.931 27.715 31.995 ;
			RECT	27.851 31.931 27.883 31.995 ;
			RECT	28.019 31.931 28.051 31.995 ;
			RECT	28.187 31.931 28.219 31.995 ;
			RECT	28.355 31.931 28.387 31.995 ;
			RECT	28.523 31.931 28.555 31.995 ;
			RECT	28.691 31.931 28.723 31.995 ;
			RECT	28.859 31.931 28.891 31.995 ;
			RECT	29.027 31.931 29.059 31.995 ;
			RECT	29.195 31.931 29.227 31.995 ;
			RECT	29.363 31.931 29.395 31.995 ;
			RECT	29.531 31.931 29.563 31.995 ;
			RECT	29.699 31.931 29.731 31.995 ;
			RECT	29.867 31.931 29.899 31.995 ;
			RECT	30.035 31.931 30.067 31.995 ;
			RECT	30.203 31.931 30.235 31.995 ;
			RECT	30.371 31.931 30.403 31.995 ;
			RECT	30.539 31.931 30.571 31.995 ;
			RECT	30.707 31.931 30.739 31.995 ;
			RECT	30.875 31.931 30.907 31.995 ;
			RECT	31.043 31.931 31.075 31.995 ;
			RECT	31.211 31.931 31.243 31.995 ;
			RECT	31.379 31.931 31.411 31.995 ;
			RECT	31.547 31.931 31.579 31.995 ;
			RECT	31.715 31.931 31.747 31.995 ;
			RECT	31.883 31.931 31.915 31.995 ;
			RECT	32.051 31.931 32.083 31.995 ;
			RECT	32.219 31.931 32.251 31.995 ;
			RECT	32.387 31.931 32.419 31.995 ;
			RECT	32.555 31.931 32.587 31.995 ;
			RECT	32.723 31.931 32.755 31.995 ;
			RECT	32.891 31.931 32.923 31.995 ;
			RECT	33.059 31.931 33.091 31.995 ;
			RECT	33.227 31.931 33.259 31.995 ;
			RECT	33.395 31.931 33.427 31.995 ;
			RECT	33.563 31.931 33.595 31.995 ;
			RECT	33.731 31.931 33.763 31.995 ;
			RECT	33.899 31.931 33.931 31.995 ;
			RECT	34.067 31.931 34.099 31.995 ;
			RECT	34.235 31.931 34.267 31.995 ;
			RECT	34.403 31.931 34.435 31.995 ;
			RECT	34.571 31.931 34.603 31.995 ;
			RECT	34.739 31.931 34.771 31.995 ;
			RECT	34.907 31.931 34.939 31.995 ;
			RECT	35.075 31.931 35.107 31.995 ;
			RECT	35.243 31.931 35.275 31.995 ;
			RECT	35.411 31.931 35.443 31.995 ;
			RECT	35.579 31.931 35.611 31.995 ;
			RECT	35.747 31.931 35.779 31.995 ;
			RECT	35.915 31.931 35.947 31.995 ;
			RECT	36.083 31.931 36.115 31.995 ;
			RECT	36.251 31.931 36.283 31.995 ;
			RECT	36.419 31.931 36.451 31.995 ;
			RECT	36.587 31.931 36.619 31.995 ;
			RECT	36.755 31.931 36.787 31.995 ;
			RECT	36.923 31.931 36.955 31.995 ;
			RECT	37.091 31.931 37.123 31.995 ;
			RECT	37.259 31.931 37.291 31.995 ;
			RECT	37.427 31.931 37.459 31.995 ;
			RECT	37.595 31.931 37.627 31.995 ;
			RECT	37.763 31.931 37.795 31.995 ;
			RECT	37.931 31.931 37.963 31.995 ;
			RECT	38.099 31.931 38.131 31.995 ;
			RECT	38.267 31.931 38.299 31.995 ;
			RECT	38.435 31.931 38.467 31.995 ;
			RECT	38.603 31.931 38.635 31.995 ;
			RECT	38.771 31.931 38.803 31.995 ;
			RECT	38.939 31.931 38.971 31.995 ;
			RECT	39.107 31.931 39.139 31.995 ;
			RECT	39.275 31.931 39.307 31.995 ;
			RECT	39.443 31.931 39.475 31.995 ;
			RECT	39.611 31.931 39.643 31.995 ;
			RECT	39.779 31.931 39.811 31.995 ;
			RECT	39.947 31.931 39.979 31.995 ;
			RECT	40.115 31.931 40.147 31.995 ;
			RECT	40.283 31.931 40.315 31.995 ;
			RECT	40.451 31.931 40.483 31.995 ;
			RECT	40.619 31.931 40.651 31.995 ;
			RECT	40.787 31.931 40.819 31.995 ;
			RECT	40.955 31.931 40.987 31.995 ;
			RECT	41.123 31.931 41.155 31.995 ;
			RECT	41.291 31.931 41.323 31.995 ;
			RECT	41.459 31.931 41.491 31.995 ;
			RECT	41.627 31.931 41.659 31.995 ;
			RECT	41.795 31.931 41.827 31.995 ;
			RECT	41.963 31.931 41.995 31.995 ;
			RECT	42.131 31.931 42.163 31.995 ;
			RECT	42.299 31.931 42.331 31.995 ;
			RECT	42.467 31.931 42.499 31.995 ;
			RECT	42.635 31.931 42.667 31.995 ;
			RECT	42.803 31.931 42.835 31.995 ;
			RECT	42.971 31.931 43.003 31.995 ;
			RECT	43.139 31.931 43.171 31.995 ;
			RECT	43.307 31.931 43.339 31.995 ;
			RECT	43.475 31.931 43.507 31.995 ;
			RECT	43.643 31.931 43.675 31.995 ;
			RECT	43.811 31.931 43.843 31.995 ;
			RECT	43.979 31.931 44.011 31.995 ;
			RECT	44.147 31.931 44.179 31.995 ;
			RECT	44.315 31.931 44.347 31.995 ;
			RECT	44.483 31.931 44.515 31.995 ;
			RECT	44.651 31.931 44.683 31.995 ;
			RECT	44.819 31.931 44.851 31.995 ;
			RECT	44.987 31.931 45.019 31.995 ;
			RECT	45.155 31.931 45.187 31.995 ;
			RECT	45.323 31.931 45.355 31.995 ;
			RECT	45.491 31.931 45.523 31.995 ;
			RECT	45.659 31.931 45.691 31.995 ;
			RECT	45.827 31.931 45.859 31.995 ;
			RECT	45.995 31.931 46.027 31.995 ;
			RECT	46.163 31.931 46.195 31.995 ;
			RECT	46.331 31.931 46.363 31.995 ;
			RECT	46.499 31.931 46.531 31.995 ;
			RECT	46.667 31.931 46.699 31.995 ;
			RECT	46.835 31.931 46.867 31.995 ;
			RECT	47.003 31.931 47.035 31.995 ;
			RECT	47.171 31.931 47.203 31.995 ;
			RECT	47.339 31.931 47.371 31.995 ;
			RECT	47.507 31.931 47.539 31.995 ;
			RECT	47.675 31.931 47.707 31.995 ;
			RECT	47.843 31.931 47.875 31.995 ;
			RECT	48.011 31.931 48.043 31.995 ;
			RECT	48.179 31.931 48.211 31.995 ;
			RECT	48.347 31.931 48.379 31.995 ;
			RECT	48.515 31.931 48.547 31.995 ;
			RECT	48.683 31.931 48.715 31.995 ;
			RECT	48.851 31.931 48.883 31.995 ;
			RECT	49.019 31.931 49.051 31.995 ;
			RECT	49.187 31.931 49.219 31.995 ;
			RECT	49.439 31.931 49.471 31.995 ;
			RECT	51.92 31.931 51.952 31.995 ;
			RECT	53.91 31.93 53.942 31.994 ;
			RECT	55.969 31.93 56.033 31.994 ;
			RECT	57.254 31.931 57.286 31.995 ;
			RECT	58.733 31.931 58.765 31.995 ;
			RECT	58.985 31.931 59.017 31.995 ;
			RECT	59.153 31.931 59.185 31.995 ;
			RECT	59.321 31.931 59.353 31.995 ;
			RECT	59.489 31.931 59.521 31.995 ;
			RECT	59.657 31.931 59.689 31.995 ;
			RECT	59.825 31.931 59.857 31.995 ;
			RECT	59.993 31.931 60.025 31.995 ;
			RECT	60.161 31.931 60.193 31.995 ;
			RECT	60.329 31.931 60.361 31.995 ;
			RECT	60.497 31.931 60.529 31.995 ;
			RECT	60.665 31.931 60.697 31.995 ;
			RECT	60.833 31.931 60.865 31.995 ;
			RECT	61.001 31.931 61.033 31.995 ;
			RECT	61.169 31.931 61.201 31.995 ;
			RECT	61.337 31.931 61.369 31.995 ;
			RECT	61.505 31.931 61.537 31.995 ;
			RECT	61.673 31.931 61.705 31.995 ;
			RECT	61.841 31.931 61.873 31.995 ;
			RECT	62.009 31.931 62.041 31.995 ;
			RECT	62.177 31.931 62.209 31.995 ;
			RECT	62.345 31.931 62.377 31.995 ;
			RECT	62.513 31.931 62.545 31.995 ;
			RECT	62.681 31.931 62.713 31.995 ;
			RECT	62.849 31.931 62.881 31.995 ;
			RECT	63.017 31.931 63.049 31.995 ;
			RECT	63.185 31.931 63.217 31.995 ;
			RECT	63.353 31.931 63.385 31.995 ;
			RECT	63.521 31.931 63.553 31.995 ;
			RECT	63.689 31.931 63.721 31.995 ;
			RECT	63.857 31.931 63.889 31.995 ;
			RECT	64.025 31.931 64.057 31.995 ;
			RECT	64.193 31.931 64.225 31.995 ;
			RECT	64.361 31.931 64.393 31.995 ;
			RECT	64.529 31.931 64.561 31.995 ;
			RECT	64.697 31.931 64.729 31.995 ;
			RECT	64.865 31.931 64.897 31.995 ;
			RECT	65.033 31.931 65.065 31.995 ;
			RECT	65.201 31.931 65.233 31.995 ;
			RECT	65.369 31.931 65.401 31.995 ;
			RECT	65.537 31.931 65.569 31.995 ;
			RECT	65.705 31.931 65.737 31.995 ;
			RECT	65.873 31.931 65.905 31.995 ;
			RECT	66.041 31.931 66.073 31.995 ;
			RECT	66.209 31.931 66.241 31.995 ;
			RECT	66.377 31.931 66.409 31.995 ;
			RECT	66.545 31.931 66.577 31.995 ;
			RECT	66.713 31.931 66.745 31.995 ;
			RECT	66.881 31.931 66.913 31.995 ;
			RECT	67.049 31.931 67.081 31.995 ;
			RECT	67.217 31.931 67.249 31.995 ;
			RECT	67.385 31.931 67.417 31.995 ;
			RECT	67.553 31.931 67.585 31.995 ;
			RECT	67.721 31.931 67.753 31.995 ;
			RECT	67.889 31.931 67.921 31.995 ;
			RECT	68.057 31.931 68.089 31.995 ;
			RECT	68.225 31.931 68.257 31.995 ;
			RECT	68.393 31.931 68.425 31.995 ;
			RECT	68.561 31.931 68.593 31.995 ;
			RECT	68.729 31.931 68.761 31.995 ;
			RECT	68.897 31.931 68.929 31.995 ;
			RECT	69.065 31.931 69.097 31.995 ;
			RECT	69.233 31.931 69.265 31.995 ;
			RECT	69.401 31.931 69.433 31.995 ;
			RECT	69.569 31.931 69.601 31.995 ;
			RECT	69.737 31.931 69.769 31.995 ;
			RECT	69.905 31.931 69.937 31.995 ;
			RECT	70.073 31.931 70.105 31.995 ;
			RECT	70.241 31.931 70.273 31.995 ;
			RECT	70.409 31.931 70.441 31.995 ;
			RECT	70.577 31.931 70.609 31.995 ;
			RECT	70.745 31.931 70.777 31.995 ;
			RECT	70.913 31.931 70.945 31.995 ;
			RECT	71.081 31.931 71.113 31.995 ;
			RECT	71.249 31.931 71.281 31.995 ;
			RECT	71.417 31.931 71.449 31.995 ;
			RECT	71.585 31.931 71.617 31.995 ;
			RECT	71.753 31.931 71.785 31.995 ;
			RECT	71.921 31.931 71.953 31.995 ;
			RECT	72.089 31.931 72.121 31.995 ;
			RECT	72.257 31.931 72.289 31.995 ;
			RECT	72.425 31.931 72.457 31.995 ;
			RECT	72.593 31.931 72.625 31.995 ;
			RECT	72.761 31.931 72.793 31.995 ;
			RECT	72.929 31.931 72.961 31.995 ;
			RECT	73.097 31.931 73.129 31.995 ;
			RECT	73.265 31.931 73.297 31.995 ;
			RECT	73.433 31.931 73.465 31.995 ;
			RECT	73.601 31.931 73.633 31.995 ;
			RECT	73.769 31.931 73.801 31.995 ;
			RECT	73.937 31.931 73.969 31.995 ;
			RECT	74.105 31.931 74.137 31.995 ;
			RECT	74.273 31.931 74.305 31.995 ;
			RECT	74.441 31.931 74.473 31.995 ;
			RECT	74.609 31.931 74.641 31.995 ;
			RECT	74.777 31.931 74.809 31.995 ;
			RECT	74.945 31.931 74.977 31.995 ;
			RECT	75.113 31.931 75.145 31.995 ;
			RECT	75.281 31.931 75.313 31.995 ;
			RECT	75.449 31.931 75.481 31.995 ;
			RECT	75.617 31.931 75.649 31.995 ;
			RECT	75.785 31.931 75.817 31.995 ;
			RECT	75.953 31.931 75.985 31.995 ;
			RECT	76.121 31.931 76.153 31.995 ;
			RECT	76.289 31.931 76.321 31.995 ;
			RECT	76.457 31.931 76.489 31.995 ;
			RECT	76.625 31.931 76.657 31.995 ;
			RECT	76.793 31.931 76.825 31.995 ;
			RECT	76.961 31.931 76.993 31.995 ;
			RECT	77.129 31.931 77.161 31.995 ;
			RECT	77.297 31.931 77.329 31.995 ;
			RECT	77.465 31.931 77.497 31.995 ;
			RECT	77.633 31.931 77.665 31.995 ;
			RECT	77.801 31.931 77.833 31.995 ;
			RECT	77.969 31.931 78.001 31.995 ;
			RECT	78.137 31.931 78.169 31.995 ;
			RECT	78.305 31.931 78.337 31.995 ;
			RECT	78.473 31.931 78.505 31.995 ;
			RECT	78.641 31.931 78.673 31.995 ;
			RECT	78.809 31.931 78.841 31.995 ;
			RECT	78.977 31.931 79.009 31.995 ;
			RECT	79.145 31.931 79.177 31.995 ;
			RECT	79.313 31.931 79.345 31.995 ;
			RECT	79.481 31.931 79.513 31.995 ;
			RECT	79.649 31.931 79.681 31.995 ;
			RECT	79.817 31.931 79.849 31.995 ;
			RECT	79.985 31.931 80.017 31.995 ;
			RECT	80.153 31.931 80.185 31.995 ;
			RECT	80.321 31.931 80.353 31.995 ;
			RECT	80.489 31.931 80.521 31.995 ;
			RECT	80.657 31.931 80.689 31.995 ;
			RECT	80.825 31.931 80.857 31.995 ;
			RECT	80.993 31.931 81.025 31.995 ;
			RECT	81.161 31.931 81.193 31.995 ;
			RECT	81.329 31.931 81.361 31.995 ;
			RECT	81.497 31.931 81.529 31.995 ;
			RECT	81.665 31.931 81.697 31.995 ;
			RECT	81.833 31.931 81.865 31.995 ;
			RECT	82.001 31.931 82.033 31.995 ;
			RECT	82.169 31.931 82.201 31.995 ;
			RECT	82.337 31.931 82.369 31.995 ;
			RECT	82.505 31.931 82.537 31.995 ;
			RECT	82.673 31.931 82.705 31.995 ;
			RECT	82.841 31.931 82.873 31.995 ;
			RECT	83.009 31.931 83.041 31.995 ;
			RECT	83.177 31.931 83.209 31.995 ;
			RECT	83.345 31.931 83.377 31.995 ;
			RECT	83.513 31.931 83.545 31.995 ;
			RECT	83.681 31.931 83.713 31.995 ;
			RECT	83.849 31.931 83.881 31.995 ;
			RECT	84.017 31.931 84.049 31.995 ;
			RECT	84.185 31.931 84.217 31.995 ;
			RECT	84.353 31.931 84.385 31.995 ;
			RECT	84.521 31.931 84.553 31.995 ;
			RECT	84.689 31.931 84.721 31.995 ;
			RECT	84.857 31.931 84.889 31.995 ;
			RECT	85.025 31.931 85.057 31.995 ;
			RECT	85.193 31.931 85.225 31.995 ;
			RECT	85.361 31.931 85.393 31.995 ;
			RECT	85.529 31.931 85.561 31.995 ;
			RECT	85.697 31.931 85.729 31.995 ;
			RECT	85.865 31.931 85.897 31.995 ;
			RECT	86.033 31.931 86.065 31.995 ;
			RECT	86.201 31.931 86.233 31.995 ;
			RECT	86.369 31.931 86.401 31.995 ;
			RECT	86.537 31.931 86.569 31.995 ;
			RECT	86.705 31.931 86.737 31.995 ;
			RECT	86.873 31.931 86.905 31.995 ;
			RECT	87.041 31.931 87.073 31.995 ;
			RECT	87.209 31.931 87.241 31.995 ;
			RECT	87.377 31.931 87.409 31.995 ;
			RECT	87.545 31.931 87.577 31.995 ;
			RECT	87.713 31.931 87.745 31.995 ;
			RECT	87.881 31.931 87.913 31.995 ;
			RECT	88.049 31.931 88.081 31.995 ;
			RECT	88.217 31.931 88.249 31.995 ;
			RECT	88.385 31.931 88.417 31.995 ;
			RECT	88.553 31.931 88.585 31.995 ;
			RECT	88.721 31.931 88.753 31.995 ;
			RECT	88.889 31.931 88.921 31.995 ;
			RECT	89.057 31.931 89.089 31.995 ;
			RECT	89.225 31.931 89.257 31.995 ;
			RECT	89.393 31.931 89.425 31.995 ;
			RECT	89.561 31.931 89.593 31.995 ;
			RECT	89.729 31.931 89.761 31.995 ;
			RECT	89.897 31.931 89.929 31.995 ;
			RECT	90.065 31.931 90.097 31.995 ;
			RECT	90.233 31.931 90.265 31.995 ;
			RECT	90.401 31.931 90.433 31.995 ;
			RECT	90.569 31.931 90.601 31.995 ;
			RECT	90.737 31.931 90.769 31.995 ;
			RECT	90.905 31.931 90.937 31.995 ;
			RECT	91.073 31.931 91.105 31.995 ;
			RECT	91.241 31.931 91.273 31.995 ;
			RECT	91.409 31.931 91.441 31.995 ;
			RECT	91.577 31.931 91.609 31.995 ;
			RECT	91.745 31.931 91.777 31.995 ;
			RECT	91.913 31.931 91.945 31.995 ;
			RECT	92.081 31.931 92.113 31.995 ;
			RECT	92.249 31.931 92.281 31.995 ;
			RECT	92.417 31.931 92.449 31.995 ;
			RECT	92.585 31.931 92.617 31.995 ;
			RECT	92.753 31.931 92.785 31.995 ;
			RECT	92.921 31.931 92.953 31.995 ;
			RECT	93.089 31.931 93.121 31.995 ;
			RECT	93.257 31.931 93.289 31.995 ;
			RECT	93.425 31.931 93.457 31.995 ;
			RECT	93.593 31.931 93.625 31.995 ;
			RECT	93.761 31.931 93.793 31.995 ;
			RECT	93.929 31.931 93.961 31.995 ;
			RECT	94.097 31.931 94.129 31.995 ;
			RECT	94.265 31.931 94.297 31.995 ;
			RECT	94.433 31.931 94.465 31.995 ;
			RECT	94.601 31.931 94.633 31.995 ;
			RECT	94.769 31.931 94.801 31.995 ;
			RECT	94.937 31.931 94.969 31.995 ;
			RECT	95.105 31.931 95.137 31.995 ;
			RECT	95.273 31.931 95.305 31.995 ;
			RECT	95.441 31.931 95.473 31.995 ;
			RECT	95.609 31.931 95.641 31.995 ;
			RECT	95.777 31.931 95.809 31.995 ;
			RECT	95.945 31.931 95.977 31.995 ;
			RECT	96.113 31.931 96.145 31.995 ;
			RECT	96.281 31.931 96.313 31.995 ;
			RECT	96.449 31.931 96.481 31.995 ;
			RECT	96.617 31.931 96.649 31.995 ;
			RECT	96.785 31.931 96.817 31.995 ;
			RECT	96.953 31.931 96.985 31.995 ;
			RECT	97.121 31.931 97.153 31.995 ;
			RECT	97.289 31.931 97.321 31.995 ;
			RECT	97.457 31.931 97.489 31.995 ;
			RECT	97.625 31.931 97.657 31.995 ;
			RECT	97.793 31.931 97.825 31.995 ;
			RECT	97.961 31.931 97.993 31.995 ;
			RECT	98.129 31.931 98.161 31.995 ;
			RECT	98.297 31.931 98.329 31.995 ;
			RECT	98.465 31.931 98.497 31.995 ;
			RECT	98.633 31.931 98.665 31.995 ;
			RECT	98.801 31.931 98.833 31.995 ;
			RECT	98.969 31.931 99.001 31.995 ;
			RECT	99.137 31.931 99.169 31.995 ;
			RECT	99.305 31.931 99.337 31.995 ;
			RECT	99.473 31.931 99.505 31.995 ;
			RECT	99.641 31.931 99.673 31.995 ;
			RECT	99.809 31.931 99.841 31.995 ;
			RECT	99.977 31.931 100.009 31.995 ;
			RECT	100.145 31.931 100.177 31.995 ;
			RECT	100.313 31.931 100.345 31.995 ;
			RECT	100.481 31.931 100.513 31.995 ;
			RECT	100.649 31.931 100.681 31.995 ;
			RECT	100.817 31.931 100.849 31.995 ;
			RECT	100.985 31.931 101.017 31.995 ;
			RECT	101.153 31.931 101.185 31.995 ;
			RECT	101.321 31.931 101.353 31.995 ;
			RECT	101.489 31.931 101.521 31.995 ;
			RECT	101.657 31.931 101.689 31.995 ;
			RECT	101.825 31.931 101.857 31.995 ;
			RECT	101.993 31.931 102.025 31.995 ;
			RECT	102.245 31.931 102.277 31.995 ;
			RECT	103.085 31.931 103.117 31.995 ;
			RECT	103.925 31.931 103.957 31.995 ;
			RECT	104.177 31.931 104.209 31.995 ;
			RECT	104.345 31.931 104.377 31.995 ;
			RECT	104.513 31.931 104.545 31.995 ;
			RECT	104.681 31.931 104.713 31.995 ;
			RECT	104.849 31.931 104.881 31.995 ;
			RECT	105.017 31.931 105.049 31.995 ;
			RECT	105.185 31.931 105.217 31.995 ;
			RECT	105.353 31.931 105.385 31.995 ;
			RECT	105.521 31.931 105.553 31.995 ;
			RECT	105.689 31.931 105.721 31.995 ;
			RECT	105.857 31.931 105.889 31.995 ;
			RECT	106.025 31.931 106.057 31.995 ;
			RECT	106.193 31.931 106.225 31.995 ;
			RECT	106.361 31.931 106.393 31.995 ;
			RECT	106.529 31.931 106.561 31.995 ;
			RECT	106.697 31.931 106.729 31.995 ;
			RECT	106.865 31.931 106.897 31.995 ;
			RECT	107.033 31.931 107.065 31.995 ;
			RECT	107.201 31.931 107.233 31.995 ;
			RECT	107.369 31.931 107.401 31.995 ;
			RECT	107.537 31.931 107.569 31.995 ;
			RECT	107.705 31.931 107.737 31.995 ;
			RECT	107.873 31.931 107.905 31.995 ;
			RECT	108.041 31.931 108.073 31.995 ;
			RECT	108.209 31.931 108.241 31.995 ;
			RECT	108.377 31.931 108.409 31.995 ;
			RECT	108.545 31.931 108.577 31.995 ;
			RECT	108.713 31.931 108.745 31.995 ;
			RECT	108.881 31.931 108.913 31.995 ;
			RECT	109.049 31.931 109.081 31.995 ;
			RECT	109.217 31.931 109.249 31.995 ;
			RECT	109.385 31.931 109.417 31.995 ;
			RECT	109.553 31.931 109.585 31.995 ;
			RECT	109.721 31.931 109.753 31.995 ;
			RECT	109.889 31.931 109.921 31.995 ;
			RECT	110.057 31.931 110.089 31.995 ;
			RECT	110.225 31.931 110.257 31.995 ;
			RECT	110.393 31.931 110.425 31.995 ;
			RECT	110.561 31.931 110.593 31.995 ;
			RECT	110.729 31.931 110.761 31.995 ;
			RECT	110.897 31.931 110.929 31.995 ;
			RECT	111.065 31.931 111.097 31.995 ;
			RECT	111.233 31.931 111.265 31.995 ;
			RECT	111.401 31.931 111.433 31.995 ;
			RECT	111.569 31.931 111.601 31.995 ;
			RECT	111.737 31.931 111.769 31.995 ;
			RECT	111.905 31.931 111.937 31.995 ;
			RECT	112.073 31.931 112.105 31.995 ;
			RECT	112.241 31.931 112.273 31.995 ;
			RECT	112.409 31.931 112.441 31.995 ;
			RECT	112.577 31.931 112.609 31.995 ;
			RECT	112.745 31.931 112.777 31.995 ;
			RECT	112.913 31.931 112.945 31.995 ;
			RECT	113.081 31.931 113.113 31.995 ;
			RECT	113.249 31.931 113.281 31.995 ;
			RECT	113.417 31.931 113.449 31.995 ;
			RECT	113.585 31.931 113.617 31.995 ;
			RECT	113.753 31.931 113.785 31.995 ;
			RECT	113.921 31.931 113.953 31.995 ;
			RECT	114.089 31.931 114.121 31.995 ;
			RECT	114.257 31.931 114.289 31.995 ;
			RECT	114.425 31.931 114.457 31.995 ;
			RECT	114.593 31.931 114.625 31.995 ;
			RECT	114.761 31.931 114.793 31.995 ;
			RECT	114.929 31.931 114.961 31.995 ;
			RECT	115.097 31.931 115.129 31.995 ;
			RECT	115.265 31.931 115.297 31.995 ;
			RECT	115.433 31.931 115.465 31.995 ;
			RECT	115.601 31.931 115.633 31.995 ;
			RECT	115.769 31.931 115.801 31.995 ;
			RECT	115.937 31.931 115.969 31.995 ;
			RECT	116.105 31.931 116.137 31.995 ;
			RECT	116.273 31.931 116.305 31.995 ;
			RECT	116.441 31.931 116.473 31.995 ;
			RECT	116.609 31.931 116.641 31.995 ;
			RECT	116.777 31.931 116.809 31.995 ;
			RECT	116.945 31.931 116.977 31.995 ;
			RECT	117.113 31.931 117.145 31.995 ;
			RECT	117.281 31.931 117.313 31.995 ;
			RECT	117.449 31.931 117.481 31.995 ;
			RECT	117.617 31.931 117.649 31.995 ;
			RECT	117.785 31.931 117.817 31.995 ;
			RECT	117.953 31.931 117.985 31.995 ;
			RECT	118.121 31.931 118.153 31.995 ;
			RECT	118.289 31.931 118.321 31.995 ;
			RECT	118.457 31.931 118.489 31.995 ;
			RECT	118.625 31.931 118.657 31.995 ;
			RECT	118.793 31.931 118.825 31.995 ;
			RECT	118.961 31.931 118.993 31.995 ;
			RECT	119.129 31.931 119.161 31.995 ;
			RECT	119.297 31.931 119.329 31.995 ;
			RECT	119.465 31.931 119.497 31.995 ;
			RECT	119.633 31.931 119.665 31.995 ;
			RECT	119.801 31.931 119.833 31.995 ;
			RECT	119.969 31.931 120.001 31.995 ;
			RECT	120.137 31.931 120.169 31.995 ;
			RECT	120.305 31.931 120.337 31.995 ;
			RECT	120.473 31.931 120.505 31.995 ;
			RECT	120.641 31.931 120.673 31.995 ;
			RECT	120.809 31.931 120.841 31.995 ;
			RECT	120.977 31.931 121.009 31.995 ;
			RECT	121.145 31.931 121.177 31.995 ;
			RECT	121.313 31.931 121.345 31.995 ;
			RECT	121.481 31.931 121.513 31.995 ;
			RECT	121.649 31.931 121.681 31.995 ;
			RECT	121.817 31.931 121.849 31.995 ;
			RECT	121.985 31.931 122.017 31.995 ;
			RECT	122.153 31.931 122.185 31.995 ;
			RECT	122.321 31.931 122.353 31.995 ;
			RECT	122.489 31.931 122.521 31.995 ;
			RECT	122.657 31.931 122.689 31.995 ;
			RECT	122.825 31.931 122.857 31.995 ;
			RECT	122.993 31.931 123.025 31.995 ;
			RECT	123.161 31.931 123.193 31.995 ;
			RECT	123.329 31.931 123.361 31.995 ;
			RECT	123.497 31.931 123.529 31.995 ;
			RECT	123.665 31.931 123.697 31.995 ;
			RECT	123.833 31.931 123.865 31.995 ;
			RECT	124.001 31.931 124.033 31.995 ;
			RECT	124.169 31.931 124.201 31.995 ;
			RECT	124.337 31.931 124.369 31.995 ;
			RECT	124.505 31.931 124.537 31.995 ;
			RECT	124.673 31.931 124.705 31.995 ;
			RECT	124.841 31.931 124.873 31.995 ;
			RECT	125.009 31.931 125.041 31.995 ;
			RECT	125.177 31.931 125.209 31.995 ;
			RECT	125.345 31.931 125.377 31.995 ;
			RECT	125.513 31.931 125.545 31.995 ;
			RECT	125.681 31.931 125.713 31.995 ;
			RECT	125.849 31.931 125.881 31.995 ;
			RECT	126.017 31.931 126.049 31.995 ;
			RECT	126.185 31.931 126.217 31.995 ;
			RECT	126.353 31.931 126.385 31.995 ;
			RECT	126.521 31.931 126.553 31.995 ;
			RECT	126.689 31.931 126.721 31.995 ;
			RECT	126.857 31.931 126.889 31.995 ;
			RECT	127.025 31.931 127.057 31.995 ;
			RECT	127.193 31.931 127.225 31.995 ;
			RECT	127.361 31.931 127.393 31.995 ;
			RECT	127.529 31.931 127.561 31.995 ;
			RECT	127.697 31.931 127.729 31.995 ;
			RECT	127.865 31.931 127.897 31.995 ;
			RECT	128.033 31.931 128.065 31.995 ;
			RECT	128.201 31.931 128.233 31.995 ;
			RECT	128.369 31.931 128.401 31.995 ;
			RECT	128.537 31.931 128.569 31.995 ;
			RECT	128.705 31.931 128.737 31.995 ;
			RECT	128.873 31.931 128.905 31.995 ;
			RECT	129.041 31.931 129.073 31.995 ;
			RECT	129.209 31.931 129.241 31.995 ;
			RECT	129.377 31.931 129.409 31.995 ;
			RECT	129.545 31.931 129.577 31.995 ;
			RECT	129.713 31.931 129.745 31.995 ;
			RECT	129.881 31.931 129.913 31.995 ;
			RECT	130.049 31.931 130.081 31.995 ;
			RECT	130.217 31.931 130.249 31.995 ;
			RECT	130.385 31.931 130.417 31.995 ;
			RECT	130.553 31.931 130.585 31.995 ;
			RECT	130.721 31.931 130.753 31.995 ;
			RECT	130.889 31.931 130.921 31.995 ;
			RECT	131.057 31.931 131.089 31.995 ;
			RECT	131.225 31.931 131.257 31.995 ;
			RECT	131.393 31.931 131.425 31.995 ;
			RECT	131.561 31.931 131.593 31.995 ;
			RECT	131.729 31.931 131.761 31.995 ;
			RECT	131.897 31.931 131.929 31.995 ;
			RECT	132.065 31.931 132.097 31.995 ;
			RECT	132.233 31.931 132.265 31.995 ;
			RECT	132.401 31.931 132.433 31.995 ;
			RECT	132.569 31.931 132.601 31.995 ;
			RECT	132.737 31.931 132.769 31.995 ;
			RECT	132.905 31.931 132.937 31.995 ;
			RECT	133.073 31.931 133.105 31.995 ;
			RECT	133.241 31.931 133.273 31.995 ;
			RECT	133.409 31.931 133.441 31.995 ;
			RECT	133.577 31.931 133.609 31.995 ;
			RECT	133.745 31.931 133.777 31.995 ;
			RECT	133.913 31.931 133.945 31.995 ;
			RECT	134.081 31.931 134.113 31.995 ;
			RECT	134.249 31.931 134.281 31.995 ;
			RECT	134.417 31.931 134.449 31.995 ;
			RECT	134.585 31.931 134.617 31.995 ;
			RECT	134.753 31.931 134.785 31.995 ;
			RECT	134.921 31.931 134.953 31.995 ;
			RECT	135.089 31.931 135.121 31.995 ;
			RECT	135.257 31.931 135.289 31.995 ;
			RECT	135.425 31.931 135.457 31.995 ;
			RECT	135.593 31.931 135.625 31.995 ;
			RECT	135.761 31.931 135.793 31.995 ;
			RECT	135.929 31.931 135.961 31.995 ;
			RECT	136.097 31.931 136.129 31.995 ;
			RECT	136.265 31.931 136.297 31.995 ;
			RECT	136.433 31.931 136.465 31.995 ;
			RECT	136.601 31.931 136.633 31.995 ;
			RECT	136.769 31.931 136.801 31.995 ;
			RECT	136.937 31.931 136.969 31.995 ;
			RECT	137.105 31.931 137.137 31.995 ;
			RECT	137.273 31.931 137.305 31.995 ;
			RECT	137.441 31.931 137.473 31.995 ;
			RECT	137.609 31.931 137.641 31.995 ;
			RECT	137.777 31.931 137.809 31.995 ;
			RECT	137.945 31.931 137.977 31.995 ;
			RECT	138.113 31.931 138.145 31.995 ;
			RECT	138.281 31.931 138.313 31.995 ;
			RECT	138.449 31.931 138.481 31.995 ;
			RECT	138.617 31.931 138.649 31.995 ;
			RECT	138.785 31.931 138.817 31.995 ;
			RECT	138.953 31.931 138.985 31.995 ;
			RECT	139.121 31.931 139.153 31.995 ;
			RECT	139.289 31.931 139.321 31.995 ;
			RECT	139.457 31.931 139.489 31.995 ;
			RECT	139.625 31.931 139.657 31.995 ;
			RECT	139.793 31.931 139.825 31.995 ;
			RECT	139.961 31.931 139.993 31.995 ;
			RECT	140.129 31.931 140.161 31.995 ;
			RECT	140.297 31.931 140.329 31.995 ;
			RECT	140.465 31.931 140.497 31.995 ;
			RECT	140.633 31.931 140.665 31.995 ;
			RECT	140.801 31.931 140.833 31.995 ;
			RECT	140.969 31.931 141.001 31.995 ;
			RECT	141.137 31.931 141.169 31.995 ;
			RECT	141.305 31.931 141.337 31.995 ;
			RECT	141.473 31.931 141.505 31.995 ;
			RECT	141.641 31.931 141.673 31.995 ;
			RECT	141.809 31.931 141.841 31.995 ;
			RECT	141.977 31.931 142.009 31.995 ;
			RECT	142.145 31.931 142.177 31.995 ;
			RECT	142.313 31.931 142.345 31.995 ;
			RECT	142.481 31.931 142.513 31.995 ;
			RECT	142.649 31.931 142.681 31.995 ;
			RECT	142.817 31.931 142.849 31.995 ;
			RECT	142.985 31.931 143.017 31.995 ;
			RECT	143.153 31.931 143.185 31.995 ;
			RECT	143.321 31.931 143.353 31.995 ;
			RECT	143.489 31.931 143.521 31.995 ;
			RECT	143.657 31.931 143.689 31.995 ;
			RECT	143.825 31.931 143.857 31.995 ;
			RECT	143.993 31.931 144.025 31.995 ;
			RECT	144.161 31.931 144.193 31.995 ;
			RECT	144.329 31.931 144.361 31.995 ;
			RECT	144.497 31.931 144.529 31.995 ;
			RECT	144.665 31.931 144.697 31.995 ;
			RECT	144.833 31.931 144.865 31.995 ;
			RECT	145.001 31.931 145.033 31.995 ;
			RECT	145.169 31.931 145.201 31.995 ;
			RECT	145.337 31.931 145.369 31.995 ;
			RECT	145.505 31.931 145.537 31.995 ;
			RECT	145.673 31.931 145.705 31.995 ;
			RECT	145.841 31.931 145.873 31.995 ;
			RECT	146.009 31.931 146.041 31.995 ;
			RECT	146.177 31.931 146.209 31.995 ;
			RECT	146.345 31.931 146.377 31.995 ;
			RECT	146.513 31.931 146.545 31.995 ;
			RECT	146.681 31.931 146.713 31.995 ;
			RECT	146.849 31.931 146.881 31.995 ;
			RECT	147.017 31.931 147.049 31.995 ;
			RECT	147.185 31.931 147.217 31.995 ;
			RECT	147.437 31.931 147.469 31.995 ;
			RECT	149.918 31.931 149.95 31.995 ;
			RECT	151.908 31.93 151.94 31.994 ;
			RECT	153.967 31.93 154.031 31.994 ;
			RECT	155.252 31.931 155.284 31.995 ;
			RECT	156.731 31.931 156.763 31.995 ;
			RECT	156.983 31.931 157.015 31.995 ;
			RECT	157.151 31.931 157.183 31.995 ;
			RECT	157.319 31.931 157.351 31.995 ;
			RECT	157.487 31.931 157.519 31.995 ;
			RECT	157.655 31.931 157.687 31.995 ;
			RECT	157.823 31.931 157.855 31.995 ;
			RECT	157.991 31.931 158.023 31.995 ;
			RECT	158.159 31.931 158.191 31.995 ;
			RECT	158.327 31.931 158.359 31.995 ;
			RECT	158.495 31.931 158.527 31.995 ;
			RECT	158.663 31.931 158.695 31.995 ;
			RECT	158.831 31.931 158.863 31.995 ;
			RECT	158.999 31.931 159.031 31.995 ;
			RECT	159.167 31.931 159.199 31.995 ;
			RECT	159.335 31.931 159.367 31.995 ;
			RECT	159.503 31.931 159.535 31.995 ;
			RECT	159.671 31.931 159.703 31.995 ;
			RECT	159.839 31.931 159.871 31.995 ;
			RECT	160.007 31.931 160.039 31.995 ;
			RECT	160.175 31.931 160.207 31.995 ;
			RECT	160.343 31.931 160.375 31.995 ;
			RECT	160.511 31.931 160.543 31.995 ;
			RECT	160.679 31.931 160.711 31.995 ;
			RECT	160.847 31.931 160.879 31.995 ;
			RECT	161.015 31.931 161.047 31.995 ;
			RECT	161.183 31.931 161.215 31.995 ;
			RECT	161.351 31.931 161.383 31.995 ;
			RECT	161.519 31.931 161.551 31.995 ;
			RECT	161.687 31.931 161.719 31.995 ;
			RECT	161.855 31.931 161.887 31.995 ;
			RECT	162.023 31.931 162.055 31.995 ;
			RECT	162.191 31.931 162.223 31.995 ;
			RECT	162.359 31.931 162.391 31.995 ;
			RECT	162.527 31.931 162.559 31.995 ;
			RECT	162.695 31.931 162.727 31.995 ;
			RECT	162.863 31.931 162.895 31.995 ;
			RECT	163.031 31.931 163.063 31.995 ;
			RECT	163.199 31.931 163.231 31.995 ;
			RECT	163.367 31.931 163.399 31.995 ;
			RECT	163.535 31.931 163.567 31.995 ;
			RECT	163.703 31.931 163.735 31.995 ;
			RECT	163.871 31.931 163.903 31.995 ;
			RECT	164.039 31.931 164.071 31.995 ;
			RECT	164.207 31.931 164.239 31.995 ;
			RECT	164.375 31.931 164.407 31.995 ;
			RECT	164.543 31.931 164.575 31.995 ;
			RECT	164.711 31.931 164.743 31.995 ;
			RECT	164.879 31.931 164.911 31.995 ;
			RECT	165.047 31.931 165.079 31.995 ;
			RECT	165.215 31.931 165.247 31.995 ;
			RECT	165.383 31.931 165.415 31.995 ;
			RECT	165.551 31.931 165.583 31.995 ;
			RECT	165.719 31.931 165.751 31.995 ;
			RECT	165.887 31.931 165.919 31.995 ;
			RECT	166.055 31.931 166.087 31.995 ;
			RECT	166.223 31.931 166.255 31.995 ;
			RECT	166.391 31.931 166.423 31.995 ;
			RECT	166.559 31.931 166.591 31.995 ;
			RECT	166.727 31.931 166.759 31.995 ;
			RECT	166.895 31.931 166.927 31.995 ;
			RECT	167.063 31.931 167.095 31.995 ;
			RECT	167.231 31.931 167.263 31.995 ;
			RECT	167.399 31.931 167.431 31.995 ;
			RECT	167.567 31.931 167.599 31.995 ;
			RECT	167.735 31.931 167.767 31.995 ;
			RECT	167.903 31.931 167.935 31.995 ;
			RECT	168.071 31.931 168.103 31.995 ;
			RECT	168.239 31.931 168.271 31.995 ;
			RECT	168.407 31.931 168.439 31.995 ;
			RECT	168.575 31.931 168.607 31.995 ;
			RECT	168.743 31.931 168.775 31.995 ;
			RECT	168.911 31.931 168.943 31.995 ;
			RECT	169.079 31.931 169.111 31.995 ;
			RECT	169.247 31.931 169.279 31.995 ;
			RECT	169.415 31.931 169.447 31.995 ;
			RECT	169.583 31.931 169.615 31.995 ;
			RECT	169.751 31.931 169.783 31.995 ;
			RECT	169.919 31.931 169.951 31.995 ;
			RECT	170.087 31.931 170.119 31.995 ;
			RECT	170.255 31.931 170.287 31.995 ;
			RECT	170.423 31.931 170.455 31.995 ;
			RECT	170.591 31.931 170.623 31.995 ;
			RECT	170.759 31.931 170.791 31.995 ;
			RECT	170.927 31.931 170.959 31.995 ;
			RECT	171.095 31.931 171.127 31.995 ;
			RECT	171.263 31.931 171.295 31.995 ;
			RECT	171.431 31.931 171.463 31.995 ;
			RECT	171.599 31.931 171.631 31.995 ;
			RECT	171.767 31.931 171.799 31.995 ;
			RECT	171.935 31.931 171.967 31.995 ;
			RECT	172.103 31.931 172.135 31.995 ;
			RECT	172.271 31.931 172.303 31.995 ;
			RECT	172.439 31.931 172.471 31.995 ;
			RECT	172.607 31.931 172.639 31.995 ;
			RECT	172.775 31.931 172.807 31.995 ;
			RECT	172.943 31.931 172.975 31.995 ;
			RECT	173.111 31.931 173.143 31.995 ;
			RECT	173.279 31.931 173.311 31.995 ;
			RECT	173.447 31.931 173.479 31.995 ;
			RECT	173.615 31.931 173.647 31.995 ;
			RECT	173.783 31.931 173.815 31.995 ;
			RECT	173.951 31.931 173.983 31.995 ;
			RECT	174.119 31.931 174.151 31.995 ;
			RECT	174.287 31.931 174.319 31.995 ;
			RECT	174.455 31.931 174.487 31.995 ;
			RECT	174.623 31.931 174.655 31.995 ;
			RECT	174.791 31.931 174.823 31.995 ;
			RECT	174.959 31.931 174.991 31.995 ;
			RECT	175.127 31.931 175.159 31.995 ;
			RECT	175.295 31.931 175.327 31.995 ;
			RECT	175.463 31.931 175.495 31.995 ;
			RECT	175.631 31.931 175.663 31.995 ;
			RECT	175.799 31.931 175.831 31.995 ;
			RECT	175.967 31.931 175.999 31.995 ;
			RECT	176.135 31.931 176.167 31.995 ;
			RECT	176.303 31.931 176.335 31.995 ;
			RECT	176.471 31.931 176.503 31.995 ;
			RECT	176.639 31.931 176.671 31.995 ;
			RECT	176.807 31.931 176.839 31.995 ;
			RECT	176.975 31.931 177.007 31.995 ;
			RECT	177.143 31.931 177.175 31.995 ;
			RECT	177.311 31.931 177.343 31.995 ;
			RECT	177.479 31.931 177.511 31.995 ;
			RECT	177.647 31.931 177.679 31.995 ;
			RECT	177.815 31.931 177.847 31.995 ;
			RECT	177.983 31.931 178.015 31.995 ;
			RECT	178.151 31.931 178.183 31.995 ;
			RECT	178.319 31.931 178.351 31.995 ;
			RECT	178.487 31.931 178.519 31.995 ;
			RECT	178.655 31.931 178.687 31.995 ;
			RECT	178.823 31.931 178.855 31.995 ;
			RECT	178.991 31.931 179.023 31.995 ;
			RECT	179.159 31.931 179.191 31.995 ;
			RECT	179.327 31.931 179.359 31.995 ;
			RECT	179.495 31.931 179.527 31.995 ;
			RECT	179.663 31.931 179.695 31.995 ;
			RECT	179.831 31.931 179.863 31.995 ;
			RECT	179.999 31.931 180.031 31.995 ;
			RECT	180.167 31.931 180.199 31.995 ;
			RECT	180.335 31.931 180.367 31.995 ;
			RECT	180.503 31.931 180.535 31.995 ;
			RECT	180.671 31.931 180.703 31.995 ;
			RECT	180.839 31.931 180.871 31.995 ;
			RECT	181.007 31.931 181.039 31.995 ;
			RECT	181.175 31.931 181.207 31.995 ;
			RECT	181.343 31.931 181.375 31.995 ;
			RECT	181.511 31.931 181.543 31.995 ;
			RECT	181.679 31.931 181.711 31.995 ;
			RECT	181.847 31.931 181.879 31.995 ;
			RECT	182.015 31.931 182.047 31.995 ;
			RECT	182.183 31.931 182.215 31.995 ;
			RECT	182.351 31.931 182.383 31.995 ;
			RECT	182.519 31.931 182.551 31.995 ;
			RECT	182.687 31.931 182.719 31.995 ;
			RECT	182.855 31.931 182.887 31.995 ;
			RECT	183.023 31.931 183.055 31.995 ;
			RECT	183.191 31.931 183.223 31.995 ;
			RECT	183.359 31.931 183.391 31.995 ;
			RECT	183.527 31.931 183.559 31.995 ;
			RECT	183.695 31.931 183.727 31.995 ;
			RECT	183.863 31.931 183.895 31.995 ;
			RECT	184.031 31.931 184.063 31.995 ;
			RECT	184.199 31.931 184.231 31.995 ;
			RECT	184.367 31.931 184.399 31.995 ;
			RECT	184.535 31.931 184.567 31.995 ;
			RECT	184.703 31.931 184.735 31.995 ;
			RECT	184.871 31.931 184.903 31.995 ;
			RECT	185.039 31.931 185.071 31.995 ;
			RECT	185.207 31.931 185.239 31.995 ;
			RECT	185.375 31.931 185.407 31.995 ;
			RECT	185.543 31.931 185.575 31.995 ;
			RECT	185.711 31.931 185.743 31.995 ;
			RECT	185.879 31.931 185.911 31.995 ;
			RECT	186.047 31.931 186.079 31.995 ;
			RECT	186.215 31.931 186.247 31.995 ;
			RECT	186.383 31.931 186.415 31.995 ;
			RECT	186.551 31.931 186.583 31.995 ;
			RECT	186.719 31.931 186.751 31.995 ;
			RECT	186.887 31.931 186.919 31.995 ;
			RECT	187.055 31.931 187.087 31.995 ;
			RECT	187.223 31.931 187.255 31.995 ;
			RECT	187.391 31.931 187.423 31.995 ;
			RECT	187.559 31.931 187.591 31.995 ;
			RECT	187.727 31.931 187.759 31.995 ;
			RECT	187.895 31.931 187.927 31.995 ;
			RECT	188.063 31.931 188.095 31.995 ;
			RECT	188.231 31.931 188.263 31.995 ;
			RECT	188.399 31.931 188.431 31.995 ;
			RECT	188.567 31.931 188.599 31.995 ;
			RECT	188.735 31.931 188.767 31.995 ;
			RECT	188.903 31.931 188.935 31.995 ;
			RECT	189.071 31.931 189.103 31.995 ;
			RECT	189.239 31.931 189.271 31.995 ;
			RECT	189.407 31.931 189.439 31.995 ;
			RECT	189.575 31.931 189.607 31.995 ;
			RECT	189.743 31.931 189.775 31.995 ;
			RECT	189.911 31.931 189.943 31.995 ;
			RECT	190.079 31.931 190.111 31.995 ;
			RECT	190.247 31.931 190.279 31.995 ;
			RECT	190.415 31.931 190.447 31.995 ;
			RECT	190.583 31.931 190.615 31.995 ;
			RECT	190.751 31.931 190.783 31.995 ;
			RECT	190.919 31.931 190.951 31.995 ;
			RECT	191.087 31.931 191.119 31.995 ;
			RECT	191.255 31.931 191.287 31.995 ;
			RECT	191.423 31.931 191.455 31.995 ;
			RECT	191.591 31.931 191.623 31.995 ;
			RECT	191.759 31.931 191.791 31.995 ;
			RECT	191.927 31.931 191.959 31.995 ;
			RECT	192.095 31.931 192.127 31.995 ;
			RECT	192.263 31.931 192.295 31.995 ;
			RECT	192.431 31.931 192.463 31.995 ;
			RECT	192.599 31.931 192.631 31.995 ;
			RECT	192.767 31.931 192.799 31.995 ;
			RECT	192.935 31.931 192.967 31.995 ;
			RECT	193.103 31.931 193.135 31.995 ;
			RECT	193.271 31.931 193.303 31.995 ;
			RECT	193.439 31.931 193.471 31.995 ;
			RECT	193.607 31.931 193.639 31.995 ;
			RECT	193.775 31.931 193.807 31.995 ;
			RECT	193.943 31.931 193.975 31.995 ;
			RECT	194.111 31.931 194.143 31.995 ;
			RECT	194.279 31.931 194.311 31.995 ;
			RECT	194.447 31.931 194.479 31.995 ;
			RECT	194.615 31.931 194.647 31.995 ;
			RECT	194.783 31.931 194.815 31.995 ;
			RECT	194.951 31.931 194.983 31.995 ;
			RECT	195.119 31.931 195.151 31.995 ;
			RECT	195.287 31.931 195.319 31.995 ;
			RECT	195.455 31.931 195.487 31.995 ;
			RECT	195.623 31.931 195.655 31.995 ;
			RECT	195.791 31.931 195.823 31.995 ;
			RECT	195.959 31.931 195.991 31.995 ;
			RECT	196.127 31.931 196.159 31.995 ;
			RECT	196.295 31.931 196.327 31.995 ;
			RECT	196.463 31.931 196.495 31.995 ;
			RECT	196.631 31.931 196.663 31.995 ;
			RECT	196.799 31.931 196.831 31.995 ;
			RECT	196.967 31.931 196.999 31.995 ;
			RECT	197.135 31.931 197.167 31.995 ;
			RECT	197.303 31.931 197.335 31.995 ;
			RECT	197.471 31.931 197.503 31.995 ;
			RECT	197.639 31.931 197.671 31.995 ;
			RECT	197.807 31.931 197.839 31.995 ;
			RECT	197.975 31.931 198.007 31.995 ;
			RECT	198.143 31.931 198.175 31.995 ;
			RECT	198.311 31.931 198.343 31.995 ;
			RECT	198.479 31.931 198.511 31.995 ;
			RECT	198.647 31.931 198.679 31.995 ;
			RECT	198.815 31.931 198.847 31.995 ;
			RECT	198.983 31.931 199.015 31.995 ;
			RECT	199.151 31.931 199.183 31.995 ;
			RECT	199.319 31.931 199.351 31.995 ;
			RECT	199.487 31.931 199.519 31.995 ;
			RECT	199.655 31.931 199.687 31.995 ;
			RECT	199.823 31.931 199.855 31.995 ;
			RECT	199.991 31.931 200.023 31.995 ;
			RECT	200.243 31.931 200.275 31.995 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 34.022 201.665 34.142 ;
			LAYER	J3 ;
			RECT	1.645 34.05 1.709 34.114 ;
			RECT	2.124 34.05 2.156 34.114 ;
			RECT	2.323 34.05 2.387 34.114 ;
			RECT	3.438 34.066 3.47 34.098 ;
			RECT	4.195 34.05 4.227 34.114 ;
			RECT	4.354 34.05 4.386 34.114 ;
			RECT	4.96 34.05 4.992 34.114 ;
			RECT	5.252 34.05 5.284 34.114 ;
			RECT	6.179 34.05 6.211 34.114 ;
			RECT	6.347 34.05 6.379 34.114 ;
			RECT	6.515 34.05 6.547 34.114 ;
			RECT	6.683 34.05 6.715 34.114 ;
			RECT	6.851 34.05 6.883 34.114 ;
			RECT	7.019 34.05 7.051 34.114 ;
			RECT	7.187 34.05 7.219 34.114 ;
			RECT	7.355 34.05 7.387 34.114 ;
			RECT	7.523 34.05 7.555 34.114 ;
			RECT	7.691 34.05 7.723 34.114 ;
			RECT	7.859 34.05 7.891 34.114 ;
			RECT	8.027 34.05 8.059 34.114 ;
			RECT	8.195 34.05 8.227 34.114 ;
			RECT	8.363 34.05 8.395 34.114 ;
			RECT	8.531 34.05 8.563 34.114 ;
			RECT	8.699 34.05 8.731 34.114 ;
			RECT	8.867 34.05 8.899 34.114 ;
			RECT	9.035 34.05 9.067 34.114 ;
			RECT	9.203 34.05 9.235 34.114 ;
			RECT	9.371 34.05 9.403 34.114 ;
			RECT	9.539 34.05 9.571 34.114 ;
			RECT	9.707 34.05 9.739 34.114 ;
			RECT	9.875 34.05 9.907 34.114 ;
			RECT	10.043 34.05 10.075 34.114 ;
			RECT	10.211 34.05 10.243 34.114 ;
			RECT	10.379 34.05 10.411 34.114 ;
			RECT	10.547 34.05 10.579 34.114 ;
			RECT	10.715 34.05 10.747 34.114 ;
			RECT	10.883 34.05 10.915 34.114 ;
			RECT	11.051 34.05 11.083 34.114 ;
			RECT	11.219 34.05 11.251 34.114 ;
			RECT	11.387 34.05 11.419 34.114 ;
			RECT	11.555 34.05 11.587 34.114 ;
			RECT	11.723 34.05 11.755 34.114 ;
			RECT	11.891 34.05 11.923 34.114 ;
			RECT	12.059 34.05 12.091 34.114 ;
			RECT	12.227 34.05 12.259 34.114 ;
			RECT	12.395 34.05 12.427 34.114 ;
			RECT	12.563 34.05 12.595 34.114 ;
			RECT	12.731 34.05 12.763 34.114 ;
			RECT	12.899 34.05 12.931 34.114 ;
			RECT	13.067 34.05 13.099 34.114 ;
			RECT	13.235 34.05 13.267 34.114 ;
			RECT	13.403 34.05 13.435 34.114 ;
			RECT	13.571 34.05 13.603 34.114 ;
			RECT	13.739 34.05 13.771 34.114 ;
			RECT	13.907 34.05 13.939 34.114 ;
			RECT	14.075 34.05 14.107 34.114 ;
			RECT	14.243 34.05 14.275 34.114 ;
			RECT	14.411 34.05 14.443 34.114 ;
			RECT	14.579 34.05 14.611 34.114 ;
			RECT	14.747 34.05 14.779 34.114 ;
			RECT	14.915 34.05 14.947 34.114 ;
			RECT	15.083 34.05 15.115 34.114 ;
			RECT	15.251 34.05 15.283 34.114 ;
			RECT	15.419 34.05 15.451 34.114 ;
			RECT	15.587 34.05 15.619 34.114 ;
			RECT	15.755 34.05 15.787 34.114 ;
			RECT	15.923 34.05 15.955 34.114 ;
			RECT	16.091 34.05 16.123 34.114 ;
			RECT	16.259 34.05 16.291 34.114 ;
			RECT	16.427 34.05 16.459 34.114 ;
			RECT	16.595 34.05 16.627 34.114 ;
			RECT	16.763 34.05 16.795 34.114 ;
			RECT	16.931 34.05 16.963 34.114 ;
			RECT	17.099 34.05 17.131 34.114 ;
			RECT	17.267 34.05 17.299 34.114 ;
			RECT	17.435 34.05 17.467 34.114 ;
			RECT	17.603 34.05 17.635 34.114 ;
			RECT	17.771 34.05 17.803 34.114 ;
			RECT	17.939 34.05 17.971 34.114 ;
			RECT	18.107 34.05 18.139 34.114 ;
			RECT	18.275 34.05 18.307 34.114 ;
			RECT	18.443 34.05 18.475 34.114 ;
			RECT	18.611 34.05 18.643 34.114 ;
			RECT	18.779 34.05 18.811 34.114 ;
			RECT	18.947 34.05 18.979 34.114 ;
			RECT	19.115 34.05 19.147 34.114 ;
			RECT	19.283 34.05 19.315 34.114 ;
			RECT	19.451 34.05 19.483 34.114 ;
			RECT	19.619 34.05 19.651 34.114 ;
			RECT	19.787 34.05 19.819 34.114 ;
			RECT	19.955 34.05 19.987 34.114 ;
			RECT	20.123 34.05 20.155 34.114 ;
			RECT	20.291 34.05 20.323 34.114 ;
			RECT	20.459 34.05 20.491 34.114 ;
			RECT	20.627 34.05 20.659 34.114 ;
			RECT	20.795 34.05 20.827 34.114 ;
			RECT	20.963 34.05 20.995 34.114 ;
			RECT	21.131 34.05 21.163 34.114 ;
			RECT	21.299 34.05 21.331 34.114 ;
			RECT	21.467 34.05 21.499 34.114 ;
			RECT	21.635 34.05 21.667 34.114 ;
			RECT	21.803 34.05 21.835 34.114 ;
			RECT	21.971 34.05 22.003 34.114 ;
			RECT	22.139 34.05 22.171 34.114 ;
			RECT	22.307 34.05 22.339 34.114 ;
			RECT	22.475 34.05 22.507 34.114 ;
			RECT	22.643 34.05 22.675 34.114 ;
			RECT	22.811 34.05 22.843 34.114 ;
			RECT	22.979 34.05 23.011 34.114 ;
			RECT	23.147 34.05 23.179 34.114 ;
			RECT	23.315 34.05 23.347 34.114 ;
			RECT	23.483 34.05 23.515 34.114 ;
			RECT	23.651 34.05 23.683 34.114 ;
			RECT	23.819 34.05 23.851 34.114 ;
			RECT	23.987 34.05 24.019 34.114 ;
			RECT	24.155 34.05 24.187 34.114 ;
			RECT	24.323 34.05 24.355 34.114 ;
			RECT	24.491 34.05 24.523 34.114 ;
			RECT	24.659 34.05 24.691 34.114 ;
			RECT	24.827 34.05 24.859 34.114 ;
			RECT	24.995 34.05 25.027 34.114 ;
			RECT	25.163 34.05 25.195 34.114 ;
			RECT	25.331 34.05 25.363 34.114 ;
			RECT	25.499 34.05 25.531 34.114 ;
			RECT	25.667 34.05 25.699 34.114 ;
			RECT	25.835 34.05 25.867 34.114 ;
			RECT	26.003 34.05 26.035 34.114 ;
			RECT	26.171 34.05 26.203 34.114 ;
			RECT	26.339 34.05 26.371 34.114 ;
			RECT	26.507 34.05 26.539 34.114 ;
			RECT	26.675 34.05 26.707 34.114 ;
			RECT	26.843 34.05 26.875 34.114 ;
			RECT	27.011 34.05 27.043 34.114 ;
			RECT	27.179 34.05 27.211 34.114 ;
			RECT	27.347 34.05 27.379 34.114 ;
			RECT	27.515 34.05 27.547 34.114 ;
			RECT	27.683 34.05 27.715 34.114 ;
			RECT	27.851 34.05 27.883 34.114 ;
			RECT	28.019 34.05 28.051 34.114 ;
			RECT	28.187 34.05 28.219 34.114 ;
			RECT	28.355 34.05 28.387 34.114 ;
			RECT	28.523 34.05 28.555 34.114 ;
			RECT	28.691 34.05 28.723 34.114 ;
			RECT	28.859 34.05 28.891 34.114 ;
			RECT	29.027 34.05 29.059 34.114 ;
			RECT	29.195 34.05 29.227 34.114 ;
			RECT	29.363 34.05 29.395 34.114 ;
			RECT	29.531 34.05 29.563 34.114 ;
			RECT	29.699 34.05 29.731 34.114 ;
			RECT	29.867 34.05 29.899 34.114 ;
			RECT	30.035 34.05 30.067 34.114 ;
			RECT	30.203 34.05 30.235 34.114 ;
			RECT	30.371 34.05 30.403 34.114 ;
			RECT	30.539 34.05 30.571 34.114 ;
			RECT	30.707 34.05 30.739 34.114 ;
			RECT	30.875 34.05 30.907 34.114 ;
			RECT	31.043 34.05 31.075 34.114 ;
			RECT	31.211 34.05 31.243 34.114 ;
			RECT	31.379 34.05 31.411 34.114 ;
			RECT	31.547 34.05 31.579 34.114 ;
			RECT	31.715 34.05 31.747 34.114 ;
			RECT	31.883 34.05 31.915 34.114 ;
			RECT	32.051 34.05 32.083 34.114 ;
			RECT	32.219 34.05 32.251 34.114 ;
			RECT	32.387 34.05 32.419 34.114 ;
			RECT	32.555 34.05 32.587 34.114 ;
			RECT	32.723 34.05 32.755 34.114 ;
			RECT	32.891 34.05 32.923 34.114 ;
			RECT	33.059 34.05 33.091 34.114 ;
			RECT	33.227 34.05 33.259 34.114 ;
			RECT	33.395 34.05 33.427 34.114 ;
			RECT	33.563 34.05 33.595 34.114 ;
			RECT	33.731 34.05 33.763 34.114 ;
			RECT	33.899 34.05 33.931 34.114 ;
			RECT	34.067 34.05 34.099 34.114 ;
			RECT	34.235 34.05 34.267 34.114 ;
			RECT	34.403 34.05 34.435 34.114 ;
			RECT	34.571 34.05 34.603 34.114 ;
			RECT	34.739 34.05 34.771 34.114 ;
			RECT	34.907 34.05 34.939 34.114 ;
			RECT	35.075 34.05 35.107 34.114 ;
			RECT	35.243 34.05 35.275 34.114 ;
			RECT	35.411 34.05 35.443 34.114 ;
			RECT	35.579 34.05 35.611 34.114 ;
			RECT	35.747 34.05 35.779 34.114 ;
			RECT	35.915 34.05 35.947 34.114 ;
			RECT	36.083 34.05 36.115 34.114 ;
			RECT	36.251 34.05 36.283 34.114 ;
			RECT	36.419 34.05 36.451 34.114 ;
			RECT	36.587 34.05 36.619 34.114 ;
			RECT	36.755 34.05 36.787 34.114 ;
			RECT	36.923 34.05 36.955 34.114 ;
			RECT	37.091 34.05 37.123 34.114 ;
			RECT	37.259 34.05 37.291 34.114 ;
			RECT	37.427 34.05 37.459 34.114 ;
			RECT	37.595 34.05 37.627 34.114 ;
			RECT	37.763 34.05 37.795 34.114 ;
			RECT	37.931 34.05 37.963 34.114 ;
			RECT	38.099 34.05 38.131 34.114 ;
			RECT	38.267 34.05 38.299 34.114 ;
			RECT	38.435 34.05 38.467 34.114 ;
			RECT	38.603 34.05 38.635 34.114 ;
			RECT	38.771 34.05 38.803 34.114 ;
			RECT	38.939 34.05 38.971 34.114 ;
			RECT	39.107 34.05 39.139 34.114 ;
			RECT	39.275 34.05 39.307 34.114 ;
			RECT	39.443 34.05 39.475 34.114 ;
			RECT	39.611 34.05 39.643 34.114 ;
			RECT	39.779 34.05 39.811 34.114 ;
			RECT	39.947 34.05 39.979 34.114 ;
			RECT	40.115 34.05 40.147 34.114 ;
			RECT	40.283 34.05 40.315 34.114 ;
			RECT	40.451 34.05 40.483 34.114 ;
			RECT	40.619 34.05 40.651 34.114 ;
			RECT	40.787 34.05 40.819 34.114 ;
			RECT	40.955 34.05 40.987 34.114 ;
			RECT	41.123 34.05 41.155 34.114 ;
			RECT	41.291 34.05 41.323 34.114 ;
			RECT	41.459 34.05 41.491 34.114 ;
			RECT	41.627 34.05 41.659 34.114 ;
			RECT	41.795 34.05 41.827 34.114 ;
			RECT	41.963 34.05 41.995 34.114 ;
			RECT	42.131 34.05 42.163 34.114 ;
			RECT	42.299 34.05 42.331 34.114 ;
			RECT	42.467 34.05 42.499 34.114 ;
			RECT	42.635 34.05 42.667 34.114 ;
			RECT	42.803 34.05 42.835 34.114 ;
			RECT	42.971 34.05 43.003 34.114 ;
			RECT	43.139 34.05 43.171 34.114 ;
			RECT	43.307 34.05 43.339 34.114 ;
			RECT	43.475 34.05 43.507 34.114 ;
			RECT	43.643 34.05 43.675 34.114 ;
			RECT	43.811 34.05 43.843 34.114 ;
			RECT	43.979 34.05 44.011 34.114 ;
			RECT	44.147 34.05 44.179 34.114 ;
			RECT	44.315 34.05 44.347 34.114 ;
			RECT	44.483 34.05 44.515 34.114 ;
			RECT	44.651 34.05 44.683 34.114 ;
			RECT	44.819 34.05 44.851 34.114 ;
			RECT	44.987 34.05 45.019 34.114 ;
			RECT	45.155 34.05 45.187 34.114 ;
			RECT	45.323 34.05 45.355 34.114 ;
			RECT	45.491 34.05 45.523 34.114 ;
			RECT	45.659 34.05 45.691 34.114 ;
			RECT	45.827 34.05 45.859 34.114 ;
			RECT	45.995 34.05 46.027 34.114 ;
			RECT	46.163 34.05 46.195 34.114 ;
			RECT	46.331 34.05 46.363 34.114 ;
			RECT	46.499 34.05 46.531 34.114 ;
			RECT	46.667 34.05 46.699 34.114 ;
			RECT	46.835 34.05 46.867 34.114 ;
			RECT	47.003 34.05 47.035 34.114 ;
			RECT	47.171 34.05 47.203 34.114 ;
			RECT	47.339 34.05 47.371 34.114 ;
			RECT	47.507 34.05 47.539 34.114 ;
			RECT	47.675 34.05 47.707 34.114 ;
			RECT	47.843 34.05 47.875 34.114 ;
			RECT	48.011 34.05 48.043 34.114 ;
			RECT	48.179 34.05 48.211 34.114 ;
			RECT	48.347 34.05 48.379 34.114 ;
			RECT	48.515 34.05 48.547 34.114 ;
			RECT	48.683 34.05 48.715 34.114 ;
			RECT	48.851 34.05 48.883 34.114 ;
			RECT	49.019 34.05 49.051 34.114 ;
			RECT	49.187 34.05 49.219 34.114 ;
			RECT	49.311 34.05 49.375 34.114 ;
			RECT	49.613 34.05 49.645 34.114 ;
			RECT	49.813 34.05 49.845 34.114 ;
			RECT	51.92 34.05 51.952 34.114 ;
			RECT	52.578 34.05 52.61 34.114 ;
			RECT	53.91 34.05 53.942 34.114 ;
			RECT	55.466 34.05 55.498 34.114 ;
			RECT	55.803 34.05 55.835 34.114 ;
			RECT	55.969 34.05 56.033 34.114 ;
			RECT	58.359 34.05 58.391 34.114 ;
			RECT	58.559 34.05 58.591 34.114 ;
			RECT	58.829 34.05 58.893 34.114 ;
			RECT	58.985 34.05 59.017 34.114 ;
			RECT	59.153 34.05 59.185 34.114 ;
			RECT	59.321 34.05 59.353 34.114 ;
			RECT	59.489 34.05 59.521 34.114 ;
			RECT	59.657 34.05 59.689 34.114 ;
			RECT	59.825 34.05 59.857 34.114 ;
			RECT	59.993 34.05 60.025 34.114 ;
			RECT	60.161 34.05 60.193 34.114 ;
			RECT	60.329 34.05 60.361 34.114 ;
			RECT	60.497 34.05 60.529 34.114 ;
			RECT	60.665 34.05 60.697 34.114 ;
			RECT	60.833 34.05 60.865 34.114 ;
			RECT	61.001 34.05 61.033 34.114 ;
			RECT	61.169 34.05 61.201 34.114 ;
			RECT	61.337 34.05 61.369 34.114 ;
			RECT	61.505 34.05 61.537 34.114 ;
			RECT	61.673 34.05 61.705 34.114 ;
			RECT	61.841 34.05 61.873 34.114 ;
			RECT	62.009 34.05 62.041 34.114 ;
			RECT	62.177 34.05 62.209 34.114 ;
			RECT	62.345 34.05 62.377 34.114 ;
			RECT	62.513 34.05 62.545 34.114 ;
			RECT	62.681 34.05 62.713 34.114 ;
			RECT	62.849 34.05 62.881 34.114 ;
			RECT	63.017 34.05 63.049 34.114 ;
			RECT	63.185 34.05 63.217 34.114 ;
			RECT	63.353 34.05 63.385 34.114 ;
			RECT	63.521 34.05 63.553 34.114 ;
			RECT	63.689 34.05 63.721 34.114 ;
			RECT	63.857 34.05 63.889 34.114 ;
			RECT	64.025 34.05 64.057 34.114 ;
			RECT	64.193 34.05 64.225 34.114 ;
			RECT	64.361 34.05 64.393 34.114 ;
			RECT	64.529 34.05 64.561 34.114 ;
			RECT	64.697 34.05 64.729 34.114 ;
			RECT	64.865 34.05 64.897 34.114 ;
			RECT	65.033 34.05 65.065 34.114 ;
			RECT	65.201 34.05 65.233 34.114 ;
			RECT	65.369 34.05 65.401 34.114 ;
			RECT	65.537 34.05 65.569 34.114 ;
			RECT	65.705 34.05 65.737 34.114 ;
			RECT	65.873 34.05 65.905 34.114 ;
			RECT	66.041 34.05 66.073 34.114 ;
			RECT	66.209 34.05 66.241 34.114 ;
			RECT	66.377 34.05 66.409 34.114 ;
			RECT	66.545 34.05 66.577 34.114 ;
			RECT	66.713 34.05 66.745 34.114 ;
			RECT	66.881 34.05 66.913 34.114 ;
			RECT	67.049 34.05 67.081 34.114 ;
			RECT	67.217 34.05 67.249 34.114 ;
			RECT	67.385 34.05 67.417 34.114 ;
			RECT	67.553 34.05 67.585 34.114 ;
			RECT	67.721 34.05 67.753 34.114 ;
			RECT	67.889 34.05 67.921 34.114 ;
			RECT	68.057 34.05 68.089 34.114 ;
			RECT	68.225 34.05 68.257 34.114 ;
			RECT	68.393 34.05 68.425 34.114 ;
			RECT	68.561 34.05 68.593 34.114 ;
			RECT	68.729 34.05 68.761 34.114 ;
			RECT	68.897 34.05 68.929 34.114 ;
			RECT	69.065 34.05 69.097 34.114 ;
			RECT	69.233 34.05 69.265 34.114 ;
			RECT	69.401 34.05 69.433 34.114 ;
			RECT	69.569 34.05 69.601 34.114 ;
			RECT	69.737 34.05 69.769 34.114 ;
			RECT	69.905 34.05 69.937 34.114 ;
			RECT	70.073 34.05 70.105 34.114 ;
			RECT	70.241 34.05 70.273 34.114 ;
			RECT	70.409 34.05 70.441 34.114 ;
			RECT	70.577 34.05 70.609 34.114 ;
			RECT	70.745 34.05 70.777 34.114 ;
			RECT	70.913 34.05 70.945 34.114 ;
			RECT	71.081 34.05 71.113 34.114 ;
			RECT	71.249 34.05 71.281 34.114 ;
			RECT	71.417 34.05 71.449 34.114 ;
			RECT	71.585 34.05 71.617 34.114 ;
			RECT	71.753 34.05 71.785 34.114 ;
			RECT	71.921 34.05 71.953 34.114 ;
			RECT	72.089 34.05 72.121 34.114 ;
			RECT	72.257 34.05 72.289 34.114 ;
			RECT	72.425 34.05 72.457 34.114 ;
			RECT	72.593 34.05 72.625 34.114 ;
			RECT	72.761 34.05 72.793 34.114 ;
			RECT	72.929 34.05 72.961 34.114 ;
			RECT	73.097 34.05 73.129 34.114 ;
			RECT	73.265 34.05 73.297 34.114 ;
			RECT	73.433 34.05 73.465 34.114 ;
			RECT	73.601 34.05 73.633 34.114 ;
			RECT	73.769 34.05 73.801 34.114 ;
			RECT	73.937 34.05 73.969 34.114 ;
			RECT	74.105 34.05 74.137 34.114 ;
			RECT	74.273 34.05 74.305 34.114 ;
			RECT	74.441 34.05 74.473 34.114 ;
			RECT	74.609 34.05 74.641 34.114 ;
			RECT	74.777 34.05 74.809 34.114 ;
			RECT	74.945 34.05 74.977 34.114 ;
			RECT	75.113 34.05 75.145 34.114 ;
			RECT	75.281 34.05 75.313 34.114 ;
			RECT	75.449 34.05 75.481 34.114 ;
			RECT	75.617 34.05 75.649 34.114 ;
			RECT	75.785 34.05 75.817 34.114 ;
			RECT	75.953 34.05 75.985 34.114 ;
			RECT	76.121 34.05 76.153 34.114 ;
			RECT	76.289 34.05 76.321 34.114 ;
			RECT	76.457 34.05 76.489 34.114 ;
			RECT	76.625 34.05 76.657 34.114 ;
			RECT	76.793 34.05 76.825 34.114 ;
			RECT	76.961 34.05 76.993 34.114 ;
			RECT	77.129 34.05 77.161 34.114 ;
			RECT	77.297 34.05 77.329 34.114 ;
			RECT	77.465 34.05 77.497 34.114 ;
			RECT	77.633 34.05 77.665 34.114 ;
			RECT	77.801 34.05 77.833 34.114 ;
			RECT	77.969 34.05 78.001 34.114 ;
			RECT	78.137 34.05 78.169 34.114 ;
			RECT	78.305 34.05 78.337 34.114 ;
			RECT	78.473 34.05 78.505 34.114 ;
			RECT	78.641 34.05 78.673 34.114 ;
			RECT	78.809 34.05 78.841 34.114 ;
			RECT	78.977 34.05 79.009 34.114 ;
			RECT	79.145 34.05 79.177 34.114 ;
			RECT	79.313 34.05 79.345 34.114 ;
			RECT	79.481 34.05 79.513 34.114 ;
			RECT	79.649 34.05 79.681 34.114 ;
			RECT	79.817 34.05 79.849 34.114 ;
			RECT	79.985 34.05 80.017 34.114 ;
			RECT	80.153 34.05 80.185 34.114 ;
			RECT	80.321 34.05 80.353 34.114 ;
			RECT	80.489 34.05 80.521 34.114 ;
			RECT	80.657 34.05 80.689 34.114 ;
			RECT	80.825 34.05 80.857 34.114 ;
			RECT	80.993 34.05 81.025 34.114 ;
			RECT	81.161 34.05 81.193 34.114 ;
			RECT	81.329 34.05 81.361 34.114 ;
			RECT	81.497 34.05 81.529 34.114 ;
			RECT	81.665 34.05 81.697 34.114 ;
			RECT	81.833 34.05 81.865 34.114 ;
			RECT	82.001 34.05 82.033 34.114 ;
			RECT	82.169 34.05 82.201 34.114 ;
			RECT	82.337 34.05 82.369 34.114 ;
			RECT	82.505 34.05 82.537 34.114 ;
			RECT	82.673 34.05 82.705 34.114 ;
			RECT	82.841 34.05 82.873 34.114 ;
			RECT	83.009 34.05 83.041 34.114 ;
			RECT	83.177 34.05 83.209 34.114 ;
			RECT	83.345 34.05 83.377 34.114 ;
			RECT	83.513 34.05 83.545 34.114 ;
			RECT	83.681 34.05 83.713 34.114 ;
			RECT	83.849 34.05 83.881 34.114 ;
			RECT	84.017 34.05 84.049 34.114 ;
			RECT	84.185 34.05 84.217 34.114 ;
			RECT	84.353 34.05 84.385 34.114 ;
			RECT	84.521 34.05 84.553 34.114 ;
			RECT	84.689 34.05 84.721 34.114 ;
			RECT	84.857 34.05 84.889 34.114 ;
			RECT	85.025 34.05 85.057 34.114 ;
			RECT	85.193 34.05 85.225 34.114 ;
			RECT	85.361 34.05 85.393 34.114 ;
			RECT	85.529 34.05 85.561 34.114 ;
			RECT	85.697 34.05 85.729 34.114 ;
			RECT	85.865 34.05 85.897 34.114 ;
			RECT	86.033 34.05 86.065 34.114 ;
			RECT	86.201 34.05 86.233 34.114 ;
			RECT	86.369 34.05 86.401 34.114 ;
			RECT	86.537 34.05 86.569 34.114 ;
			RECT	86.705 34.05 86.737 34.114 ;
			RECT	86.873 34.05 86.905 34.114 ;
			RECT	87.041 34.05 87.073 34.114 ;
			RECT	87.209 34.05 87.241 34.114 ;
			RECT	87.377 34.05 87.409 34.114 ;
			RECT	87.545 34.05 87.577 34.114 ;
			RECT	87.713 34.05 87.745 34.114 ;
			RECT	87.881 34.05 87.913 34.114 ;
			RECT	88.049 34.05 88.081 34.114 ;
			RECT	88.217 34.05 88.249 34.114 ;
			RECT	88.385 34.05 88.417 34.114 ;
			RECT	88.553 34.05 88.585 34.114 ;
			RECT	88.721 34.05 88.753 34.114 ;
			RECT	88.889 34.05 88.921 34.114 ;
			RECT	89.057 34.05 89.089 34.114 ;
			RECT	89.225 34.05 89.257 34.114 ;
			RECT	89.393 34.05 89.425 34.114 ;
			RECT	89.561 34.05 89.593 34.114 ;
			RECT	89.729 34.05 89.761 34.114 ;
			RECT	89.897 34.05 89.929 34.114 ;
			RECT	90.065 34.05 90.097 34.114 ;
			RECT	90.233 34.05 90.265 34.114 ;
			RECT	90.401 34.05 90.433 34.114 ;
			RECT	90.569 34.05 90.601 34.114 ;
			RECT	90.737 34.05 90.769 34.114 ;
			RECT	90.905 34.05 90.937 34.114 ;
			RECT	91.073 34.05 91.105 34.114 ;
			RECT	91.241 34.05 91.273 34.114 ;
			RECT	91.409 34.05 91.441 34.114 ;
			RECT	91.577 34.05 91.609 34.114 ;
			RECT	91.745 34.05 91.777 34.114 ;
			RECT	91.913 34.05 91.945 34.114 ;
			RECT	92.081 34.05 92.113 34.114 ;
			RECT	92.249 34.05 92.281 34.114 ;
			RECT	92.417 34.05 92.449 34.114 ;
			RECT	92.585 34.05 92.617 34.114 ;
			RECT	92.753 34.05 92.785 34.114 ;
			RECT	92.921 34.05 92.953 34.114 ;
			RECT	93.089 34.05 93.121 34.114 ;
			RECT	93.257 34.05 93.289 34.114 ;
			RECT	93.425 34.05 93.457 34.114 ;
			RECT	93.593 34.05 93.625 34.114 ;
			RECT	93.761 34.05 93.793 34.114 ;
			RECT	93.929 34.05 93.961 34.114 ;
			RECT	94.097 34.05 94.129 34.114 ;
			RECT	94.265 34.05 94.297 34.114 ;
			RECT	94.433 34.05 94.465 34.114 ;
			RECT	94.601 34.05 94.633 34.114 ;
			RECT	94.769 34.05 94.801 34.114 ;
			RECT	94.937 34.05 94.969 34.114 ;
			RECT	95.105 34.05 95.137 34.114 ;
			RECT	95.273 34.05 95.305 34.114 ;
			RECT	95.441 34.05 95.473 34.114 ;
			RECT	95.609 34.05 95.641 34.114 ;
			RECT	95.777 34.05 95.809 34.114 ;
			RECT	95.945 34.05 95.977 34.114 ;
			RECT	96.113 34.05 96.145 34.114 ;
			RECT	96.281 34.05 96.313 34.114 ;
			RECT	96.449 34.05 96.481 34.114 ;
			RECT	96.617 34.05 96.649 34.114 ;
			RECT	96.785 34.05 96.817 34.114 ;
			RECT	96.953 34.05 96.985 34.114 ;
			RECT	97.121 34.05 97.153 34.114 ;
			RECT	97.289 34.05 97.321 34.114 ;
			RECT	97.457 34.05 97.489 34.114 ;
			RECT	97.625 34.05 97.657 34.114 ;
			RECT	97.793 34.05 97.825 34.114 ;
			RECT	97.961 34.05 97.993 34.114 ;
			RECT	98.129 34.05 98.161 34.114 ;
			RECT	98.297 34.05 98.329 34.114 ;
			RECT	98.465 34.05 98.497 34.114 ;
			RECT	98.633 34.05 98.665 34.114 ;
			RECT	98.801 34.05 98.833 34.114 ;
			RECT	98.969 34.05 99.001 34.114 ;
			RECT	99.137 34.05 99.169 34.114 ;
			RECT	99.305 34.05 99.337 34.114 ;
			RECT	99.473 34.05 99.505 34.114 ;
			RECT	99.641 34.05 99.673 34.114 ;
			RECT	99.809 34.05 99.841 34.114 ;
			RECT	99.977 34.05 100.009 34.114 ;
			RECT	100.145 34.05 100.177 34.114 ;
			RECT	100.313 34.05 100.345 34.114 ;
			RECT	100.481 34.05 100.513 34.114 ;
			RECT	100.649 34.05 100.681 34.114 ;
			RECT	100.817 34.05 100.849 34.114 ;
			RECT	100.985 34.05 101.017 34.114 ;
			RECT	101.153 34.05 101.185 34.114 ;
			RECT	101.321 34.05 101.353 34.114 ;
			RECT	101.489 34.05 101.521 34.114 ;
			RECT	101.657 34.05 101.689 34.114 ;
			RECT	101.825 34.05 101.857 34.114 ;
			RECT	101.993 34.05 102.025 34.114 ;
			RECT	104.177 34.05 104.209 34.114 ;
			RECT	104.345 34.05 104.377 34.114 ;
			RECT	104.513 34.05 104.545 34.114 ;
			RECT	104.681 34.05 104.713 34.114 ;
			RECT	104.849 34.05 104.881 34.114 ;
			RECT	105.017 34.05 105.049 34.114 ;
			RECT	105.185 34.05 105.217 34.114 ;
			RECT	105.353 34.05 105.385 34.114 ;
			RECT	105.521 34.05 105.553 34.114 ;
			RECT	105.689 34.05 105.721 34.114 ;
			RECT	105.857 34.05 105.889 34.114 ;
			RECT	106.025 34.05 106.057 34.114 ;
			RECT	106.193 34.05 106.225 34.114 ;
			RECT	106.361 34.05 106.393 34.114 ;
			RECT	106.529 34.05 106.561 34.114 ;
			RECT	106.697 34.05 106.729 34.114 ;
			RECT	106.865 34.05 106.897 34.114 ;
			RECT	107.033 34.05 107.065 34.114 ;
			RECT	107.201 34.05 107.233 34.114 ;
			RECT	107.369 34.05 107.401 34.114 ;
			RECT	107.537 34.05 107.569 34.114 ;
			RECT	107.705 34.05 107.737 34.114 ;
			RECT	107.873 34.05 107.905 34.114 ;
			RECT	108.041 34.05 108.073 34.114 ;
			RECT	108.209 34.05 108.241 34.114 ;
			RECT	108.377 34.05 108.409 34.114 ;
			RECT	108.545 34.05 108.577 34.114 ;
			RECT	108.713 34.05 108.745 34.114 ;
			RECT	108.881 34.05 108.913 34.114 ;
			RECT	109.049 34.05 109.081 34.114 ;
			RECT	109.217 34.05 109.249 34.114 ;
			RECT	109.385 34.05 109.417 34.114 ;
			RECT	109.553 34.05 109.585 34.114 ;
			RECT	109.721 34.05 109.753 34.114 ;
			RECT	109.889 34.05 109.921 34.114 ;
			RECT	110.057 34.05 110.089 34.114 ;
			RECT	110.225 34.05 110.257 34.114 ;
			RECT	110.393 34.05 110.425 34.114 ;
			RECT	110.561 34.05 110.593 34.114 ;
			RECT	110.729 34.05 110.761 34.114 ;
			RECT	110.897 34.05 110.929 34.114 ;
			RECT	111.065 34.05 111.097 34.114 ;
			RECT	111.233 34.05 111.265 34.114 ;
			RECT	111.401 34.05 111.433 34.114 ;
			RECT	111.569 34.05 111.601 34.114 ;
			RECT	111.737 34.05 111.769 34.114 ;
			RECT	111.905 34.05 111.937 34.114 ;
			RECT	112.073 34.05 112.105 34.114 ;
			RECT	112.241 34.05 112.273 34.114 ;
			RECT	112.409 34.05 112.441 34.114 ;
			RECT	112.577 34.05 112.609 34.114 ;
			RECT	112.745 34.05 112.777 34.114 ;
			RECT	112.913 34.05 112.945 34.114 ;
			RECT	113.081 34.05 113.113 34.114 ;
			RECT	113.249 34.05 113.281 34.114 ;
			RECT	113.417 34.05 113.449 34.114 ;
			RECT	113.585 34.05 113.617 34.114 ;
			RECT	113.753 34.05 113.785 34.114 ;
			RECT	113.921 34.05 113.953 34.114 ;
			RECT	114.089 34.05 114.121 34.114 ;
			RECT	114.257 34.05 114.289 34.114 ;
			RECT	114.425 34.05 114.457 34.114 ;
			RECT	114.593 34.05 114.625 34.114 ;
			RECT	114.761 34.05 114.793 34.114 ;
			RECT	114.929 34.05 114.961 34.114 ;
			RECT	115.097 34.05 115.129 34.114 ;
			RECT	115.265 34.05 115.297 34.114 ;
			RECT	115.433 34.05 115.465 34.114 ;
			RECT	115.601 34.05 115.633 34.114 ;
			RECT	115.769 34.05 115.801 34.114 ;
			RECT	115.937 34.05 115.969 34.114 ;
			RECT	116.105 34.05 116.137 34.114 ;
			RECT	116.273 34.05 116.305 34.114 ;
			RECT	116.441 34.05 116.473 34.114 ;
			RECT	116.609 34.05 116.641 34.114 ;
			RECT	116.777 34.05 116.809 34.114 ;
			RECT	116.945 34.05 116.977 34.114 ;
			RECT	117.113 34.05 117.145 34.114 ;
			RECT	117.281 34.05 117.313 34.114 ;
			RECT	117.449 34.05 117.481 34.114 ;
			RECT	117.617 34.05 117.649 34.114 ;
			RECT	117.785 34.05 117.817 34.114 ;
			RECT	117.953 34.05 117.985 34.114 ;
			RECT	118.121 34.05 118.153 34.114 ;
			RECT	118.289 34.05 118.321 34.114 ;
			RECT	118.457 34.05 118.489 34.114 ;
			RECT	118.625 34.05 118.657 34.114 ;
			RECT	118.793 34.05 118.825 34.114 ;
			RECT	118.961 34.05 118.993 34.114 ;
			RECT	119.129 34.05 119.161 34.114 ;
			RECT	119.297 34.05 119.329 34.114 ;
			RECT	119.465 34.05 119.497 34.114 ;
			RECT	119.633 34.05 119.665 34.114 ;
			RECT	119.801 34.05 119.833 34.114 ;
			RECT	119.969 34.05 120.001 34.114 ;
			RECT	120.137 34.05 120.169 34.114 ;
			RECT	120.305 34.05 120.337 34.114 ;
			RECT	120.473 34.05 120.505 34.114 ;
			RECT	120.641 34.05 120.673 34.114 ;
			RECT	120.809 34.05 120.841 34.114 ;
			RECT	120.977 34.05 121.009 34.114 ;
			RECT	121.145 34.05 121.177 34.114 ;
			RECT	121.313 34.05 121.345 34.114 ;
			RECT	121.481 34.05 121.513 34.114 ;
			RECT	121.649 34.05 121.681 34.114 ;
			RECT	121.817 34.05 121.849 34.114 ;
			RECT	121.985 34.05 122.017 34.114 ;
			RECT	122.153 34.05 122.185 34.114 ;
			RECT	122.321 34.05 122.353 34.114 ;
			RECT	122.489 34.05 122.521 34.114 ;
			RECT	122.657 34.05 122.689 34.114 ;
			RECT	122.825 34.05 122.857 34.114 ;
			RECT	122.993 34.05 123.025 34.114 ;
			RECT	123.161 34.05 123.193 34.114 ;
			RECT	123.329 34.05 123.361 34.114 ;
			RECT	123.497 34.05 123.529 34.114 ;
			RECT	123.665 34.05 123.697 34.114 ;
			RECT	123.833 34.05 123.865 34.114 ;
			RECT	124.001 34.05 124.033 34.114 ;
			RECT	124.169 34.05 124.201 34.114 ;
			RECT	124.337 34.05 124.369 34.114 ;
			RECT	124.505 34.05 124.537 34.114 ;
			RECT	124.673 34.05 124.705 34.114 ;
			RECT	124.841 34.05 124.873 34.114 ;
			RECT	125.009 34.05 125.041 34.114 ;
			RECT	125.177 34.05 125.209 34.114 ;
			RECT	125.345 34.05 125.377 34.114 ;
			RECT	125.513 34.05 125.545 34.114 ;
			RECT	125.681 34.05 125.713 34.114 ;
			RECT	125.849 34.05 125.881 34.114 ;
			RECT	126.017 34.05 126.049 34.114 ;
			RECT	126.185 34.05 126.217 34.114 ;
			RECT	126.353 34.05 126.385 34.114 ;
			RECT	126.521 34.05 126.553 34.114 ;
			RECT	126.689 34.05 126.721 34.114 ;
			RECT	126.857 34.05 126.889 34.114 ;
			RECT	127.025 34.05 127.057 34.114 ;
			RECT	127.193 34.05 127.225 34.114 ;
			RECT	127.361 34.05 127.393 34.114 ;
			RECT	127.529 34.05 127.561 34.114 ;
			RECT	127.697 34.05 127.729 34.114 ;
			RECT	127.865 34.05 127.897 34.114 ;
			RECT	128.033 34.05 128.065 34.114 ;
			RECT	128.201 34.05 128.233 34.114 ;
			RECT	128.369 34.05 128.401 34.114 ;
			RECT	128.537 34.05 128.569 34.114 ;
			RECT	128.705 34.05 128.737 34.114 ;
			RECT	128.873 34.05 128.905 34.114 ;
			RECT	129.041 34.05 129.073 34.114 ;
			RECT	129.209 34.05 129.241 34.114 ;
			RECT	129.377 34.05 129.409 34.114 ;
			RECT	129.545 34.05 129.577 34.114 ;
			RECT	129.713 34.05 129.745 34.114 ;
			RECT	129.881 34.05 129.913 34.114 ;
			RECT	130.049 34.05 130.081 34.114 ;
			RECT	130.217 34.05 130.249 34.114 ;
			RECT	130.385 34.05 130.417 34.114 ;
			RECT	130.553 34.05 130.585 34.114 ;
			RECT	130.721 34.05 130.753 34.114 ;
			RECT	130.889 34.05 130.921 34.114 ;
			RECT	131.057 34.05 131.089 34.114 ;
			RECT	131.225 34.05 131.257 34.114 ;
			RECT	131.393 34.05 131.425 34.114 ;
			RECT	131.561 34.05 131.593 34.114 ;
			RECT	131.729 34.05 131.761 34.114 ;
			RECT	131.897 34.05 131.929 34.114 ;
			RECT	132.065 34.05 132.097 34.114 ;
			RECT	132.233 34.05 132.265 34.114 ;
			RECT	132.401 34.05 132.433 34.114 ;
			RECT	132.569 34.05 132.601 34.114 ;
			RECT	132.737 34.05 132.769 34.114 ;
			RECT	132.905 34.05 132.937 34.114 ;
			RECT	133.073 34.05 133.105 34.114 ;
			RECT	133.241 34.05 133.273 34.114 ;
			RECT	133.409 34.05 133.441 34.114 ;
			RECT	133.577 34.05 133.609 34.114 ;
			RECT	133.745 34.05 133.777 34.114 ;
			RECT	133.913 34.05 133.945 34.114 ;
			RECT	134.081 34.05 134.113 34.114 ;
			RECT	134.249 34.05 134.281 34.114 ;
			RECT	134.417 34.05 134.449 34.114 ;
			RECT	134.585 34.05 134.617 34.114 ;
			RECT	134.753 34.05 134.785 34.114 ;
			RECT	134.921 34.05 134.953 34.114 ;
			RECT	135.089 34.05 135.121 34.114 ;
			RECT	135.257 34.05 135.289 34.114 ;
			RECT	135.425 34.05 135.457 34.114 ;
			RECT	135.593 34.05 135.625 34.114 ;
			RECT	135.761 34.05 135.793 34.114 ;
			RECT	135.929 34.05 135.961 34.114 ;
			RECT	136.097 34.05 136.129 34.114 ;
			RECT	136.265 34.05 136.297 34.114 ;
			RECT	136.433 34.05 136.465 34.114 ;
			RECT	136.601 34.05 136.633 34.114 ;
			RECT	136.769 34.05 136.801 34.114 ;
			RECT	136.937 34.05 136.969 34.114 ;
			RECT	137.105 34.05 137.137 34.114 ;
			RECT	137.273 34.05 137.305 34.114 ;
			RECT	137.441 34.05 137.473 34.114 ;
			RECT	137.609 34.05 137.641 34.114 ;
			RECT	137.777 34.05 137.809 34.114 ;
			RECT	137.945 34.05 137.977 34.114 ;
			RECT	138.113 34.05 138.145 34.114 ;
			RECT	138.281 34.05 138.313 34.114 ;
			RECT	138.449 34.05 138.481 34.114 ;
			RECT	138.617 34.05 138.649 34.114 ;
			RECT	138.785 34.05 138.817 34.114 ;
			RECT	138.953 34.05 138.985 34.114 ;
			RECT	139.121 34.05 139.153 34.114 ;
			RECT	139.289 34.05 139.321 34.114 ;
			RECT	139.457 34.05 139.489 34.114 ;
			RECT	139.625 34.05 139.657 34.114 ;
			RECT	139.793 34.05 139.825 34.114 ;
			RECT	139.961 34.05 139.993 34.114 ;
			RECT	140.129 34.05 140.161 34.114 ;
			RECT	140.297 34.05 140.329 34.114 ;
			RECT	140.465 34.05 140.497 34.114 ;
			RECT	140.633 34.05 140.665 34.114 ;
			RECT	140.801 34.05 140.833 34.114 ;
			RECT	140.969 34.05 141.001 34.114 ;
			RECT	141.137 34.05 141.169 34.114 ;
			RECT	141.305 34.05 141.337 34.114 ;
			RECT	141.473 34.05 141.505 34.114 ;
			RECT	141.641 34.05 141.673 34.114 ;
			RECT	141.809 34.05 141.841 34.114 ;
			RECT	141.977 34.05 142.009 34.114 ;
			RECT	142.145 34.05 142.177 34.114 ;
			RECT	142.313 34.05 142.345 34.114 ;
			RECT	142.481 34.05 142.513 34.114 ;
			RECT	142.649 34.05 142.681 34.114 ;
			RECT	142.817 34.05 142.849 34.114 ;
			RECT	142.985 34.05 143.017 34.114 ;
			RECT	143.153 34.05 143.185 34.114 ;
			RECT	143.321 34.05 143.353 34.114 ;
			RECT	143.489 34.05 143.521 34.114 ;
			RECT	143.657 34.05 143.689 34.114 ;
			RECT	143.825 34.05 143.857 34.114 ;
			RECT	143.993 34.05 144.025 34.114 ;
			RECT	144.161 34.05 144.193 34.114 ;
			RECT	144.329 34.05 144.361 34.114 ;
			RECT	144.497 34.05 144.529 34.114 ;
			RECT	144.665 34.05 144.697 34.114 ;
			RECT	144.833 34.05 144.865 34.114 ;
			RECT	145.001 34.05 145.033 34.114 ;
			RECT	145.169 34.05 145.201 34.114 ;
			RECT	145.337 34.05 145.369 34.114 ;
			RECT	145.505 34.05 145.537 34.114 ;
			RECT	145.673 34.05 145.705 34.114 ;
			RECT	145.841 34.05 145.873 34.114 ;
			RECT	146.009 34.05 146.041 34.114 ;
			RECT	146.177 34.05 146.209 34.114 ;
			RECT	146.345 34.05 146.377 34.114 ;
			RECT	146.513 34.05 146.545 34.114 ;
			RECT	146.681 34.05 146.713 34.114 ;
			RECT	146.849 34.05 146.881 34.114 ;
			RECT	147.017 34.05 147.049 34.114 ;
			RECT	147.185 34.05 147.217 34.114 ;
			RECT	147.309 34.05 147.373 34.114 ;
			RECT	147.611 34.05 147.643 34.114 ;
			RECT	147.811 34.05 147.843 34.114 ;
			RECT	149.918 34.05 149.95 34.114 ;
			RECT	150.576 34.05 150.608 34.114 ;
			RECT	151.908 34.05 151.94 34.114 ;
			RECT	153.464 34.05 153.496 34.114 ;
			RECT	153.801 34.05 153.833 34.114 ;
			RECT	153.967 34.05 154.031 34.114 ;
			RECT	156.357 34.05 156.389 34.114 ;
			RECT	156.557 34.05 156.589 34.114 ;
			RECT	156.827 34.05 156.891 34.114 ;
			RECT	156.983 34.05 157.015 34.114 ;
			RECT	157.151 34.05 157.183 34.114 ;
			RECT	157.319 34.05 157.351 34.114 ;
			RECT	157.487 34.05 157.519 34.114 ;
			RECT	157.655 34.05 157.687 34.114 ;
			RECT	157.823 34.05 157.855 34.114 ;
			RECT	157.991 34.05 158.023 34.114 ;
			RECT	158.159 34.05 158.191 34.114 ;
			RECT	158.327 34.05 158.359 34.114 ;
			RECT	158.495 34.05 158.527 34.114 ;
			RECT	158.663 34.05 158.695 34.114 ;
			RECT	158.831 34.05 158.863 34.114 ;
			RECT	158.999 34.05 159.031 34.114 ;
			RECT	159.167 34.05 159.199 34.114 ;
			RECT	159.335 34.05 159.367 34.114 ;
			RECT	159.503 34.05 159.535 34.114 ;
			RECT	159.671 34.05 159.703 34.114 ;
			RECT	159.839 34.05 159.871 34.114 ;
			RECT	160.007 34.05 160.039 34.114 ;
			RECT	160.175 34.05 160.207 34.114 ;
			RECT	160.343 34.05 160.375 34.114 ;
			RECT	160.511 34.05 160.543 34.114 ;
			RECT	160.679 34.05 160.711 34.114 ;
			RECT	160.847 34.05 160.879 34.114 ;
			RECT	161.015 34.05 161.047 34.114 ;
			RECT	161.183 34.05 161.215 34.114 ;
			RECT	161.351 34.05 161.383 34.114 ;
			RECT	161.519 34.05 161.551 34.114 ;
			RECT	161.687 34.05 161.719 34.114 ;
			RECT	161.855 34.05 161.887 34.114 ;
			RECT	162.023 34.05 162.055 34.114 ;
			RECT	162.191 34.05 162.223 34.114 ;
			RECT	162.359 34.05 162.391 34.114 ;
			RECT	162.527 34.05 162.559 34.114 ;
			RECT	162.695 34.05 162.727 34.114 ;
			RECT	162.863 34.05 162.895 34.114 ;
			RECT	163.031 34.05 163.063 34.114 ;
			RECT	163.199 34.05 163.231 34.114 ;
			RECT	163.367 34.05 163.399 34.114 ;
			RECT	163.535 34.05 163.567 34.114 ;
			RECT	163.703 34.05 163.735 34.114 ;
			RECT	163.871 34.05 163.903 34.114 ;
			RECT	164.039 34.05 164.071 34.114 ;
			RECT	164.207 34.05 164.239 34.114 ;
			RECT	164.375 34.05 164.407 34.114 ;
			RECT	164.543 34.05 164.575 34.114 ;
			RECT	164.711 34.05 164.743 34.114 ;
			RECT	164.879 34.05 164.911 34.114 ;
			RECT	165.047 34.05 165.079 34.114 ;
			RECT	165.215 34.05 165.247 34.114 ;
			RECT	165.383 34.05 165.415 34.114 ;
			RECT	165.551 34.05 165.583 34.114 ;
			RECT	165.719 34.05 165.751 34.114 ;
			RECT	165.887 34.05 165.919 34.114 ;
			RECT	166.055 34.05 166.087 34.114 ;
			RECT	166.223 34.05 166.255 34.114 ;
			RECT	166.391 34.05 166.423 34.114 ;
			RECT	166.559 34.05 166.591 34.114 ;
			RECT	166.727 34.05 166.759 34.114 ;
			RECT	166.895 34.05 166.927 34.114 ;
			RECT	167.063 34.05 167.095 34.114 ;
			RECT	167.231 34.05 167.263 34.114 ;
			RECT	167.399 34.05 167.431 34.114 ;
			RECT	167.567 34.05 167.599 34.114 ;
			RECT	167.735 34.05 167.767 34.114 ;
			RECT	167.903 34.05 167.935 34.114 ;
			RECT	168.071 34.05 168.103 34.114 ;
			RECT	168.239 34.05 168.271 34.114 ;
			RECT	168.407 34.05 168.439 34.114 ;
			RECT	168.575 34.05 168.607 34.114 ;
			RECT	168.743 34.05 168.775 34.114 ;
			RECT	168.911 34.05 168.943 34.114 ;
			RECT	169.079 34.05 169.111 34.114 ;
			RECT	169.247 34.05 169.279 34.114 ;
			RECT	169.415 34.05 169.447 34.114 ;
			RECT	169.583 34.05 169.615 34.114 ;
			RECT	169.751 34.05 169.783 34.114 ;
			RECT	169.919 34.05 169.951 34.114 ;
			RECT	170.087 34.05 170.119 34.114 ;
			RECT	170.255 34.05 170.287 34.114 ;
			RECT	170.423 34.05 170.455 34.114 ;
			RECT	170.591 34.05 170.623 34.114 ;
			RECT	170.759 34.05 170.791 34.114 ;
			RECT	170.927 34.05 170.959 34.114 ;
			RECT	171.095 34.05 171.127 34.114 ;
			RECT	171.263 34.05 171.295 34.114 ;
			RECT	171.431 34.05 171.463 34.114 ;
			RECT	171.599 34.05 171.631 34.114 ;
			RECT	171.767 34.05 171.799 34.114 ;
			RECT	171.935 34.05 171.967 34.114 ;
			RECT	172.103 34.05 172.135 34.114 ;
			RECT	172.271 34.05 172.303 34.114 ;
			RECT	172.439 34.05 172.471 34.114 ;
			RECT	172.607 34.05 172.639 34.114 ;
			RECT	172.775 34.05 172.807 34.114 ;
			RECT	172.943 34.05 172.975 34.114 ;
			RECT	173.111 34.05 173.143 34.114 ;
			RECT	173.279 34.05 173.311 34.114 ;
			RECT	173.447 34.05 173.479 34.114 ;
			RECT	173.615 34.05 173.647 34.114 ;
			RECT	173.783 34.05 173.815 34.114 ;
			RECT	173.951 34.05 173.983 34.114 ;
			RECT	174.119 34.05 174.151 34.114 ;
			RECT	174.287 34.05 174.319 34.114 ;
			RECT	174.455 34.05 174.487 34.114 ;
			RECT	174.623 34.05 174.655 34.114 ;
			RECT	174.791 34.05 174.823 34.114 ;
			RECT	174.959 34.05 174.991 34.114 ;
			RECT	175.127 34.05 175.159 34.114 ;
			RECT	175.295 34.05 175.327 34.114 ;
			RECT	175.463 34.05 175.495 34.114 ;
			RECT	175.631 34.05 175.663 34.114 ;
			RECT	175.799 34.05 175.831 34.114 ;
			RECT	175.967 34.05 175.999 34.114 ;
			RECT	176.135 34.05 176.167 34.114 ;
			RECT	176.303 34.05 176.335 34.114 ;
			RECT	176.471 34.05 176.503 34.114 ;
			RECT	176.639 34.05 176.671 34.114 ;
			RECT	176.807 34.05 176.839 34.114 ;
			RECT	176.975 34.05 177.007 34.114 ;
			RECT	177.143 34.05 177.175 34.114 ;
			RECT	177.311 34.05 177.343 34.114 ;
			RECT	177.479 34.05 177.511 34.114 ;
			RECT	177.647 34.05 177.679 34.114 ;
			RECT	177.815 34.05 177.847 34.114 ;
			RECT	177.983 34.05 178.015 34.114 ;
			RECT	178.151 34.05 178.183 34.114 ;
			RECT	178.319 34.05 178.351 34.114 ;
			RECT	178.487 34.05 178.519 34.114 ;
			RECT	178.655 34.05 178.687 34.114 ;
			RECT	178.823 34.05 178.855 34.114 ;
			RECT	178.991 34.05 179.023 34.114 ;
			RECT	179.159 34.05 179.191 34.114 ;
			RECT	179.327 34.05 179.359 34.114 ;
			RECT	179.495 34.05 179.527 34.114 ;
			RECT	179.663 34.05 179.695 34.114 ;
			RECT	179.831 34.05 179.863 34.114 ;
			RECT	179.999 34.05 180.031 34.114 ;
			RECT	180.167 34.05 180.199 34.114 ;
			RECT	180.335 34.05 180.367 34.114 ;
			RECT	180.503 34.05 180.535 34.114 ;
			RECT	180.671 34.05 180.703 34.114 ;
			RECT	180.839 34.05 180.871 34.114 ;
			RECT	181.007 34.05 181.039 34.114 ;
			RECT	181.175 34.05 181.207 34.114 ;
			RECT	181.343 34.05 181.375 34.114 ;
			RECT	181.511 34.05 181.543 34.114 ;
			RECT	181.679 34.05 181.711 34.114 ;
			RECT	181.847 34.05 181.879 34.114 ;
			RECT	182.015 34.05 182.047 34.114 ;
			RECT	182.183 34.05 182.215 34.114 ;
			RECT	182.351 34.05 182.383 34.114 ;
			RECT	182.519 34.05 182.551 34.114 ;
			RECT	182.687 34.05 182.719 34.114 ;
			RECT	182.855 34.05 182.887 34.114 ;
			RECT	183.023 34.05 183.055 34.114 ;
			RECT	183.191 34.05 183.223 34.114 ;
			RECT	183.359 34.05 183.391 34.114 ;
			RECT	183.527 34.05 183.559 34.114 ;
			RECT	183.695 34.05 183.727 34.114 ;
			RECT	183.863 34.05 183.895 34.114 ;
			RECT	184.031 34.05 184.063 34.114 ;
			RECT	184.199 34.05 184.231 34.114 ;
			RECT	184.367 34.05 184.399 34.114 ;
			RECT	184.535 34.05 184.567 34.114 ;
			RECT	184.703 34.05 184.735 34.114 ;
			RECT	184.871 34.05 184.903 34.114 ;
			RECT	185.039 34.05 185.071 34.114 ;
			RECT	185.207 34.05 185.239 34.114 ;
			RECT	185.375 34.05 185.407 34.114 ;
			RECT	185.543 34.05 185.575 34.114 ;
			RECT	185.711 34.05 185.743 34.114 ;
			RECT	185.879 34.05 185.911 34.114 ;
			RECT	186.047 34.05 186.079 34.114 ;
			RECT	186.215 34.05 186.247 34.114 ;
			RECT	186.383 34.05 186.415 34.114 ;
			RECT	186.551 34.05 186.583 34.114 ;
			RECT	186.719 34.05 186.751 34.114 ;
			RECT	186.887 34.05 186.919 34.114 ;
			RECT	187.055 34.05 187.087 34.114 ;
			RECT	187.223 34.05 187.255 34.114 ;
			RECT	187.391 34.05 187.423 34.114 ;
			RECT	187.559 34.05 187.591 34.114 ;
			RECT	187.727 34.05 187.759 34.114 ;
			RECT	187.895 34.05 187.927 34.114 ;
			RECT	188.063 34.05 188.095 34.114 ;
			RECT	188.231 34.05 188.263 34.114 ;
			RECT	188.399 34.05 188.431 34.114 ;
			RECT	188.567 34.05 188.599 34.114 ;
			RECT	188.735 34.05 188.767 34.114 ;
			RECT	188.903 34.05 188.935 34.114 ;
			RECT	189.071 34.05 189.103 34.114 ;
			RECT	189.239 34.05 189.271 34.114 ;
			RECT	189.407 34.05 189.439 34.114 ;
			RECT	189.575 34.05 189.607 34.114 ;
			RECT	189.743 34.05 189.775 34.114 ;
			RECT	189.911 34.05 189.943 34.114 ;
			RECT	190.079 34.05 190.111 34.114 ;
			RECT	190.247 34.05 190.279 34.114 ;
			RECT	190.415 34.05 190.447 34.114 ;
			RECT	190.583 34.05 190.615 34.114 ;
			RECT	190.751 34.05 190.783 34.114 ;
			RECT	190.919 34.05 190.951 34.114 ;
			RECT	191.087 34.05 191.119 34.114 ;
			RECT	191.255 34.05 191.287 34.114 ;
			RECT	191.423 34.05 191.455 34.114 ;
			RECT	191.591 34.05 191.623 34.114 ;
			RECT	191.759 34.05 191.791 34.114 ;
			RECT	191.927 34.05 191.959 34.114 ;
			RECT	192.095 34.05 192.127 34.114 ;
			RECT	192.263 34.05 192.295 34.114 ;
			RECT	192.431 34.05 192.463 34.114 ;
			RECT	192.599 34.05 192.631 34.114 ;
			RECT	192.767 34.05 192.799 34.114 ;
			RECT	192.935 34.05 192.967 34.114 ;
			RECT	193.103 34.05 193.135 34.114 ;
			RECT	193.271 34.05 193.303 34.114 ;
			RECT	193.439 34.05 193.471 34.114 ;
			RECT	193.607 34.05 193.639 34.114 ;
			RECT	193.775 34.05 193.807 34.114 ;
			RECT	193.943 34.05 193.975 34.114 ;
			RECT	194.111 34.05 194.143 34.114 ;
			RECT	194.279 34.05 194.311 34.114 ;
			RECT	194.447 34.05 194.479 34.114 ;
			RECT	194.615 34.05 194.647 34.114 ;
			RECT	194.783 34.05 194.815 34.114 ;
			RECT	194.951 34.05 194.983 34.114 ;
			RECT	195.119 34.05 195.151 34.114 ;
			RECT	195.287 34.05 195.319 34.114 ;
			RECT	195.455 34.05 195.487 34.114 ;
			RECT	195.623 34.05 195.655 34.114 ;
			RECT	195.791 34.05 195.823 34.114 ;
			RECT	195.959 34.05 195.991 34.114 ;
			RECT	196.127 34.05 196.159 34.114 ;
			RECT	196.295 34.05 196.327 34.114 ;
			RECT	196.463 34.05 196.495 34.114 ;
			RECT	196.631 34.05 196.663 34.114 ;
			RECT	196.799 34.05 196.831 34.114 ;
			RECT	196.967 34.05 196.999 34.114 ;
			RECT	197.135 34.05 197.167 34.114 ;
			RECT	197.303 34.05 197.335 34.114 ;
			RECT	197.471 34.05 197.503 34.114 ;
			RECT	197.639 34.05 197.671 34.114 ;
			RECT	197.807 34.05 197.839 34.114 ;
			RECT	197.975 34.05 198.007 34.114 ;
			RECT	198.143 34.05 198.175 34.114 ;
			RECT	198.311 34.05 198.343 34.114 ;
			RECT	198.479 34.05 198.511 34.114 ;
			RECT	198.647 34.05 198.679 34.114 ;
			RECT	198.815 34.05 198.847 34.114 ;
			RECT	198.983 34.05 199.015 34.114 ;
			RECT	199.151 34.05 199.183 34.114 ;
			RECT	199.319 34.05 199.351 34.114 ;
			RECT	199.487 34.05 199.519 34.114 ;
			RECT	199.655 34.05 199.687 34.114 ;
			RECT	199.823 34.05 199.855 34.114 ;
			RECT	199.991 34.05 200.023 34.114 ;
			RECT	200.9 34.05 200.932 34.114 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 34.432 201.665 34.552 ;
			LAYER	J3 ;
			RECT	1.645 34.46 1.709 34.524 ;
			RECT	2.323 34.46 2.387 34.524 ;
			RECT	3.438 34.476 3.47 34.508 ;
			RECT	4.195 34.46 4.227 34.524 ;
			RECT	4.354 34.46 4.386 34.524 ;
			RECT	4.959 34.46 4.991 34.524 ;
			RECT	6.179 34.46 6.211 34.524 ;
			RECT	6.347 34.46 6.379 34.524 ;
			RECT	6.515 34.46 6.547 34.524 ;
			RECT	6.683 34.46 6.715 34.524 ;
			RECT	6.851 34.46 6.883 34.524 ;
			RECT	7.019 34.46 7.051 34.524 ;
			RECT	7.187 34.46 7.219 34.524 ;
			RECT	7.355 34.46 7.387 34.524 ;
			RECT	7.523 34.46 7.555 34.524 ;
			RECT	7.691 34.46 7.723 34.524 ;
			RECT	7.859 34.46 7.891 34.524 ;
			RECT	8.027 34.46 8.059 34.524 ;
			RECT	8.195 34.46 8.227 34.524 ;
			RECT	8.363 34.46 8.395 34.524 ;
			RECT	8.531 34.46 8.563 34.524 ;
			RECT	8.699 34.46 8.731 34.524 ;
			RECT	8.867 34.46 8.899 34.524 ;
			RECT	9.035 34.46 9.067 34.524 ;
			RECT	9.203 34.46 9.235 34.524 ;
			RECT	9.371 34.46 9.403 34.524 ;
			RECT	9.539 34.46 9.571 34.524 ;
			RECT	9.707 34.46 9.739 34.524 ;
			RECT	9.875 34.46 9.907 34.524 ;
			RECT	10.043 34.46 10.075 34.524 ;
			RECT	10.211 34.46 10.243 34.524 ;
			RECT	10.379 34.46 10.411 34.524 ;
			RECT	10.547 34.46 10.579 34.524 ;
			RECT	10.715 34.46 10.747 34.524 ;
			RECT	10.883 34.46 10.915 34.524 ;
			RECT	11.051 34.46 11.083 34.524 ;
			RECT	11.219 34.46 11.251 34.524 ;
			RECT	11.387 34.46 11.419 34.524 ;
			RECT	11.555 34.46 11.587 34.524 ;
			RECT	11.723 34.46 11.755 34.524 ;
			RECT	11.891 34.46 11.923 34.524 ;
			RECT	12.059 34.46 12.091 34.524 ;
			RECT	12.227 34.46 12.259 34.524 ;
			RECT	12.395 34.46 12.427 34.524 ;
			RECT	12.563 34.46 12.595 34.524 ;
			RECT	12.731 34.46 12.763 34.524 ;
			RECT	12.899 34.46 12.931 34.524 ;
			RECT	13.067 34.46 13.099 34.524 ;
			RECT	13.235 34.46 13.267 34.524 ;
			RECT	13.403 34.46 13.435 34.524 ;
			RECT	13.571 34.46 13.603 34.524 ;
			RECT	13.739 34.46 13.771 34.524 ;
			RECT	13.907 34.46 13.939 34.524 ;
			RECT	14.075 34.46 14.107 34.524 ;
			RECT	14.243 34.46 14.275 34.524 ;
			RECT	14.411 34.46 14.443 34.524 ;
			RECT	14.579 34.46 14.611 34.524 ;
			RECT	14.747 34.46 14.779 34.524 ;
			RECT	14.915 34.46 14.947 34.524 ;
			RECT	15.083 34.46 15.115 34.524 ;
			RECT	15.251 34.46 15.283 34.524 ;
			RECT	15.419 34.46 15.451 34.524 ;
			RECT	15.587 34.46 15.619 34.524 ;
			RECT	15.755 34.46 15.787 34.524 ;
			RECT	15.923 34.46 15.955 34.524 ;
			RECT	16.091 34.46 16.123 34.524 ;
			RECT	16.259 34.46 16.291 34.524 ;
			RECT	16.427 34.46 16.459 34.524 ;
			RECT	16.595 34.46 16.627 34.524 ;
			RECT	16.763 34.46 16.795 34.524 ;
			RECT	16.931 34.46 16.963 34.524 ;
			RECT	17.099 34.46 17.131 34.524 ;
			RECT	17.267 34.46 17.299 34.524 ;
			RECT	17.435 34.46 17.467 34.524 ;
			RECT	17.603 34.46 17.635 34.524 ;
			RECT	17.771 34.46 17.803 34.524 ;
			RECT	17.939 34.46 17.971 34.524 ;
			RECT	18.107 34.46 18.139 34.524 ;
			RECT	18.275 34.46 18.307 34.524 ;
			RECT	18.443 34.46 18.475 34.524 ;
			RECT	18.611 34.46 18.643 34.524 ;
			RECT	18.779 34.46 18.811 34.524 ;
			RECT	18.947 34.46 18.979 34.524 ;
			RECT	19.115 34.46 19.147 34.524 ;
			RECT	19.283 34.46 19.315 34.524 ;
			RECT	19.451 34.46 19.483 34.524 ;
			RECT	19.619 34.46 19.651 34.524 ;
			RECT	19.787 34.46 19.819 34.524 ;
			RECT	19.955 34.46 19.987 34.524 ;
			RECT	20.123 34.46 20.155 34.524 ;
			RECT	20.291 34.46 20.323 34.524 ;
			RECT	20.459 34.46 20.491 34.524 ;
			RECT	20.627 34.46 20.659 34.524 ;
			RECT	20.795 34.46 20.827 34.524 ;
			RECT	20.963 34.46 20.995 34.524 ;
			RECT	21.131 34.46 21.163 34.524 ;
			RECT	21.299 34.46 21.331 34.524 ;
			RECT	21.467 34.46 21.499 34.524 ;
			RECT	21.635 34.46 21.667 34.524 ;
			RECT	21.803 34.46 21.835 34.524 ;
			RECT	21.971 34.46 22.003 34.524 ;
			RECT	22.139 34.46 22.171 34.524 ;
			RECT	22.307 34.46 22.339 34.524 ;
			RECT	22.475 34.46 22.507 34.524 ;
			RECT	22.643 34.46 22.675 34.524 ;
			RECT	22.811 34.46 22.843 34.524 ;
			RECT	22.979 34.46 23.011 34.524 ;
			RECT	23.147 34.46 23.179 34.524 ;
			RECT	23.315 34.46 23.347 34.524 ;
			RECT	23.483 34.46 23.515 34.524 ;
			RECT	23.651 34.46 23.683 34.524 ;
			RECT	23.819 34.46 23.851 34.524 ;
			RECT	23.987 34.46 24.019 34.524 ;
			RECT	24.155 34.46 24.187 34.524 ;
			RECT	24.323 34.46 24.355 34.524 ;
			RECT	24.491 34.46 24.523 34.524 ;
			RECT	24.659 34.46 24.691 34.524 ;
			RECT	24.827 34.46 24.859 34.524 ;
			RECT	24.995 34.46 25.027 34.524 ;
			RECT	25.163 34.46 25.195 34.524 ;
			RECT	25.331 34.46 25.363 34.524 ;
			RECT	25.499 34.46 25.531 34.524 ;
			RECT	25.667 34.46 25.699 34.524 ;
			RECT	25.835 34.46 25.867 34.524 ;
			RECT	26.003 34.46 26.035 34.524 ;
			RECT	26.171 34.46 26.203 34.524 ;
			RECT	26.339 34.46 26.371 34.524 ;
			RECT	26.507 34.46 26.539 34.524 ;
			RECT	26.675 34.46 26.707 34.524 ;
			RECT	26.843 34.46 26.875 34.524 ;
			RECT	27.011 34.46 27.043 34.524 ;
			RECT	27.179 34.46 27.211 34.524 ;
			RECT	27.347 34.46 27.379 34.524 ;
			RECT	27.515 34.46 27.547 34.524 ;
			RECT	27.683 34.46 27.715 34.524 ;
			RECT	27.851 34.46 27.883 34.524 ;
			RECT	28.019 34.46 28.051 34.524 ;
			RECT	28.187 34.46 28.219 34.524 ;
			RECT	28.355 34.46 28.387 34.524 ;
			RECT	28.523 34.46 28.555 34.524 ;
			RECT	28.691 34.46 28.723 34.524 ;
			RECT	28.859 34.46 28.891 34.524 ;
			RECT	29.027 34.46 29.059 34.524 ;
			RECT	29.195 34.46 29.227 34.524 ;
			RECT	29.363 34.46 29.395 34.524 ;
			RECT	29.531 34.46 29.563 34.524 ;
			RECT	29.699 34.46 29.731 34.524 ;
			RECT	29.867 34.46 29.899 34.524 ;
			RECT	30.035 34.46 30.067 34.524 ;
			RECT	30.203 34.46 30.235 34.524 ;
			RECT	30.371 34.46 30.403 34.524 ;
			RECT	30.539 34.46 30.571 34.524 ;
			RECT	30.707 34.46 30.739 34.524 ;
			RECT	30.875 34.46 30.907 34.524 ;
			RECT	31.043 34.46 31.075 34.524 ;
			RECT	31.211 34.46 31.243 34.524 ;
			RECT	31.379 34.46 31.411 34.524 ;
			RECT	31.547 34.46 31.579 34.524 ;
			RECT	31.715 34.46 31.747 34.524 ;
			RECT	31.883 34.46 31.915 34.524 ;
			RECT	32.051 34.46 32.083 34.524 ;
			RECT	32.219 34.46 32.251 34.524 ;
			RECT	32.387 34.46 32.419 34.524 ;
			RECT	32.555 34.46 32.587 34.524 ;
			RECT	32.723 34.46 32.755 34.524 ;
			RECT	32.891 34.46 32.923 34.524 ;
			RECT	33.059 34.46 33.091 34.524 ;
			RECT	33.227 34.46 33.259 34.524 ;
			RECT	33.395 34.46 33.427 34.524 ;
			RECT	33.563 34.46 33.595 34.524 ;
			RECT	33.731 34.46 33.763 34.524 ;
			RECT	33.899 34.46 33.931 34.524 ;
			RECT	34.067 34.46 34.099 34.524 ;
			RECT	34.235 34.46 34.267 34.524 ;
			RECT	34.403 34.46 34.435 34.524 ;
			RECT	34.571 34.46 34.603 34.524 ;
			RECT	34.739 34.46 34.771 34.524 ;
			RECT	34.907 34.46 34.939 34.524 ;
			RECT	35.075 34.46 35.107 34.524 ;
			RECT	35.243 34.46 35.275 34.524 ;
			RECT	35.411 34.46 35.443 34.524 ;
			RECT	35.579 34.46 35.611 34.524 ;
			RECT	35.747 34.46 35.779 34.524 ;
			RECT	35.915 34.46 35.947 34.524 ;
			RECT	36.083 34.46 36.115 34.524 ;
			RECT	36.251 34.46 36.283 34.524 ;
			RECT	36.419 34.46 36.451 34.524 ;
			RECT	36.587 34.46 36.619 34.524 ;
			RECT	36.755 34.46 36.787 34.524 ;
			RECT	36.923 34.46 36.955 34.524 ;
			RECT	37.091 34.46 37.123 34.524 ;
			RECT	37.259 34.46 37.291 34.524 ;
			RECT	37.427 34.46 37.459 34.524 ;
			RECT	37.595 34.46 37.627 34.524 ;
			RECT	37.763 34.46 37.795 34.524 ;
			RECT	37.931 34.46 37.963 34.524 ;
			RECT	38.099 34.46 38.131 34.524 ;
			RECT	38.267 34.46 38.299 34.524 ;
			RECT	38.435 34.46 38.467 34.524 ;
			RECT	38.603 34.46 38.635 34.524 ;
			RECT	38.771 34.46 38.803 34.524 ;
			RECT	38.939 34.46 38.971 34.524 ;
			RECT	39.107 34.46 39.139 34.524 ;
			RECT	39.275 34.46 39.307 34.524 ;
			RECT	39.443 34.46 39.475 34.524 ;
			RECT	39.611 34.46 39.643 34.524 ;
			RECT	39.779 34.46 39.811 34.524 ;
			RECT	39.947 34.46 39.979 34.524 ;
			RECT	40.115 34.46 40.147 34.524 ;
			RECT	40.283 34.46 40.315 34.524 ;
			RECT	40.451 34.46 40.483 34.524 ;
			RECT	40.619 34.46 40.651 34.524 ;
			RECT	40.787 34.46 40.819 34.524 ;
			RECT	40.955 34.46 40.987 34.524 ;
			RECT	41.123 34.46 41.155 34.524 ;
			RECT	41.291 34.46 41.323 34.524 ;
			RECT	41.459 34.46 41.491 34.524 ;
			RECT	41.627 34.46 41.659 34.524 ;
			RECT	41.795 34.46 41.827 34.524 ;
			RECT	41.963 34.46 41.995 34.524 ;
			RECT	42.131 34.46 42.163 34.524 ;
			RECT	42.299 34.46 42.331 34.524 ;
			RECT	42.467 34.46 42.499 34.524 ;
			RECT	42.635 34.46 42.667 34.524 ;
			RECT	42.803 34.46 42.835 34.524 ;
			RECT	42.971 34.46 43.003 34.524 ;
			RECT	43.139 34.46 43.171 34.524 ;
			RECT	43.307 34.46 43.339 34.524 ;
			RECT	43.475 34.46 43.507 34.524 ;
			RECT	43.643 34.46 43.675 34.524 ;
			RECT	43.811 34.46 43.843 34.524 ;
			RECT	43.979 34.46 44.011 34.524 ;
			RECT	44.147 34.46 44.179 34.524 ;
			RECT	44.315 34.46 44.347 34.524 ;
			RECT	44.483 34.46 44.515 34.524 ;
			RECT	44.651 34.46 44.683 34.524 ;
			RECT	44.819 34.46 44.851 34.524 ;
			RECT	44.987 34.46 45.019 34.524 ;
			RECT	45.155 34.46 45.187 34.524 ;
			RECT	45.323 34.46 45.355 34.524 ;
			RECT	45.491 34.46 45.523 34.524 ;
			RECT	45.659 34.46 45.691 34.524 ;
			RECT	45.827 34.46 45.859 34.524 ;
			RECT	45.995 34.46 46.027 34.524 ;
			RECT	46.163 34.46 46.195 34.524 ;
			RECT	46.331 34.46 46.363 34.524 ;
			RECT	46.499 34.46 46.531 34.524 ;
			RECT	46.667 34.46 46.699 34.524 ;
			RECT	46.835 34.46 46.867 34.524 ;
			RECT	47.003 34.46 47.035 34.524 ;
			RECT	47.171 34.46 47.203 34.524 ;
			RECT	47.339 34.46 47.371 34.524 ;
			RECT	47.507 34.46 47.539 34.524 ;
			RECT	47.675 34.46 47.707 34.524 ;
			RECT	47.843 34.46 47.875 34.524 ;
			RECT	48.011 34.46 48.043 34.524 ;
			RECT	48.179 34.46 48.211 34.524 ;
			RECT	48.347 34.46 48.379 34.524 ;
			RECT	48.515 34.46 48.547 34.524 ;
			RECT	48.683 34.46 48.715 34.524 ;
			RECT	48.851 34.46 48.883 34.524 ;
			RECT	49.019 34.46 49.051 34.524 ;
			RECT	49.187 34.46 49.219 34.524 ;
			RECT	49.311 34.46 49.375 34.524 ;
			RECT	49.613 34.46 49.645 34.524 ;
			RECT	51.92 34.46 51.952 34.524 ;
			RECT	52.221 34.46 52.253 34.524 ;
			RECT	52.968 34.46 53.032 34.524 ;
			RECT	53.91 34.46 53.942 34.524 ;
			RECT	55.969 34.46 56.033 34.524 ;
			RECT	58.559 34.46 58.591 34.524 ;
			RECT	58.829 34.46 58.893 34.524 ;
			RECT	58.985 34.46 59.017 34.524 ;
			RECT	59.153 34.46 59.185 34.524 ;
			RECT	59.321 34.46 59.353 34.524 ;
			RECT	59.489 34.46 59.521 34.524 ;
			RECT	59.657 34.46 59.689 34.524 ;
			RECT	59.825 34.46 59.857 34.524 ;
			RECT	59.993 34.46 60.025 34.524 ;
			RECT	60.161 34.46 60.193 34.524 ;
			RECT	60.329 34.46 60.361 34.524 ;
			RECT	60.497 34.46 60.529 34.524 ;
			RECT	60.665 34.46 60.697 34.524 ;
			RECT	60.833 34.46 60.865 34.524 ;
			RECT	61.001 34.46 61.033 34.524 ;
			RECT	61.169 34.46 61.201 34.524 ;
			RECT	61.337 34.46 61.369 34.524 ;
			RECT	61.505 34.46 61.537 34.524 ;
			RECT	61.673 34.46 61.705 34.524 ;
			RECT	61.841 34.46 61.873 34.524 ;
			RECT	62.009 34.46 62.041 34.524 ;
			RECT	62.177 34.46 62.209 34.524 ;
			RECT	62.345 34.46 62.377 34.524 ;
			RECT	62.513 34.46 62.545 34.524 ;
			RECT	62.681 34.46 62.713 34.524 ;
			RECT	62.849 34.46 62.881 34.524 ;
			RECT	63.017 34.46 63.049 34.524 ;
			RECT	63.185 34.46 63.217 34.524 ;
			RECT	63.353 34.46 63.385 34.524 ;
			RECT	63.521 34.46 63.553 34.524 ;
			RECT	63.689 34.46 63.721 34.524 ;
			RECT	63.857 34.46 63.889 34.524 ;
			RECT	64.025 34.46 64.057 34.524 ;
			RECT	64.193 34.46 64.225 34.524 ;
			RECT	64.361 34.46 64.393 34.524 ;
			RECT	64.529 34.46 64.561 34.524 ;
			RECT	64.697 34.46 64.729 34.524 ;
			RECT	64.865 34.46 64.897 34.524 ;
			RECT	65.033 34.46 65.065 34.524 ;
			RECT	65.201 34.46 65.233 34.524 ;
			RECT	65.369 34.46 65.401 34.524 ;
			RECT	65.537 34.46 65.569 34.524 ;
			RECT	65.705 34.46 65.737 34.524 ;
			RECT	65.873 34.46 65.905 34.524 ;
			RECT	66.041 34.46 66.073 34.524 ;
			RECT	66.209 34.46 66.241 34.524 ;
			RECT	66.377 34.46 66.409 34.524 ;
			RECT	66.545 34.46 66.577 34.524 ;
			RECT	66.713 34.46 66.745 34.524 ;
			RECT	66.881 34.46 66.913 34.524 ;
			RECT	67.049 34.46 67.081 34.524 ;
			RECT	67.217 34.46 67.249 34.524 ;
			RECT	67.385 34.46 67.417 34.524 ;
			RECT	67.553 34.46 67.585 34.524 ;
			RECT	67.721 34.46 67.753 34.524 ;
			RECT	67.889 34.46 67.921 34.524 ;
			RECT	68.057 34.46 68.089 34.524 ;
			RECT	68.225 34.46 68.257 34.524 ;
			RECT	68.393 34.46 68.425 34.524 ;
			RECT	68.561 34.46 68.593 34.524 ;
			RECT	68.729 34.46 68.761 34.524 ;
			RECT	68.897 34.46 68.929 34.524 ;
			RECT	69.065 34.46 69.097 34.524 ;
			RECT	69.233 34.46 69.265 34.524 ;
			RECT	69.401 34.46 69.433 34.524 ;
			RECT	69.569 34.46 69.601 34.524 ;
			RECT	69.737 34.46 69.769 34.524 ;
			RECT	69.905 34.46 69.937 34.524 ;
			RECT	70.073 34.46 70.105 34.524 ;
			RECT	70.241 34.46 70.273 34.524 ;
			RECT	70.409 34.46 70.441 34.524 ;
			RECT	70.577 34.46 70.609 34.524 ;
			RECT	70.745 34.46 70.777 34.524 ;
			RECT	70.913 34.46 70.945 34.524 ;
			RECT	71.081 34.46 71.113 34.524 ;
			RECT	71.249 34.46 71.281 34.524 ;
			RECT	71.417 34.46 71.449 34.524 ;
			RECT	71.585 34.46 71.617 34.524 ;
			RECT	71.753 34.46 71.785 34.524 ;
			RECT	71.921 34.46 71.953 34.524 ;
			RECT	72.089 34.46 72.121 34.524 ;
			RECT	72.257 34.46 72.289 34.524 ;
			RECT	72.425 34.46 72.457 34.524 ;
			RECT	72.593 34.46 72.625 34.524 ;
			RECT	72.761 34.46 72.793 34.524 ;
			RECT	72.929 34.46 72.961 34.524 ;
			RECT	73.097 34.46 73.129 34.524 ;
			RECT	73.265 34.46 73.297 34.524 ;
			RECT	73.433 34.46 73.465 34.524 ;
			RECT	73.601 34.46 73.633 34.524 ;
			RECT	73.769 34.46 73.801 34.524 ;
			RECT	73.937 34.46 73.969 34.524 ;
			RECT	74.105 34.46 74.137 34.524 ;
			RECT	74.273 34.46 74.305 34.524 ;
			RECT	74.441 34.46 74.473 34.524 ;
			RECT	74.609 34.46 74.641 34.524 ;
			RECT	74.777 34.46 74.809 34.524 ;
			RECT	74.945 34.46 74.977 34.524 ;
			RECT	75.113 34.46 75.145 34.524 ;
			RECT	75.281 34.46 75.313 34.524 ;
			RECT	75.449 34.46 75.481 34.524 ;
			RECT	75.617 34.46 75.649 34.524 ;
			RECT	75.785 34.46 75.817 34.524 ;
			RECT	75.953 34.46 75.985 34.524 ;
			RECT	76.121 34.46 76.153 34.524 ;
			RECT	76.289 34.46 76.321 34.524 ;
			RECT	76.457 34.46 76.489 34.524 ;
			RECT	76.625 34.46 76.657 34.524 ;
			RECT	76.793 34.46 76.825 34.524 ;
			RECT	76.961 34.46 76.993 34.524 ;
			RECT	77.129 34.46 77.161 34.524 ;
			RECT	77.297 34.46 77.329 34.524 ;
			RECT	77.465 34.46 77.497 34.524 ;
			RECT	77.633 34.46 77.665 34.524 ;
			RECT	77.801 34.46 77.833 34.524 ;
			RECT	77.969 34.46 78.001 34.524 ;
			RECT	78.137 34.46 78.169 34.524 ;
			RECT	78.305 34.46 78.337 34.524 ;
			RECT	78.473 34.46 78.505 34.524 ;
			RECT	78.641 34.46 78.673 34.524 ;
			RECT	78.809 34.46 78.841 34.524 ;
			RECT	78.977 34.46 79.009 34.524 ;
			RECT	79.145 34.46 79.177 34.524 ;
			RECT	79.313 34.46 79.345 34.524 ;
			RECT	79.481 34.46 79.513 34.524 ;
			RECT	79.649 34.46 79.681 34.524 ;
			RECT	79.817 34.46 79.849 34.524 ;
			RECT	79.985 34.46 80.017 34.524 ;
			RECT	80.153 34.46 80.185 34.524 ;
			RECT	80.321 34.46 80.353 34.524 ;
			RECT	80.489 34.46 80.521 34.524 ;
			RECT	80.657 34.46 80.689 34.524 ;
			RECT	80.825 34.46 80.857 34.524 ;
			RECT	80.993 34.46 81.025 34.524 ;
			RECT	81.161 34.46 81.193 34.524 ;
			RECT	81.329 34.46 81.361 34.524 ;
			RECT	81.497 34.46 81.529 34.524 ;
			RECT	81.665 34.46 81.697 34.524 ;
			RECT	81.833 34.46 81.865 34.524 ;
			RECT	82.001 34.46 82.033 34.524 ;
			RECT	82.169 34.46 82.201 34.524 ;
			RECT	82.337 34.46 82.369 34.524 ;
			RECT	82.505 34.46 82.537 34.524 ;
			RECT	82.673 34.46 82.705 34.524 ;
			RECT	82.841 34.46 82.873 34.524 ;
			RECT	83.009 34.46 83.041 34.524 ;
			RECT	83.177 34.46 83.209 34.524 ;
			RECT	83.345 34.46 83.377 34.524 ;
			RECT	83.513 34.46 83.545 34.524 ;
			RECT	83.681 34.46 83.713 34.524 ;
			RECT	83.849 34.46 83.881 34.524 ;
			RECT	84.017 34.46 84.049 34.524 ;
			RECT	84.185 34.46 84.217 34.524 ;
			RECT	84.353 34.46 84.385 34.524 ;
			RECT	84.521 34.46 84.553 34.524 ;
			RECT	84.689 34.46 84.721 34.524 ;
			RECT	84.857 34.46 84.889 34.524 ;
			RECT	85.025 34.46 85.057 34.524 ;
			RECT	85.193 34.46 85.225 34.524 ;
			RECT	85.361 34.46 85.393 34.524 ;
			RECT	85.529 34.46 85.561 34.524 ;
			RECT	85.697 34.46 85.729 34.524 ;
			RECT	85.865 34.46 85.897 34.524 ;
			RECT	86.033 34.46 86.065 34.524 ;
			RECT	86.201 34.46 86.233 34.524 ;
			RECT	86.369 34.46 86.401 34.524 ;
			RECT	86.537 34.46 86.569 34.524 ;
			RECT	86.705 34.46 86.737 34.524 ;
			RECT	86.873 34.46 86.905 34.524 ;
			RECT	87.041 34.46 87.073 34.524 ;
			RECT	87.209 34.46 87.241 34.524 ;
			RECT	87.377 34.46 87.409 34.524 ;
			RECT	87.545 34.46 87.577 34.524 ;
			RECT	87.713 34.46 87.745 34.524 ;
			RECT	87.881 34.46 87.913 34.524 ;
			RECT	88.049 34.46 88.081 34.524 ;
			RECT	88.217 34.46 88.249 34.524 ;
			RECT	88.385 34.46 88.417 34.524 ;
			RECT	88.553 34.46 88.585 34.524 ;
			RECT	88.721 34.46 88.753 34.524 ;
			RECT	88.889 34.46 88.921 34.524 ;
			RECT	89.057 34.46 89.089 34.524 ;
			RECT	89.225 34.46 89.257 34.524 ;
			RECT	89.393 34.46 89.425 34.524 ;
			RECT	89.561 34.46 89.593 34.524 ;
			RECT	89.729 34.46 89.761 34.524 ;
			RECT	89.897 34.46 89.929 34.524 ;
			RECT	90.065 34.46 90.097 34.524 ;
			RECT	90.233 34.46 90.265 34.524 ;
			RECT	90.401 34.46 90.433 34.524 ;
			RECT	90.569 34.46 90.601 34.524 ;
			RECT	90.737 34.46 90.769 34.524 ;
			RECT	90.905 34.46 90.937 34.524 ;
			RECT	91.073 34.46 91.105 34.524 ;
			RECT	91.241 34.46 91.273 34.524 ;
			RECT	91.409 34.46 91.441 34.524 ;
			RECT	91.577 34.46 91.609 34.524 ;
			RECT	91.745 34.46 91.777 34.524 ;
			RECT	91.913 34.46 91.945 34.524 ;
			RECT	92.081 34.46 92.113 34.524 ;
			RECT	92.249 34.46 92.281 34.524 ;
			RECT	92.417 34.46 92.449 34.524 ;
			RECT	92.585 34.46 92.617 34.524 ;
			RECT	92.753 34.46 92.785 34.524 ;
			RECT	92.921 34.46 92.953 34.524 ;
			RECT	93.089 34.46 93.121 34.524 ;
			RECT	93.257 34.46 93.289 34.524 ;
			RECT	93.425 34.46 93.457 34.524 ;
			RECT	93.593 34.46 93.625 34.524 ;
			RECT	93.761 34.46 93.793 34.524 ;
			RECT	93.929 34.46 93.961 34.524 ;
			RECT	94.097 34.46 94.129 34.524 ;
			RECT	94.265 34.46 94.297 34.524 ;
			RECT	94.433 34.46 94.465 34.524 ;
			RECT	94.601 34.46 94.633 34.524 ;
			RECT	94.769 34.46 94.801 34.524 ;
			RECT	94.937 34.46 94.969 34.524 ;
			RECT	95.105 34.46 95.137 34.524 ;
			RECT	95.273 34.46 95.305 34.524 ;
			RECT	95.441 34.46 95.473 34.524 ;
			RECT	95.609 34.46 95.641 34.524 ;
			RECT	95.777 34.46 95.809 34.524 ;
			RECT	95.945 34.46 95.977 34.524 ;
			RECT	96.113 34.46 96.145 34.524 ;
			RECT	96.281 34.46 96.313 34.524 ;
			RECT	96.449 34.46 96.481 34.524 ;
			RECT	96.617 34.46 96.649 34.524 ;
			RECT	96.785 34.46 96.817 34.524 ;
			RECT	96.953 34.46 96.985 34.524 ;
			RECT	97.121 34.46 97.153 34.524 ;
			RECT	97.289 34.46 97.321 34.524 ;
			RECT	97.457 34.46 97.489 34.524 ;
			RECT	97.625 34.46 97.657 34.524 ;
			RECT	97.793 34.46 97.825 34.524 ;
			RECT	97.961 34.46 97.993 34.524 ;
			RECT	98.129 34.46 98.161 34.524 ;
			RECT	98.297 34.46 98.329 34.524 ;
			RECT	98.465 34.46 98.497 34.524 ;
			RECT	98.633 34.46 98.665 34.524 ;
			RECT	98.801 34.46 98.833 34.524 ;
			RECT	98.969 34.46 99.001 34.524 ;
			RECT	99.137 34.46 99.169 34.524 ;
			RECT	99.305 34.46 99.337 34.524 ;
			RECT	99.473 34.46 99.505 34.524 ;
			RECT	99.641 34.46 99.673 34.524 ;
			RECT	99.809 34.46 99.841 34.524 ;
			RECT	99.977 34.46 100.009 34.524 ;
			RECT	100.145 34.46 100.177 34.524 ;
			RECT	100.313 34.46 100.345 34.524 ;
			RECT	100.481 34.46 100.513 34.524 ;
			RECT	100.649 34.46 100.681 34.524 ;
			RECT	100.817 34.46 100.849 34.524 ;
			RECT	100.985 34.46 101.017 34.524 ;
			RECT	101.153 34.46 101.185 34.524 ;
			RECT	101.321 34.46 101.353 34.524 ;
			RECT	101.489 34.46 101.521 34.524 ;
			RECT	101.657 34.46 101.689 34.524 ;
			RECT	101.825 34.46 101.857 34.524 ;
			RECT	101.993 34.46 102.025 34.524 ;
			RECT	104.177 34.46 104.209 34.524 ;
			RECT	104.345 34.46 104.377 34.524 ;
			RECT	104.513 34.46 104.545 34.524 ;
			RECT	104.681 34.46 104.713 34.524 ;
			RECT	104.849 34.46 104.881 34.524 ;
			RECT	105.017 34.46 105.049 34.524 ;
			RECT	105.185 34.46 105.217 34.524 ;
			RECT	105.353 34.46 105.385 34.524 ;
			RECT	105.521 34.46 105.553 34.524 ;
			RECT	105.689 34.46 105.721 34.524 ;
			RECT	105.857 34.46 105.889 34.524 ;
			RECT	106.025 34.46 106.057 34.524 ;
			RECT	106.193 34.46 106.225 34.524 ;
			RECT	106.361 34.46 106.393 34.524 ;
			RECT	106.529 34.46 106.561 34.524 ;
			RECT	106.697 34.46 106.729 34.524 ;
			RECT	106.865 34.46 106.897 34.524 ;
			RECT	107.033 34.46 107.065 34.524 ;
			RECT	107.201 34.46 107.233 34.524 ;
			RECT	107.369 34.46 107.401 34.524 ;
			RECT	107.537 34.46 107.569 34.524 ;
			RECT	107.705 34.46 107.737 34.524 ;
			RECT	107.873 34.46 107.905 34.524 ;
			RECT	108.041 34.46 108.073 34.524 ;
			RECT	108.209 34.46 108.241 34.524 ;
			RECT	108.377 34.46 108.409 34.524 ;
			RECT	108.545 34.46 108.577 34.524 ;
			RECT	108.713 34.46 108.745 34.524 ;
			RECT	108.881 34.46 108.913 34.524 ;
			RECT	109.049 34.46 109.081 34.524 ;
			RECT	109.217 34.46 109.249 34.524 ;
			RECT	109.385 34.46 109.417 34.524 ;
			RECT	109.553 34.46 109.585 34.524 ;
			RECT	109.721 34.46 109.753 34.524 ;
			RECT	109.889 34.46 109.921 34.524 ;
			RECT	110.057 34.46 110.089 34.524 ;
			RECT	110.225 34.46 110.257 34.524 ;
			RECT	110.393 34.46 110.425 34.524 ;
			RECT	110.561 34.46 110.593 34.524 ;
			RECT	110.729 34.46 110.761 34.524 ;
			RECT	110.897 34.46 110.929 34.524 ;
			RECT	111.065 34.46 111.097 34.524 ;
			RECT	111.233 34.46 111.265 34.524 ;
			RECT	111.401 34.46 111.433 34.524 ;
			RECT	111.569 34.46 111.601 34.524 ;
			RECT	111.737 34.46 111.769 34.524 ;
			RECT	111.905 34.46 111.937 34.524 ;
			RECT	112.073 34.46 112.105 34.524 ;
			RECT	112.241 34.46 112.273 34.524 ;
			RECT	112.409 34.46 112.441 34.524 ;
			RECT	112.577 34.46 112.609 34.524 ;
			RECT	112.745 34.46 112.777 34.524 ;
			RECT	112.913 34.46 112.945 34.524 ;
			RECT	113.081 34.46 113.113 34.524 ;
			RECT	113.249 34.46 113.281 34.524 ;
			RECT	113.417 34.46 113.449 34.524 ;
			RECT	113.585 34.46 113.617 34.524 ;
			RECT	113.753 34.46 113.785 34.524 ;
			RECT	113.921 34.46 113.953 34.524 ;
			RECT	114.089 34.46 114.121 34.524 ;
			RECT	114.257 34.46 114.289 34.524 ;
			RECT	114.425 34.46 114.457 34.524 ;
			RECT	114.593 34.46 114.625 34.524 ;
			RECT	114.761 34.46 114.793 34.524 ;
			RECT	114.929 34.46 114.961 34.524 ;
			RECT	115.097 34.46 115.129 34.524 ;
			RECT	115.265 34.46 115.297 34.524 ;
			RECT	115.433 34.46 115.465 34.524 ;
			RECT	115.601 34.46 115.633 34.524 ;
			RECT	115.769 34.46 115.801 34.524 ;
			RECT	115.937 34.46 115.969 34.524 ;
			RECT	116.105 34.46 116.137 34.524 ;
			RECT	116.273 34.46 116.305 34.524 ;
			RECT	116.441 34.46 116.473 34.524 ;
			RECT	116.609 34.46 116.641 34.524 ;
			RECT	116.777 34.46 116.809 34.524 ;
			RECT	116.945 34.46 116.977 34.524 ;
			RECT	117.113 34.46 117.145 34.524 ;
			RECT	117.281 34.46 117.313 34.524 ;
			RECT	117.449 34.46 117.481 34.524 ;
			RECT	117.617 34.46 117.649 34.524 ;
			RECT	117.785 34.46 117.817 34.524 ;
			RECT	117.953 34.46 117.985 34.524 ;
			RECT	118.121 34.46 118.153 34.524 ;
			RECT	118.289 34.46 118.321 34.524 ;
			RECT	118.457 34.46 118.489 34.524 ;
			RECT	118.625 34.46 118.657 34.524 ;
			RECT	118.793 34.46 118.825 34.524 ;
			RECT	118.961 34.46 118.993 34.524 ;
			RECT	119.129 34.46 119.161 34.524 ;
			RECT	119.297 34.46 119.329 34.524 ;
			RECT	119.465 34.46 119.497 34.524 ;
			RECT	119.633 34.46 119.665 34.524 ;
			RECT	119.801 34.46 119.833 34.524 ;
			RECT	119.969 34.46 120.001 34.524 ;
			RECT	120.137 34.46 120.169 34.524 ;
			RECT	120.305 34.46 120.337 34.524 ;
			RECT	120.473 34.46 120.505 34.524 ;
			RECT	120.641 34.46 120.673 34.524 ;
			RECT	120.809 34.46 120.841 34.524 ;
			RECT	120.977 34.46 121.009 34.524 ;
			RECT	121.145 34.46 121.177 34.524 ;
			RECT	121.313 34.46 121.345 34.524 ;
			RECT	121.481 34.46 121.513 34.524 ;
			RECT	121.649 34.46 121.681 34.524 ;
			RECT	121.817 34.46 121.849 34.524 ;
			RECT	121.985 34.46 122.017 34.524 ;
			RECT	122.153 34.46 122.185 34.524 ;
			RECT	122.321 34.46 122.353 34.524 ;
			RECT	122.489 34.46 122.521 34.524 ;
			RECT	122.657 34.46 122.689 34.524 ;
			RECT	122.825 34.46 122.857 34.524 ;
			RECT	122.993 34.46 123.025 34.524 ;
			RECT	123.161 34.46 123.193 34.524 ;
			RECT	123.329 34.46 123.361 34.524 ;
			RECT	123.497 34.46 123.529 34.524 ;
			RECT	123.665 34.46 123.697 34.524 ;
			RECT	123.833 34.46 123.865 34.524 ;
			RECT	124.001 34.46 124.033 34.524 ;
			RECT	124.169 34.46 124.201 34.524 ;
			RECT	124.337 34.46 124.369 34.524 ;
			RECT	124.505 34.46 124.537 34.524 ;
			RECT	124.673 34.46 124.705 34.524 ;
			RECT	124.841 34.46 124.873 34.524 ;
			RECT	125.009 34.46 125.041 34.524 ;
			RECT	125.177 34.46 125.209 34.524 ;
			RECT	125.345 34.46 125.377 34.524 ;
			RECT	125.513 34.46 125.545 34.524 ;
			RECT	125.681 34.46 125.713 34.524 ;
			RECT	125.849 34.46 125.881 34.524 ;
			RECT	126.017 34.46 126.049 34.524 ;
			RECT	126.185 34.46 126.217 34.524 ;
			RECT	126.353 34.46 126.385 34.524 ;
			RECT	126.521 34.46 126.553 34.524 ;
			RECT	126.689 34.46 126.721 34.524 ;
			RECT	126.857 34.46 126.889 34.524 ;
			RECT	127.025 34.46 127.057 34.524 ;
			RECT	127.193 34.46 127.225 34.524 ;
			RECT	127.361 34.46 127.393 34.524 ;
			RECT	127.529 34.46 127.561 34.524 ;
			RECT	127.697 34.46 127.729 34.524 ;
			RECT	127.865 34.46 127.897 34.524 ;
			RECT	128.033 34.46 128.065 34.524 ;
			RECT	128.201 34.46 128.233 34.524 ;
			RECT	128.369 34.46 128.401 34.524 ;
			RECT	128.537 34.46 128.569 34.524 ;
			RECT	128.705 34.46 128.737 34.524 ;
			RECT	128.873 34.46 128.905 34.524 ;
			RECT	129.041 34.46 129.073 34.524 ;
			RECT	129.209 34.46 129.241 34.524 ;
			RECT	129.377 34.46 129.409 34.524 ;
			RECT	129.545 34.46 129.577 34.524 ;
			RECT	129.713 34.46 129.745 34.524 ;
			RECT	129.881 34.46 129.913 34.524 ;
			RECT	130.049 34.46 130.081 34.524 ;
			RECT	130.217 34.46 130.249 34.524 ;
			RECT	130.385 34.46 130.417 34.524 ;
			RECT	130.553 34.46 130.585 34.524 ;
			RECT	130.721 34.46 130.753 34.524 ;
			RECT	130.889 34.46 130.921 34.524 ;
			RECT	131.057 34.46 131.089 34.524 ;
			RECT	131.225 34.46 131.257 34.524 ;
			RECT	131.393 34.46 131.425 34.524 ;
			RECT	131.561 34.46 131.593 34.524 ;
			RECT	131.729 34.46 131.761 34.524 ;
			RECT	131.897 34.46 131.929 34.524 ;
			RECT	132.065 34.46 132.097 34.524 ;
			RECT	132.233 34.46 132.265 34.524 ;
			RECT	132.401 34.46 132.433 34.524 ;
			RECT	132.569 34.46 132.601 34.524 ;
			RECT	132.737 34.46 132.769 34.524 ;
			RECT	132.905 34.46 132.937 34.524 ;
			RECT	133.073 34.46 133.105 34.524 ;
			RECT	133.241 34.46 133.273 34.524 ;
			RECT	133.409 34.46 133.441 34.524 ;
			RECT	133.577 34.46 133.609 34.524 ;
			RECT	133.745 34.46 133.777 34.524 ;
			RECT	133.913 34.46 133.945 34.524 ;
			RECT	134.081 34.46 134.113 34.524 ;
			RECT	134.249 34.46 134.281 34.524 ;
			RECT	134.417 34.46 134.449 34.524 ;
			RECT	134.585 34.46 134.617 34.524 ;
			RECT	134.753 34.46 134.785 34.524 ;
			RECT	134.921 34.46 134.953 34.524 ;
			RECT	135.089 34.46 135.121 34.524 ;
			RECT	135.257 34.46 135.289 34.524 ;
			RECT	135.425 34.46 135.457 34.524 ;
			RECT	135.593 34.46 135.625 34.524 ;
			RECT	135.761 34.46 135.793 34.524 ;
			RECT	135.929 34.46 135.961 34.524 ;
			RECT	136.097 34.46 136.129 34.524 ;
			RECT	136.265 34.46 136.297 34.524 ;
			RECT	136.433 34.46 136.465 34.524 ;
			RECT	136.601 34.46 136.633 34.524 ;
			RECT	136.769 34.46 136.801 34.524 ;
			RECT	136.937 34.46 136.969 34.524 ;
			RECT	137.105 34.46 137.137 34.524 ;
			RECT	137.273 34.46 137.305 34.524 ;
			RECT	137.441 34.46 137.473 34.524 ;
			RECT	137.609 34.46 137.641 34.524 ;
			RECT	137.777 34.46 137.809 34.524 ;
			RECT	137.945 34.46 137.977 34.524 ;
			RECT	138.113 34.46 138.145 34.524 ;
			RECT	138.281 34.46 138.313 34.524 ;
			RECT	138.449 34.46 138.481 34.524 ;
			RECT	138.617 34.46 138.649 34.524 ;
			RECT	138.785 34.46 138.817 34.524 ;
			RECT	138.953 34.46 138.985 34.524 ;
			RECT	139.121 34.46 139.153 34.524 ;
			RECT	139.289 34.46 139.321 34.524 ;
			RECT	139.457 34.46 139.489 34.524 ;
			RECT	139.625 34.46 139.657 34.524 ;
			RECT	139.793 34.46 139.825 34.524 ;
			RECT	139.961 34.46 139.993 34.524 ;
			RECT	140.129 34.46 140.161 34.524 ;
			RECT	140.297 34.46 140.329 34.524 ;
			RECT	140.465 34.46 140.497 34.524 ;
			RECT	140.633 34.46 140.665 34.524 ;
			RECT	140.801 34.46 140.833 34.524 ;
			RECT	140.969 34.46 141.001 34.524 ;
			RECT	141.137 34.46 141.169 34.524 ;
			RECT	141.305 34.46 141.337 34.524 ;
			RECT	141.473 34.46 141.505 34.524 ;
			RECT	141.641 34.46 141.673 34.524 ;
			RECT	141.809 34.46 141.841 34.524 ;
			RECT	141.977 34.46 142.009 34.524 ;
			RECT	142.145 34.46 142.177 34.524 ;
			RECT	142.313 34.46 142.345 34.524 ;
			RECT	142.481 34.46 142.513 34.524 ;
			RECT	142.649 34.46 142.681 34.524 ;
			RECT	142.817 34.46 142.849 34.524 ;
			RECT	142.985 34.46 143.017 34.524 ;
			RECT	143.153 34.46 143.185 34.524 ;
			RECT	143.321 34.46 143.353 34.524 ;
			RECT	143.489 34.46 143.521 34.524 ;
			RECT	143.657 34.46 143.689 34.524 ;
			RECT	143.825 34.46 143.857 34.524 ;
			RECT	143.993 34.46 144.025 34.524 ;
			RECT	144.161 34.46 144.193 34.524 ;
			RECT	144.329 34.46 144.361 34.524 ;
			RECT	144.497 34.46 144.529 34.524 ;
			RECT	144.665 34.46 144.697 34.524 ;
			RECT	144.833 34.46 144.865 34.524 ;
			RECT	145.001 34.46 145.033 34.524 ;
			RECT	145.169 34.46 145.201 34.524 ;
			RECT	145.337 34.46 145.369 34.524 ;
			RECT	145.505 34.46 145.537 34.524 ;
			RECT	145.673 34.46 145.705 34.524 ;
			RECT	145.841 34.46 145.873 34.524 ;
			RECT	146.009 34.46 146.041 34.524 ;
			RECT	146.177 34.46 146.209 34.524 ;
			RECT	146.345 34.46 146.377 34.524 ;
			RECT	146.513 34.46 146.545 34.524 ;
			RECT	146.681 34.46 146.713 34.524 ;
			RECT	146.849 34.46 146.881 34.524 ;
			RECT	147.017 34.46 147.049 34.524 ;
			RECT	147.185 34.46 147.217 34.524 ;
			RECT	147.309 34.46 147.373 34.524 ;
			RECT	147.611 34.46 147.643 34.524 ;
			RECT	149.918 34.46 149.95 34.524 ;
			RECT	150.219 34.46 150.251 34.524 ;
			RECT	150.966 34.46 151.03 34.524 ;
			RECT	151.908 34.46 151.94 34.524 ;
			RECT	153.967 34.46 154.031 34.524 ;
			RECT	156.557 34.46 156.589 34.524 ;
			RECT	156.827 34.46 156.891 34.524 ;
			RECT	156.983 34.46 157.015 34.524 ;
			RECT	157.151 34.46 157.183 34.524 ;
			RECT	157.319 34.46 157.351 34.524 ;
			RECT	157.487 34.46 157.519 34.524 ;
			RECT	157.655 34.46 157.687 34.524 ;
			RECT	157.823 34.46 157.855 34.524 ;
			RECT	157.991 34.46 158.023 34.524 ;
			RECT	158.159 34.46 158.191 34.524 ;
			RECT	158.327 34.46 158.359 34.524 ;
			RECT	158.495 34.46 158.527 34.524 ;
			RECT	158.663 34.46 158.695 34.524 ;
			RECT	158.831 34.46 158.863 34.524 ;
			RECT	158.999 34.46 159.031 34.524 ;
			RECT	159.167 34.46 159.199 34.524 ;
			RECT	159.335 34.46 159.367 34.524 ;
			RECT	159.503 34.46 159.535 34.524 ;
			RECT	159.671 34.46 159.703 34.524 ;
			RECT	159.839 34.46 159.871 34.524 ;
			RECT	160.007 34.46 160.039 34.524 ;
			RECT	160.175 34.46 160.207 34.524 ;
			RECT	160.343 34.46 160.375 34.524 ;
			RECT	160.511 34.46 160.543 34.524 ;
			RECT	160.679 34.46 160.711 34.524 ;
			RECT	160.847 34.46 160.879 34.524 ;
			RECT	161.015 34.46 161.047 34.524 ;
			RECT	161.183 34.46 161.215 34.524 ;
			RECT	161.351 34.46 161.383 34.524 ;
			RECT	161.519 34.46 161.551 34.524 ;
			RECT	161.687 34.46 161.719 34.524 ;
			RECT	161.855 34.46 161.887 34.524 ;
			RECT	162.023 34.46 162.055 34.524 ;
			RECT	162.191 34.46 162.223 34.524 ;
			RECT	162.359 34.46 162.391 34.524 ;
			RECT	162.527 34.46 162.559 34.524 ;
			RECT	162.695 34.46 162.727 34.524 ;
			RECT	162.863 34.46 162.895 34.524 ;
			RECT	163.031 34.46 163.063 34.524 ;
			RECT	163.199 34.46 163.231 34.524 ;
			RECT	163.367 34.46 163.399 34.524 ;
			RECT	163.535 34.46 163.567 34.524 ;
			RECT	163.703 34.46 163.735 34.524 ;
			RECT	163.871 34.46 163.903 34.524 ;
			RECT	164.039 34.46 164.071 34.524 ;
			RECT	164.207 34.46 164.239 34.524 ;
			RECT	164.375 34.46 164.407 34.524 ;
			RECT	164.543 34.46 164.575 34.524 ;
			RECT	164.711 34.46 164.743 34.524 ;
			RECT	164.879 34.46 164.911 34.524 ;
			RECT	165.047 34.46 165.079 34.524 ;
			RECT	165.215 34.46 165.247 34.524 ;
			RECT	165.383 34.46 165.415 34.524 ;
			RECT	165.551 34.46 165.583 34.524 ;
			RECT	165.719 34.46 165.751 34.524 ;
			RECT	165.887 34.46 165.919 34.524 ;
			RECT	166.055 34.46 166.087 34.524 ;
			RECT	166.223 34.46 166.255 34.524 ;
			RECT	166.391 34.46 166.423 34.524 ;
			RECT	166.559 34.46 166.591 34.524 ;
			RECT	166.727 34.46 166.759 34.524 ;
			RECT	166.895 34.46 166.927 34.524 ;
			RECT	167.063 34.46 167.095 34.524 ;
			RECT	167.231 34.46 167.263 34.524 ;
			RECT	167.399 34.46 167.431 34.524 ;
			RECT	167.567 34.46 167.599 34.524 ;
			RECT	167.735 34.46 167.767 34.524 ;
			RECT	167.903 34.46 167.935 34.524 ;
			RECT	168.071 34.46 168.103 34.524 ;
			RECT	168.239 34.46 168.271 34.524 ;
			RECT	168.407 34.46 168.439 34.524 ;
			RECT	168.575 34.46 168.607 34.524 ;
			RECT	168.743 34.46 168.775 34.524 ;
			RECT	168.911 34.46 168.943 34.524 ;
			RECT	169.079 34.46 169.111 34.524 ;
			RECT	169.247 34.46 169.279 34.524 ;
			RECT	169.415 34.46 169.447 34.524 ;
			RECT	169.583 34.46 169.615 34.524 ;
			RECT	169.751 34.46 169.783 34.524 ;
			RECT	169.919 34.46 169.951 34.524 ;
			RECT	170.087 34.46 170.119 34.524 ;
			RECT	170.255 34.46 170.287 34.524 ;
			RECT	170.423 34.46 170.455 34.524 ;
			RECT	170.591 34.46 170.623 34.524 ;
			RECT	170.759 34.46 170.791 34.524 ;
			RECT	170.927 34.46 170.959 34.524 ;
			RECT	171.095 34.46 171.127 34.524 ;
			RECT	171.263 34.46 171.295 34.524 ;
			RECT	171.431 34.46 171.463 34.524 ;
			RECT	171.599 34.46 171.631 34.524 ;
			RECT	171.767 34.46 171.799 34.524 ;
			RECT	171.935 34.46 171.967 34.524 ;
			RECT	172.103 34.46 172.135 34.524 ;
			RECT	172.271 34.46 172.303 34.524 ;
			RECT	172.439 34.46 172.471 34.524 ;
			RECT	172.607 34.46 172.639 34.524 ;
			RECT	172.775 34.46 172.807 34.524 ;
			RECT	172.943 34.46 172.975 34.524 ;
			RECT	173.111 34.46 173.143 34.524 ;
			RECT	173.279 34.46 173.311 34.524 ;
			RECT	173.447 34.46 173.479 34.524 ;
			RECT	173.615 34.46 173.647 34.524 ;
			RECT	173.783 34.46 173.815 34.524 ;
			RECT	173.951 34.46 173.983 34.524 ;
			RECT	174.119 34.46 174.151 34.524 ;
			RECT	174.287 34.46 174.319 34.524 ;
			RECT	174.455 34.46 174.487 34.524 ;
			RECT	174.623 34.46 174.655 34.524 ;
			RECT	174.791 34.46 174.823 34.524 ;
			RECT	174.959 34.46 174.991 34.524 ;
			RECT	175.127 34.46 175.159 34.524 ;
			RECT	175.295 34.46 175.327 34.524 ;
			RECT	175.463 34.46 175.495 34.524 ;
			RECT	175.631 34.46 175.663 34.524 ;
			RECT	175.799 34.46 175.831 34.524 ;
			RECT	175.967 34.46 175.999 34.524 ;
			RECT	176.135 34.46 176.167 34.524 ;
			RECT	176.303 34.46 176.335 34.524 ;
			RECT	176.471 34.46 176.503 34.524 ;
			RECT	176.639 34.46 176.671 34.524 ;
			RECT	176.807 34.46 176.839 34.524 ;
			RECT	176.975 34.46 177.007 34.524 ;
			RECT	177.143 34.46 177.175 34.524 ;
			RECT	177.311 34.46 177.343 34.524 ;
			RECT	177.479 34.46 177.511 34.524 ;
			RECT	177.647 34.46 177.679 34.524 ;
			RECT	177.815 34.46 177.847 34.524 ;
			RECT	177.983 34.46 178.015 34.524 ;
			RECT	178.151 34.46 178.183 34.524 ;
			RECT	178.319 34.46 178.351 34.524 ;
			RECT	178.487 34.46 178.519 34.524 ;
			RECT	178.655 34.46 178.687 34.524 ;
			RECT	178.823 34.46 178.855 34.524 ;
			RECT	178.991 34.46 179.023 34.524 ;
			RECT	179.159 34.46 179.191 34.524 ;
			RECT	179.327 34.46 179.359 34.524 ;
			RECT	179.495 34.46 179.527 34.524 ;
			RECT	179.663 34.46 179.695 34.524 ;
			RECT	179.831 34.46 179.863 34.524 ;
			RECT	179.999 34.46 180.031 34.524 ;
			RECT	180.167 34.46 180.199 34.524 ;
			RECT	180.335 34.46 180.367 34.524 ;
			RECT	180.503 34.46 180.535 34.524 ;
			RECT	180.671 34.46 180.703 34.524 ;
			RECT	180.839 34.46 180.871 34.524 ;
			RECT	181.007 34.46 181.039 34.524 ;
			RECT	181.175 34.46 181.207 34.524 ;
			RECT	181.343 34.46 181.375 34.524 ;
			RECT	181.511 34.46 181.543 34.524 ;
			RECT	181.679 34.46 181.711 34.524 ;
			RECT	181.847 34.46 181.879 34.524 ;
			RECT	182.015 34.46 182.047 34.524 ;
			RECT	182.183 34.46 182.215 34.524 ;
			RECT	182.351 34.46 182.383 34.524 ;
			RECT	182.519 34.46 182.551 34.524 ;
			RECT	182.687 34.46 182.719 34.524 ;
			RECT	182.855 34.46 182.887 34.524 ;
			RECT	183.023 34.46 183.055 34.524 ;
			RECT	183.191 34.46 183.223 34.524 ;
			RECT	183.359 34.46 183.391 34.524 ;
			RECT	183.527 34.46 183.559 34.524 ;
			RECT	183.695 34.46 183.727 34.524 ;
			RECT	183.863 34.46 183.895 34.524 ;
			RECT	184.031 34.46 184.063 34.524 ;
			RECT	184.199 34.46 184.231 34.524 ;
			RECT	184.367 34.46 184.399 34.524 ;
			RECT	184.535 34.46 184.567 34.524 ;
			RECT	184.703 34.46 184.735 34.524 ;
			RECT	184.871 34.46 184.903 34.524 ;
			RECT	185.039 34.46 185.071 34.524 ;
			RECT	185.207 34.46 185.239 34.524 ;
			RECT	185.375 34.46 185.407 34.524 ;
			RECT	185.543 34.46 185.575 34.524 ;
			RECT	185.711 34.46 185.743 34.524 ;
			RECT	185.879 34.46 185.911 34.524 ;
			RECT	186.047 34.46 186.079 34.524 ;
			RECT	186.215 34.46 186.247 34.524 ;
			RECT	186.383 34.46 186.415 34.524 ;
			RECT	186.551 34.46 186.583 34.524 ;
			RECT	186.719 34.46 186.751 34.524 ;
			RECT	186.887 34.46 186.919 34.524 ;
			RECT	187.055 34.46 187.087 34.524 ;
			RECT	187.223 34.46 187.255 34.524 ;
			RECT	187.391 34.46 187.423 34.524 ;
			RECT	187.559 34.46 187.591 34.524 ;
			RECT	187.727 34.46 187.759 34.524 ;
			RECT	187.895 34.46 187.927 34.524 ;
			RECT	188.063 34.46 188.095 34.524 ;
			RECT	188.231 34.46 188.263 34.524 ;
			RECT	188.399 34.46 188.431 34.524 ;
			RECT	188.567 34.46 188.599 34.524 ;
			RECT	188.735 34.46 188.767 34.524 ;
			RECT	188.903 34.46 188.935 34.524 ;
			RECT	189.071 34.46 189.103 34.524 ;
			RECT	189.239 34.46 189.271 34.524 ;
			RECT	189.407 34.46 189.439 34.524 ;
			RECT	189.575 34.46 189.607 34.524 ;
			RECT	189.743 34.46 189.775 34.524 ;
			RECT	189.911 34.46 189.943 34.524 ;
			RECT	190.079 34.46 190.111 34.524 ;
			RECT	190.247 34.46 190.279 34.524 ;
			RECT	190.415 34.46 190.447 34.524 ;
			RECT	190.583 34.46 190.615 34.524 ;
			RECT	190.751 34.46 190.783 34.524 ;
			RECT	190.919 34.46 190.951 34.524 ;
			RECT	191.087 34.46 191.119 34.524 ;
			RECT	191.255 34.46 191.287 34.524 ;
			RECT	191.423 34.46 191.455 34.524 ;
			RECT	191.591 34.46 191.623 34.524 ;
			RECT	191.759 34.46 191.791 34.524 ;
			RECT	191.927 34.46 191.959 34.524 ;
			RECT	192.095 34.46 192.127 34.524 ;
			RECT	192.263 34.46 192.295 34.524 ;
			RECT	192.431 34.46 192.463 34.524 ;
			RECT	192.599 34.46 192.631 34.524 ;
			RECT	192.767 34.46 192.799 34.524 ;
			RECT	192.935 34.46 192.967 34.524 ;
			RECT	193.103 34.46 193.135 34.524 ;
			RECT	193.271 34.46 193.303 34.524 ;
			RECT	193.439 34.46 193.471 34.524 ;
			RECT	193.607 34.46 193.639 34.524 ;
			RECT	193.775 34.46 193.807 34.524 ;
			RECT	193.943 34.46 193.975 34.524 ;
			RECT	194.111 34.46 194.143 34.524 ;
			RECT	194.279 34.46 194.311 34.524 ;
			RECT	194.447 34.46 194.479 34.524 ;
			RECT	194.615 34.46 194.647 34.524 ;
			RECT	194.783 34.46 194.815 34.524 ;
			RECT	194.951 34.46 194.983 34.524 ;
			RECT	195.119 34.46 195.151 34.524 ;
			RECT	195.287 34.46 195.319 34.524 ;
			RECT	195.455 34.46 195.487 34.524 ;
			RECT	195.623 34.46 195.655 34.524 ;
			RECT	195.791 34.46 195.823 34.524 ;
			RECT	195.959 34.46 195.991 34.524 ;
			RECT	196.127 34.46 196.159 34.524 ;
			RECT	196.295 34.46 196.327 34.524 ;
			RECT	196.463 34.46 196.495 34.524 ;
			RECT	196.631 34.46 196.663 34.524 ;
			RECT	196.799 34.46 196.831 34.524 ;
			RECT	196.967 34.46 196.999 34.524 ;
			RECT	197.135 34.46 197.167 34.524 ;
			RECT	197.303 34.46 197.335 34.524 ;
			RECT	197.471 34.46 197.503 34.524 ;
			RECT	197.639 34.46 197.671 34.524 ;
			RECT	197.807 34.46 197.839 34.524 ;
			RECT	197.975 34.46 198.007 34.524 ;
			RECT	198.143 34.46 198.175 34.524 ;
			RECT	198.311 34.46 198.343 34.524 ;
			RECT	198.479 34.46 198.511 34.524 ;
			RECT	198.647 34.46 198.679 34.524 ;
			RECT	198.815 34.46 198.847 34.524 ;
			RECT	198.983 34.46 199.015 34.524 ;
			RECT	199.151 34.46 199.183 34.524 ;
			RECT	199.319 34.46 199.351 34.524 ;
			RECT	199.487 34.46 199.519 34.524 ;
			RECT	199.655 34.46 199.687 34.524 ;
			RECT	199.823 34.46 199.855 34.524 ;
			RECT	199.991 34.46 200.023 34.524 ;
			RECT	200.9 34.46 200.932 34.524 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 35.567 201.665 35.657 ;
			LAYER	J3 ;
			RECT	1.645 35.596 1.709 35.628 ;
			RECT	2.323 35.596 2.387 35.628 ;
			RECT	2.957 35.58 2.989 35.644 ;
			RECT	3.438 35.58 3.47 35.644 ;
			RECT	4.138 35.596 4.202 35.628 ;
			RECT	4.354 35.58 4.386 35.644 ;
			RECT	5.252 35.58 5.284 35.644 ;
			RECT	5.758 35.58 5.79 35.644 ;
			RECT	49.311 35.596 49.375 35.628 ;
			RECT	49.613 35.58 49.645 35.644 ;
			RECT	51.92 35.58 51.952 35.644 ;
			RECT	52.968 35.596 53.032 35.628 ;
			RECT	53.91 35.58 53.942 35.644 ;
			RECT	55.969 35.596 56.033 35.628 ;
			RECT	58.559 35.58 58.591 35.644 ;
			RECT	58.829 35.596 58.893 35.628 ;
			RECT	102.414 35.58 102.446 35.644 ;
			RECT	103.756 35.58 103.788 35.644 ;
			RECT	147.309 35.596 147.373 35.628 ;
			RECT	147.611 35.58 147.643 35.644 ;
			RECT	149.918 35.58 149.95 35.644 ;
			RECT	150.966 35.596 151.03 35.628 ;
			RECT	151.908 35.58 151.94 35.644 ;
			RECT	153.967 35.596 154.031 35.628 ;
			RECT	156.557 35.58 156.589 35.644 ;
			RECT	156.827 35.596 156.891 35.628 ;
			RECT	200.412 35.58 200.444 35.644 ;
			RECT	200.9 35.58 200.932 35.644 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 36.67 201.665 36.76 ;
			LAYER	J3 ;
			RECT	1.661 36.683 1.693 36.747 ;
			RECT	2.323 36.699 2.387 36.731 ;
			RECT	3.438 36.683 3.47 36.747 ;
			RECT	4.354 36.683 4.386 36.747 ;
			RECT	4.539 36.683 4.571 36.747 ;
			RECT	4.805 36.683 4.837 36.747 ;
			RECT	5.252 36.683 5.284 36.747 ;
			RECT	5.758 36.683 5.79 36.747 ;
			RECT	49.311 36.699 49.375 36.731 ;
			RECT	49.613 36.683 49.645 36.747 ;
			RECT	51.921 36.698 51.953 36.73 ;
			RECT	52.968 36.699 53.032 36.731 ;
			RECT	53.91 36.683 53.942 36.747 ;
			RECT	54.812 36.699 54.844 36.731 ;
			RECT	55.969 36.699 56.033 36.731 ;
			RECT	58.559 36.683 58.591 36.747 ;
			RECT	58.829 36.699 58.893 36.731 ;
			RECT	102.414 36.683 102.446 36.747 ;
			RECT	103.756 36.683 103.788 36.747 ;
			RECT	147.309 36.699 147.373 36.731 ;
			RECT	147.611 36.683 147.643 36.747 ;
			RECT	149.919 36.698 149.951 36.73 ;
			RECT	150.966 36.699 151.03 36.731 ;
			RECT	151.908 36.683 151.94 36.747 ;
			RECT	152.81 36.699 152.842 36.731 ;
			RECT	153.967 36.699 154.031 36.731 ;
			RECT	156.557 36.683 156.589 36.747 ;
			RECT	156.827 36.699 156.891 36.731 ;
			RECT	200.412 36.683 200.444 36.747 ;
			RECT	200.9 36.683 200.932 36.747 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 37.255 201.665 37.375 ;
			LAYER	J3 ;
			RECT	1.645 37.283 1.709 37.347 ;
			RECT	2.197 37.283 2.229 37.347 ;
			RECT	2.323 37.283 2.387 37.347 ;
			RECT	3.438 37.283 3.47 37.347 ;
			RECT	4.539 37.283 4.571 37.347 ;
			RECT	4.805 37.283 4.837 37.347 ;
			RECT	4.982 37.283 5.014 37.347 ;
			RECT	5.758 37.283 5.79 37.347 ;
			RECT	6.389 37.283 6.421 37.347 ;
			RECT	6.725 37.283 6.757 37.347 ;
			RECT	7.061 37.283 7.093 37.347 ;
			RECT	7.397 37.283 7.429 37.347 ;
			RECT	7.733 37.283 7.765 37.347 ;
			RECT	8.069 37.283 8.101 37.347 ;
			RECT	8.405 37.283 8.437 37.347 ;
			RECT	8.741 37.283 8.773 37.347 ;
			RECT	9.077 37.283 9.109 37.347 ;
			RECT	9.413 37.283 9.445 37.347 ;
			RECT	9.749 37.283 9.781 37.347 ;
			RECT	10.085 37.283 10.117 37.347 ;
			RECT	10.421 37.283 10.453 37.347 ;
			RECT	10.757 37.283 10.789 37.347 ;
			RECT	11.093 37.283 11.125 37.347 ;
			RECT	11.429 37.283 11.461 37.347 ;
			RECT	11.765 37.283 11.797 37.347 ;
			RECT	12.101 37.283 12.133 37.347 ;
			RECT	12.437 37.283 12.469 37.347 ;
			RECT	12.773 37.283 12.805 37.347 ;
			RECT	13.109 37.283 13.141 37.347 ;
			RECT	13.445 37.283 13.477 37.347 ;
			RECT	13.781 37.283 13.813 37.347 ;
			RECT	14.117 37.283 14.149 37.347 ;
			RECT	14.453 37.283 14.485 37.347 ;
			RECT	14.789 37.283 14.821 37.347 ;
			RECT	15.125 37.283 15.157 37.347 ;
			RECT	15.461 37.283 15.493 37.347 ;
			RECT	15.797 37.283 15.829 37.347 ;
			RECT	16.133 37.283 16.165 37.347 ;
			RECT	16.469 37.283 16.501 37.347 ;
			RECT	16.805 37.283 16.837 37.347 ;
			RECT	17.141 37.283 17.173 37.347 ;
			RECT	17.477 37.283 17.509 37.347 ;
			RECT	17.813 37.283 17.845 37.347 ;
			RECT	18.149 37.283 18.181 37.347 ;
			RECT	18.485 37.283 18.517 37.347 ;
			RECT	18.821 37.283 18.853 37.347 ;
			RECT	19.157 37.283 19.189 37.347 ;
			RECT	19.493 37.283 19.525 37.347 ;
			RECT	19.829 37.283 19.861 37.347 ;
			RECT	20.165 37.283 20.197 37.347 ;
			RECT	20.501 37.283 20.533 37.347 ;
			RECT	20.837 37.283 20.869 37.347 ;
			RECT	21.173 37.283 21.205 37.347 ;
			RECT	21.509 37.283 21.541 37.347 ;
			RECT	21.845 37.283 21.877 37.347 ;
			RECT	22.181 37.283 22.213 37.347 ;
			RECT	22.517 37.283 22.549 37.347 ;
			RECT	22.853 37.283 22.885 37.347 ;
			RECT	23.189 37.283 23.221 37.347 ;
			RECT	23.525 37.283 23.557 37.347 ;
			RECT	23.861 37.283 23.893 37.347 ;
			RECT	24.197 37.283 24.229 37.347 ;
			RECT	24.533 37.283 24.565 37.347 ;
			RECT	24.869 37.283 24.901 37.347 ;
			RECT	25.205 37.283 25.237 37.347 ;
			RECT	25.541 37.283 25.573 37.347 ;
			RECT	25.877 37.283 25.909 37.347 ;
			RECT	26.213 37.283 26.245 37.347 ;
			RECT	26.549 37.283 26.581 37.347 ;
			RECT	26.885 37.283 26.917 37.347 ;
			RECT	27.221 37.283 27.253 37.347 ;
			RECT	27.557 37.283 27.589 37.347 ;
			RECT	27.888 37.283 27.92 37.347 ;
			RECT	28.224 37.283 28.256 37.347 ;
			RECT	28.56 37.283 28.592 37.347 ;
			RECT	28.896 37.283 28.928 37.347 ;
			RECT	29.232 37.283 29.264 37.347 ;
			RECT	29.568 37.283 29.6 37.347 ;
			RECT	29.904 37.283 29.936 37.347 ;
			RECT	30.24 37.283 30.272 37.347 ;
			RECT	30.576 37.283 30.608 37.347 ;
			RECT	30.912 37.283 30.944 37.347 ;
			RECT	31.248 37.283 31.28 37.347 ;
			RECT	31.584 37.283 31.616 37.347 ;
			RECT	31.92 37.283 31.952 37.347 ;
			RECT	32.256 37.283 32.288 37.347 ;
			RECT	32.592 37.283 32.624 37.347 ;
			RECT	32.928 37.283 32.96 37.347 ;
			RECT	34.608 37.283 34.64 37.347 ;
			RECT	34.944 37.283 34.976 37.347 ;
			RECT	35.28 37.283 35.312 37.347 ;
			RECT	35.616 37.283 35.648 37.347 ;
			RECT	36.288 37.283 36.32 37.347 ;
			RECT	36.96 37.283 36.992 37.347 ;
			RECT	37.632 37.283 37.664 37.347 ;
			RECT	37.968 37.283 38 37.347 ;
			RECT	38.304 37.283 38.336 37.347 ;
			RECT	38.64 37.283 38.672 37.347 ;
			RECT	38.976 37.283 39.008 37.347 ;
			RECT	39.648 37.283 39.68 37.347 ;
			RECT	39.984 37.283 40.016 37.347 ;
			RECT	40.32 37.283 40.352 37.347 ;
			RECT	40.992 37.283 41.024 37.347 ;
			RECT	41.664 37.283 41.696 37.347 ;
			RECT	42 37.283 42.032 37.347 ;
			RECT	42.336 37.283 42.368 37.347 ;
			RECT	42.672 37.283 42.704 37.347 ;
			RECT	43.008 37.283 43.04 37.347 ;
			RECT	43.344 37.283 43.376 37.347 ;
			RECT	43.68 37.283 43.712 37.347 ;
			RECT	44.68 37.283 44.712 37.347 ;
			RECT	45.024 37.283 45.056 37.347 ;
			RECT	46.032 37.283 46.064 37.347 ;
			RECT	46.368 37.283 46.4 37.347 ;
			RECT	47.04 37.283 47.072 37.347 ;
			RECT	47.376 37.283 47.408 37.347 ;
			RECT	48.048 37.283 48.08 37.347 ;
			RECT	48.384 37.283 48.416 37.347 ;
			RECT	48.72 37.283 48.752 37.347 ;
			RECT	49.056 37.283 49.088 37.347 ;
			RECT	49.311 37.283 49.375 37.347 ;
			RECT	49.613 37.283 49.645 37.347 ;
			RECT	51.92 37.299 51.952 37.331 ;
			RECT	52.968 37.283 53.032 37.347 ;
			RECT	53.91 37.283 53.942 37.347 ;
			RECT	54.812 37.283 54.844 37.347 ;
			RECT	55.969 37.283 56.033 37.347 ;
			RECT	57.911 37.283 57.943 37.347 ;
			RECT	58.559 37.283 58.591 37.347 ;
			RECT	58.829 37.283 58.893 37.347 ;
			RECT	59.116 37.283 59.148 37.347 ;
			RECT	59.452 37.283 59.484 37.347 ;
			RECT	59.788 37.283 59.82 37.347 ;
			RECT	60.124 37.283 60.156 37.347 ;
			RECT	60.796 37.283 60.828 37.347 ;
			RECT	61.132 37.283 61.164 37.347 ;
			RECT	61.804 37.283 61.836 37.347 ;
			RECT	62.14 37.283 62.172 37.347 ;
			RECT	63.148 37.283 63.18 37.347 ;
			RECT	63.492 37.283 63.524 37.347 ;
			RECT	64.492 37.283 64.524 37.347 ;
			RECT	64.828 37.283 64.86 37.347 ;
			RECT	65.164 37.283 65.196 37.347 ;
			RECT	65.5 37.283 65.532 37.347 ;
			RECT	65.836 37.283 65.868 37.347 ;
			RECT	66.172 37.283 66.204 37.347 ;
			RECT	66.508 37.283 66.54 37.347 ;
			RECT	67.18 37.283 67.212 37.347 ;
			RECT	67.852 37.283 67.884 37.347 ;
			RECT	68.188 37.283 68.22 37.347 ;
			RECT	68.524 37.283 68.556 37.347 ;
			RECT	69.196 37.283 69.228 37.347 ;
			RECT	69.532 37.283 69.564 37.347 ;
			RECT	69.868 37.283 69.9 37.347 ;
			RECT	70.204 37.283 70.236 37.347 ;
			RECT	70.54 37.283 70.572 37.347 ;
			RECT	71.212 37.283 71.244 37.347 ;
			RECT	71.884 37.283 71.916 37.347 ;
			RECT	72.556 37.283 72.588 37.347 ;
			RECT	72.892 37.283 72.924 37.347 ;
			RECT	73.228 37.283 73.26 37.347 ;
			RECT	73.564 37.283 73.596 37.347 ;
			RECT	75.244 37.283 75.276 37.347 ;
			RECT	75.58 37.283 75.612 37.347 ;
			RECT	75.916 37.283 75.948 37.347 ;
			RECT	76.252 37.283 76.284 37.347 ;
			RECT	76.588 37.283 76.62 37.347 ;
			RECT	76.924 37.283 76.956 37.347 ;
			RECT	77.26 37.283 77.292 37.347 ;
			RECT	77.596 37.283 77.628 37.347 ;
			RECT	77.932 37.283 77.964 37.347 ;
			RECT	78.268 37.283 78.3 37.347 ;
			RECT	78.604 37.283 78.636 37.347 ;
			RECT	78.94 37.283 78.972 37.347 ;
			RECT	79.276 37.283 79.308 37.347 ;
			RECT	79.612 37.283 79.644 37.347 ;
			RECT	79.948 37.283 79.98 37.347 ;
			RECT	80.284 37.283 80.316 37.347 ;
			RECT	80.615 37.283 80.647 37.347 ;
			RECT	80.951 37.283 80.983 37.347 ;
			RECT	81.287 37.283 81.319 37.347 ;
			RECT	81.623 37.283 81.655 37.347 ;
			RECT	81.959 37.283 81.991 37.347 ;
			RECT	82.295 37.283 82.327 37.347 ;
			RECT	82.631 37.283 82.663 37.347 ;
			RECT	82.967 37.283 82.999 37.347 ;
			RECT	83.303 37.283 83.335 37.347 ;
			RECT	83.639 37.283 83.671 37.347 ;
			RECT	83.975 37.283 84.007 37.347 ;
			RECT	84.311 37.283 84.343 37.347 ;
			RECT	84.647 37.283 84.679 37.347 ;
			RECT	84.983 37.283 85.015 37.347 ;
			RECT	85.319 37.283 85.351 37.347 ;
			RECT	85.655 37.283 85.687 37.347 ;
			RECT	85.991 37.283 86.023 37.347 ;
			RECT	86.327 37.283 86.359 37.347 ;
			RECT	86.663 37.283 86.695 37.347 ;
			RECT	86.999 37.283 87.031 37.347 ;
			RECT	87.335 37.283 87.367 37.347 ;
			RECT	87.671 37.283 87.703 37.347 ;
			RECT	88.007 37.283 88.039 37.347 ;
			RECT	88.343 37.283 88.375 37.347 ;
			RECT	88.679 37.283 88.711 37.347 ;
			RECT	89.015 37.283 89.047 37.347 ;
			RECT	89.351 37.283 89.383 37.347 ;
			RECT	89.687 37.283 89.719 37.347 ;
			RECT	90.023 37.283 90.055 37.347 ;
			RECT	90.359 37.283 90.391 37.347 ;
			RECT	90.695 37.283 90.727 37.347 ;
			RECT	91.031 37.283 91.063 37.347 ;
			RECT	91.367 37.283 91.399 37.347 ;
			RECT	91.703 37.283 91.735 37.347 ;
			RECT	92.039 37.283 92.071 37.347 ;
			RECT	92.375 37.283 92.407 37.347 ;
			RECT	92.711 37.283 92.743 37.347 ;
			RECT	93.047 37.283 93.079 37.347 ;
			RECT	93.383 37.283 93.415 37.347 ;
			RECT	93.719 37.283 93.751 37.347 ;
			RECT	94.055 37.283 94.087 37.347 ;
			RECT	94.391 37.283 94.423 37.347 ;
			RECT	94.727 37.283 94.759 37.347 ;
			RECT	95.063 37.283 95.095 37.347 ;
			RECT	95.399 37.283 95.431 37.347 ;
			RECT	95.735 37.283 95.767 37.347 ;
			RECT	96.071 37.283 96.103 37.347 ;
			RECT	96.407 37.283 96.439 37.347 ;
			RECT	96.743 37.283 96.775 37.347 ;
			RECT	97.079 37.283 97.111 37.347 ;
			RECT	97.415 37.283 97.447 37.347 ;
			RECT	97.751 37.283 97.783 37.347 ;
			RECT	98.087 37.283 98.119 37.347 ;
			RECT	98.423 37.283 98.455 37.347 ;
			RECT	98.759 37.283 98.791 37.347 ;
			RECT	99.095 37.283 99.127 37.347 ;
			RECT	99.431 37.283 99.463 37.347 ;
			RECT	99.767 37.283 99.799 37.347 ;
			RECT	100.103 37.283 100.135 37.347 ;
			RECT	100.439 37.283 100.471 37.347 ;
			RECT	100.775 37.283 100.807 37.347 ;
			RECT	101.111 37.283 101.143 37.347 ;
			RECT	101.447 37.283 101.479 37.347 ;
			RECT	101.783 37.283 101.815 37.347 ;
			RECT	102.414 37.283 102.446 37.347 ;
			RECT	103.756 37.283 103.788 37.347 ;
			RECT	104.387 37.283 104.419 37.347 ;
			RECT	104.723 37.283 104.755 37.347 ;
			RECT	105.059 37.283 105.091 37.347 ;
			RECT	105.395 37.283 105.427 37.347 ;
			RECT	105.731 37.283 105.763 37.347 ;
			RECT	106.067 37.283 106.099 37.347 ;
			RECT	106.403 37.283 106.435 37.347 ;
			RECT	106.739 37.283 106.771 37.347 ;
			RECT	107.075 37.283 107.107 37.347 ;
			RECT	107.411 37.283 107.443 37.347 ;
			RECT	107.747 37.283 107.779 37.347 ;
			RECT	108.083 37.283 108.115 37.347 ;
			RECT	108.419 37.283 108.451 37.347 ;
			RECT	108.755 37.283 108.787 37.347 ;
			RECT	109.091 37.283 109.123 37.347 ;
			RECT	109.427 37.283 109.459 37.347 ;
			RECT	109.763 37.283 109.795 37.347 ;
			RECT	110.099 37.283 110.131 37.347 ;
			RECT	110.435 37.283 110.467 37.347 ;
			RECT	110.771 37.283 110.803 37.347 ;
			RECT	111.107 37.283 111.139 37.347 ;
			RECT	111.443 37.283 111.475 37.347 ;
			RECT	111.779 37.283 111.811 37.347 ;
			RECT	112.115 37.283 112.147 37.347 ;
			RECT	112.451 37.283 112.483 37.347 ;
			RECT	112.787 37.283 112.819 37.347 ;
			RECT	113.123 37.283 113.155 37.347 ;
			RECT	113.459 37.283 113.491 37.347 ;
			RECT	113.795 37.283 113.827 37.347 ;
			RECT	114.131 37.283 114.163 37.347 ;
			RECT	114.467 37.283 114.499 37.347 ;
			RECT	114.803 37.283 114.835 37.347 ;
			RECT	115.139 37.283 115.171 37.347 ;
			RECT	115.475 37.283 115.507 37.347 ;
			RECT	115.811 37.283 115.843 37.347 ;
			RECT	116.147 37.283 116.179 37.347 ;
			RECT	116.483 37.283 116.515 37.347 ;
			RECT	116.819 37.283 116.851 37.347 ;
			RECT	117.155 37.283 117.187 37.347 ;
			RECT	117.491 37.283 117.523 37.347 ;
			RECT	117.827 37.283 117.859 37.347 ;
			RECT	118.163 37.283 118.195 37.347 ;
			RECT	118.499 37.283 118.531 37.347 ;
			RECT	118.835 37.283 118.867 37.347 ;
			RECT	119.171 37.283 119.203 37.347 ;
			RECT	119.507 37.283 119.539 37.347 ;
			RECT	119.843 37.283 119.875 37.347 ;
			RECT	120.179 37.283 120.211 37.347 ;
			RECT	120.515 37.283 120.547 37.347 ;
			RECT	120.851 37.283 120.883 37.347 ;
			RECT	121.187 37.283 121.219 37.347 ;
			RECT	121.523 37.283 121.555 37.347 ;
			RECT	121.859 37.283 121.891 37.347 ;
			RECT	122.195 37.283 122.227 37.347 ;
			RECT	122.531 37.283 122.563 37.347 ;
			RECT	122.867 37.283 122.899 37.347 ;
			RECT	123.203 37.283 123.235 37.347 ;
			RECT	123.539 37.283 123.571 37.347 ;
			RECT	123.875 37.283 123.907 37.347 ;
			RECT	124.211 37.283 124.243 37.347 ;
			RECT	124.547 37.283 124.579 37.347 ;
			RECT	124.883 37.283 124.915 37.347 ;
			RECT	125.219 37.283 125.251 37.347 ;
			RECT	125.555 37.283 125.587 37.347 ;
			RECT	125.886 37.283 125.918 37.347 ;
			RECT	126.222 37.283 126.254 37.347 ;
			RECT	126.558 37.283 126.59 37.347 ;
			RECT	126.894 37.283 126.926 37.347 ;
			RECT	127.23 37.283 127.262 37.347 ;
			RECT	127.566 37.283 127.598 37.347 ;
			RECT	127.902 37.283 127.934 37.347 ;
			RECT	128.238 37.283 128.27 37.347 ;
			RECT	128.574 37.283 128.606 37.347 ;
			RECT	128.91 37.283 128.942 37.347 ;
			RECT	129.246 37.283 129.278 37.347 ;
			RECT	129.582 37.283 129.614 37.347 ;
			RECT	129.918 37.283 129.95 37.347 ;
			RECT	130.254 37.283 130.286 37.347 ;
			RECT	130.59 37.283 130.622 37.347 ;
			RECT	130.926 37.283 130.958 37.347 ;
			RECT	132.606 37.283 132.638 37.347 ;
			RECT	132.942 37.283 132.974 37.347 ;
			RECT	133.278 37.283 133.31 37.347 ;
			RECT	133.614 37.283 133.646 37.347 ;
			RECT	134.286 37.283 134.318 37.347 ;
			RECT	134.958 37.283 134.99 37.347 ;
			RECT	135.63 37.283 135.662 37.347 ;
			RECT	135.966 37.283 135.998 37.347 ;
			RECT	136.302 37.283 136.334 37.347 ;
			RECT	136.638 37.283 136.67 37.347 ;
			RECT	136.974 37.283 137.006 37.347 ;
			RECT	137.646 37.283 137.678 37.347 ;
			RECT	137.982 37.283 138.014 37.347 ;
			RECT	138.318 37.283 138.35 37.347 ;
			RECT	138.99 37.283 139.022 37.347 ;
			RECT	139.662 37.283 139.694 37.347 ;
			RECT	139.998 37.283 140.03 37.347 ;
			RECT	140.334 37.283 140.366 37.347 ;
			RECT	140.67 37.283 140.702 37.347 ;
			RECT	141.006 37.283 141.038 37.347 ;
			RECT	141.342 37.283 141.374 37.347 ;
			RECT	141.678 37.283 141.71 37.347 ;
			RECT	142.678 37.283 142.71 37.347 ;
			RECT	143.022 37.283 143.054 37.347 ;
			RECT	144.03 37.283 144.062 37.347 ;
			RECT	144.366 37.283 144.398 37.347 ;
			RECT	145.038 37.283 145.07 37.347 ;
			RECT	145.374 37.283 145.406 37.347 ;
			RECT	146.046 37.283 146.078 37.347 ;
			RECT	146.382 37.283 146.414 37.347 ;
			RECT	146.718 37.283 146.75 37.347 ;
			RECT	147.054 37.283 147.086 37.347 ;
			RECT	147.309 37.283 147.373 37.347 ;
			RECT	147.611 37.283 147.643 37.347 ;
			RECT	149.918 37.299 149.95 37.331 ;
			RECT	150.966 37.283 151.03 37.347 ;
			RECT	151.908 37.283 151.94 37.347 ;
			RECT	152.81 37.283 152.842 37.347 ;
			RECT	153.967 37.283 154.031 37.347 ;
			RECT	155.909 37.283 155.941 37.347 ;
			RECT	156.557 37.283 156.589 37.347 ;
			RECT	156.827 37.283 156.891 37.347 ;
			RECT	157.114 37.283 157.146 37.347 ;
			RECT	157.45 37.283 157.482 37.347 ;
			RECT	157.786 37.283 157.818 37.347 ;
			RECT	158.122 37.283 158.154 37.347 ;
			RECT	158.794 37.283 158.826 37.347 ;
			RECT	159.13 37.283 159.162 37.347 ;
			RECT	159.802 37.283 159.834 37.347 ;
			RECT	160.138 37.283 160.17 37.347 ;
			RECT	161.146 37.283 161.178 37.347 ;
			RECT	161.49 37.283 161.522 37.347 ;
			RECT	162.49 37.283 162.522 37.347 ;
			RECT	162.826 37.283 162.858 37.347 ;
			RECT	163.162 37.283 163.194 37.347 ;
			RECT	163.498 37.283 163.53 37.347 ;
			RECT	163.834 37.283 163.866 37.347 ;
			RECT	164.17 37.283 164.202 37.347 ;
			RECT	164.506 37.283 164.538 37.347 ;
			RECT	165.178 37.283 165.21 37.347 ;
			RECT	165.85 37.283 165.882 37.347 ;
			RECT	166.186 37.283 166.218 37.347 ;
			RECT	166.522 37.283 166.554 37.347 ;
			RECT	167.194 37.283 167.226 37.347 ;
			RECT	167.53 37.283 167.562 37.347 ;
			RECT	167.866 37.283 167.898 37.347 ;
			RECT	168.202 37.283 168.234 37.347 ;
			RECT	168.538 37.283 168.57 37.347 ;
			RECT	169.21 37.283 169.242 37.347 ;
			RECT	169.882 37.283 169.914 37.347 ;
			RECT	170.554 37.283 170.586 37.347 ;
			RECT	170.89 37.283 170.922 37.347 ;
			RECT	171.226 37.283 171.258 37.347 ;
			RECT	171.562 37.283 171.594 37.347 ;
			RECT	173.242 37.283 173.274 37.347 ;
			RECT	173.578 37.283 173.61 37.347 ;
			RECT	173.914 37.283 173.946 37.347 ;
			RECT	174.25 37.283 174.282 37.347 ;
			RECT	174.586 37.283 174.618 37.347 ;
			RECT	174.922 37.283 174.954 37.347 ;
			RECT	175.258 37.283 175.29 37.347 ;
			RECT	175.594 37.283 175.626 37.347 ;
			RECT	175.93 37.283 175.962 37.347 ;
			RECT	176.266 37.283 176.298 37.347 ;
			RECT	176.602 37.283 176.634 37.347 ;
			RECT	176.938 37.283 176.97 37.347 ;
			RECT	177.274 37.283 177.306 37.347 ;
			RECT	177.61 37.283 177.642 37.347 ;
			RECT	177.946 37.283 177.978 37.347 ;
			RECT	178.282 37.283 178.314 37.347 ;
			RECT	178.613 37.283 178.645 37.347 ;
			RECT	178.949 37.283 178.981 37.347 ;
			RECT	179.285 37.283 179.317 37.347 ;
			RECT	179.621 37.283 179.653 37.347 ;
			RECT	179.957 37.283 179.989 37.347 ;
			RECT	180.293 37.283 180.325 37.347 ;
			RECT	180.629 37.283 180.661 37.347 ;
			RECT	180.965 37.283 180.997 37.347 ;
			RECT	181.301 37.283 181.333 37.347 ;
			RECT	181.637 37.283 181.669 37.347 ;
			RECT	181.973 37.283 182.005 37.347 ;
			RECT	182.309 37.283 182.341 37.347 ;
			RECT	182.645 37.283 182.677 37.347 ;
			RECT	182.981 37.283 183.013 37.347 ;
			RECT	183.317 37.283 183.349 37.347 ;
			RECT	183.653 37.283 183.685 37.347 ;
			RECT	183.989 37.283 184.021 37.347 ;
			RECT	184.325 37.283 184.357 37.347 ;
			RECT	184.661 37.283 184.693 37.347 ;
			RECT	184.997 37.283 185.029 37.347 ;
			RECT	185.333 37.283 185.365 37.347 ;
			RECT	185.669 37.283 185.701 37.347 ;
			RECT	186.005 37.283 186.037 37.347 ;
			RECT	186.341 37.283 186.373 37.347 ;
			RECT	186.677 37.283 186.709 37.347 ;
			RECT	187.013 37.283 187.045 37.347 ;
			RECT	187.349 37.283 187.381 37.347 ;
			RECT	187.685 37.283 187.717 37.347 ;
			RECT	188.021 37.283 188.053 37.347 ;
			RECT	188.357 37.283 188.389 37.347 ;
			RECT	188.693 37.283 188.725 37.347 ;
			RECT	189.029 37.283 189.061 37.347 ;
			RECT	189.365 37.283 189.397 37.347 ;
			RECT	189.701 37.283 189.733 37.347 ;
			RECT	190.037 37.283 190.069 37.347 ;
			RECT	190.373 37.283 190.405 37.347 ;
			RECT	190.709 37.283 190.741 37.347 ;
			RECT	191.045 37.283 191.077 37.347 ;
			RECT	191.381 37.283 191.413 37.347 ;
			RECT	191.717 37.283 191.749 37.347 ;
			RECT	192.053 37.283 192.085 37.347 ;
			RECT	192.389 37.283 192.421 37.347 ;
			RECT	192.725 37.283 192.757 37.347 ;
			RECT	193.061 37.283 193.093 37.347 ;
			RECT	193.397 37.283 193.429 37.347 ;
			RECT	193.733 37.283 193.765 37.347 ;
			RECT	194.069 37.283 194.101 37.347 ;
			RECT	194.405 37.283 194.437 37.347 ;
			RECT	194.741 37.283 194.773 37.347 ;
			RECT	195.077 37.283 195.109 37.347 ;
			RECT	195.413 37.283 195.445 37.347 ;
			RECT	195.749 37.283 195.781 37.347 ;
			RECT	196.085 37.283 196.117 37.347 ;
			RECT	196.421 37.283 196.453 37.347 ;
			RECT	196.757 37.283 196.789 37.347 ;
			RECT	197.093 37.283 197.125 37.347 ;
			RECT	197.429 37.283 197.461 37.347 ;
			RECT	197.765 37.283 197.797 37.347 ;
			RECT	198.101 37.283 198.133 37.347 ;
			RECT	198.437 37.283 198.469 37.347 ;
			RECT	198.773 37.283 198.805 37.347 ;
			RECT	199.109 37.283 199.141 37.347 ;
			RECT	199.445 37.283 199.477 37.347 ;
			RECT	199.781 37.283 199.813 37.347 ;
			RECT	200.412 37.283 200.444 37.347 ;
			RECT	200.9 37.283 200.932 37.347 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 37.995 201.665 38.085 ;
			LAYER	J3 ;
			RECT	1.661 38.008 1.693 38.072 ;
			RECT	2.323 38.024 2.387 38.056 ;
			RECT	3.438 38.024 3.47 38.056 ;
			RECT	4.539 38.008 4.571 38.072 ;
			RECT	4.805 38.008 4.837 38.072 ;
			RECT	5.252 38.008 5.284 38.072 ;
			RECT	5.758 38.007 5.79 38.071 ;
			RECT	6.389 38.008 6.421 38.072 ;
			RECT	6.725 38.008 6.757 38.072 ;
			RECT	7.061 38.008 7.093 38.072 ;
			RECT	7.397 38.008 7.429 38.072 ;
			RECT	7.733 38.008 7.765 38.072 ;
			RECT	8.069 38.008 8.101 38.072 ;
			RECT	8.405 38.008 8.437 38.072 ;
			RECT	8.741 38.008 8.773 38.072 ;
			RECT	9.077 38.008 9.109 38.072 ;
			RECT	9.413 38.008 9.445 38.072 ;
			RECT	9.749 38.008 9.781 38.072 ;
			RECT	10.085 38.008 10.117 38.072 ;
			RECT	10.421 38.008 10.453 38.072 ;
			RECT	10.757 38.008 10.789 38.072 ;
			RECT	11.093 38.008 11.125 38.072 ;
			RECT	11.429 38.008 11.461 38.072 ;
			RECT	11.765 38.008 11.797 38.072 ;
			RECT	12.101 38.008 12.133 38.072 ;
			RECT	12.437 38.008 12.469 38.072 ;
			RECT	12.773 38.008 12.805 38.072 ;
			RECT	13.109 38.008 13.141 38.072 ;
			RECT	13.445 38.008 13.477 38.072 ;
			RECT	13.781 38.008 13.813 38.072 ;
			RECT	14.117 38.008 14.149 38.072 ;
			RECT	14.453 38.008 14.485 38.072 ;
			RECT	14.789 38.008 14.821 38.072 ;
			RECT	15.125 38.008 15.157 38.072 ;
			RECT	15.461 38.008 15.493 38.072 ;
			RECT	15.797 38.008 15.829 38.072 ;
			RECT	16.133 38.008 16.165 38.072 ;
			RECT	16.469 38.008 16.501 38.072 ;
			RECT	16.805 38.008 16.837 38.072 ;
			RECT	17.141 38.008 17.173 38.072 ;
			RECT	17.477 38.008 17.509 38.072 ;
			RECT	17.813 38.008 17.845 38.072 ;
			RECT	18.149 38.008 18.181 38.072 ;
			RECT	18.485 38.008 18.517 38.072 ;
			RECT	18.821 38.008 18.853 38.072 ;
			RECT	19.157 38.008 19.189 38.072 ;
			RECT	19.493 38.008 19.525 38.072 ;
			RECT	19.829 38.008 19.861 38.072 ;
			RECT	20.165 38.008 20.197 38.072 ;
			RECT	20.501 38.008 20.533 38.072 ;
			RECT	20.837 38.008 20.869 38.072 ;
			RECT	21.173 38.008 21.205 38.072 ;
			RECT	21.509 38.008 21.541 38.072 ;
			RECT	21.845 38.008 21.877 38.072 ;
			RECT	22.181 38.008 22.213 38.072 ;
			RECT	22.517 38.008 22.549 38.072 ;
			RECT	22.853 38.008 22.885 38.072 ;
			RECT	23.189 38.008 23.221 38.072 ;
			RECT	23.525 38.008 23.557 38.072 ;
			RECT	23.861 38.008 23.893 38.072 ;
			RECT	24.197 38.008 24.229 38.072 ;
			RECT	24.533 38.008 24.565 38.072 ;
			RECT	24.869 38.008 24.901 38.072 ;
			RECT	25.205 38.008 25.237 38.072 ;
			RECT	25.541 38.008 25.573 38.072 ;
			RECT	25.877 38.008 25.909 38.072 ;
			RECT	26.213 38.008 26.245 38.072 ;
			RECT	26.549 38.008 26.581 38.072 ;
			RECT	26.885 38.008 26.917 38.072 ;
			RECT	27.221 38.008 27.253 38.072 ;
			RECT	27.557 38.008 27.589 38.072 ;
			RECT	27.888 38.024 27.92 38.056 ;
			RECT	28.224 38.024 28.256 38.056 ;
			RECT	28.56 38.024 28.592 38.056 ;
			RECT	28.896 38.008 28.928 38.072 ;
			RECT	29.232 38.024 29.264 38.056 ;
			RECT	29.568 38.024 29.6 38.056 ;
			RECT	29.904 38.024 29.936 38.056 ;
			RECT	30.24 38.024 30.272 38.056 ;
			RECT	30.576 38.008 30.608 38.072 ;
			RECT	30.912 38.024 30.944 38.056 ;
			RECT	31.248 38.024 31.28 38.056 ;
			RECT	31.584 38.024 31.616 38.056 ;
			RECT	31.92 38.008 31.952 38.072 ;
			RECT	32.256 38.024 32.288 38.056 ;
			RECT	32.592 38.024 32.624 38.056 ;
			RECT	32.928 38.024 32.96 38.056 ;
			RECT	34.608 38.024 34.64 38.056 ;
			RECT	34.944 38.024 34.976 38.056 ;
			RECT	35.28 38.008 35.312 38.072 ;
			RECT	35.616 38.024 35.648 38.056 ;
			RECT	37.632 38.024 37.664 38.056 ;
			RECT	37.968 38.024 38 38.056 ;
			RECT	38.304 38.024 38.336 38.056 ;
			RECT	38.64 38.008 38.672 38.072 ;
			RECT	38.976 38.024 39.008 38.056 ;
			RECT	39.648 38.024 39.68 38.056 ;
			RECT	39.984 38.024 40.016 38.056 ;
			RECT	41.664 38.024 41.696 38.056 ;
			RECT	42 38.024 42.032 38.056 ;
			RECT	42.336 38.024 42.368 38.056 ;
			RECT	42.672 38.008 42.704 38.072 ;
			RECT	43.008 38.024 43.04 38.056 ;
			RECT	43.344 38.024 43.376 38.056 ;
			RECT	43.68 38.024 43.712 38.056 ;
			RECT	44.68 38.024 44.712 38.056 ;
			RECT	45.024 38.024 45.056 38.056 ;
			RECT	46.032 38.024 46.064 38.056 ;
			RECT	46.368 38.008 46.4 38.072 ;
			RECT	47.04 38.024 47.072 38.056 ;
			RECT	47.376 38.024 47.408 38.056 ;
			RECT	48.048 38.024 48.08 38.056 ;
			RECT	48.384 38.008 48.416 38.072 ;
			RECT	48.72 38.024 48.752 38.056 ;
			RECT	49.056 38.024 49.088 38.056 ;
			RECT	49.311 38.024 49.375 38.056 ;
			RECT	51.92 38.008 51.952 38.072 ;
			RECT	52.968 38.024 53.032 38.056 ;
			RECT	53.894 38.008 53.926 38.072 ;
			RECT	54.812 38.004 54.844 38.068 ;
			RECT	55.969 38.024 56.033 38.056 ;
			RECT	57.18 38.008 57.212 38.072 ;
			RECT	57.363 38.008 57.395 38.072 ;
			RECT	57.911 38.008 57.943 38.072 ;
			RECT	58.829 38.024 58.893 38.056 ;
			RECT	59.116 38.024 59.148 38.056 ;
			RECT	59.452 38.024 59.484 38.056 ;
			RECT	59.788 38.008 59.82 38.072 ;
			RECT	60.124 38.024 60.156 38.056 ;
			RECT	60.796 38.024 60.828 38.056 ;
			RECT	61.132 38.024 61.164 38.056 ;
			RECT	61.804 38.008 61.836 38.072 ;
			RECT	62.14 38.024 62.172 38.056 ;
			RECT	63.148 38.024 63.18 38.056 ;
			RECT	63.492 38.024 63.524 38.056 ;
			RECT	64.492 38.024 64.524 38.056 ;
			RECT	64.828 38.024 64.86 38.056 ;
			RECT	65.164 38.024 65.196 38.056 ;
			RECT	65.5 38.008 65.532 38.072 ;
			RECT	65.836 38.024 65.868 38.056 ;
			RECT	66.172 38.024 66.204 38.056 ;
			RECT	66.508 38.024 66.54 38.056 ;
			RECT	68.188 38.024 68.22 38.056 ;
			RECT	68.524 38.024 68.556 38.056 ;
			RECT	69.196 38.024 69.228 38.056 ;
			RECT	69.532 38.008 69.564 38.072 ;
			RECT	69.868 38.024 69.9 38.056 ;
			RECT	70.204 38.024 70.236 38.056 ;
			RECT	70.54 38.024 70.572 38.056 ;
			RECT	72.556 38.024 72.588 38.056 ;
			RECT	72.892 38.008 72.924 38.072 ;
			RECT	73.228 38.024 73.26 38.056 ;
			RECT	73.564 38.024 73.596 38.056 ;
			RECT	75.244 38.024 75.276 38.056 ;
			RECT	75.58 38.024 75.612 38.056 ;
			RECT	75.916 38.024 75.948 38.056 ;
			RECT	76.252 38.008 76.284 38.072 ;
			RECT	76.588 38.024 76.62 38.056 ;
			RECT	76.924 38.024 76.956 38.056 ;
			RECT	77.26 38.024 77.292 38.056 ;
			RECT	77.596 38.008 77.628 38.072 ;
			RECT	77.932 38.024 77.964 38.056 ;
			RECT	78.268 38.024 78.3 38.056 ;
			RECT	78.604 38.024 78.636 38.056 ;
			RECT	78.94 38.024 78.972 38.056 ;
			RECT	79.276 38.008 79.308 38.072 ;
			RECT	79.612 38.024 79.644 38.056 ;
			RECT	79.948 38.024 79.98 38.056 ;
			RECT	80.284 38.024 80.316 38.056 ;
			RECT	80.615 38.008 80.647 38.072 ;
			RECT	80.951 38.008 80.983 38.072 ;
			RECT	81.287 38.008 81.319 38.072 ;
			RECT	81.623 38.008 81.655 38.072 ;
			RECT	81.959 38.008 81.991 38.072 ;
			RECT	82.295 38.008 82.327 38.072 ;
			RECT	82.631 38.008 82.663 38.072 ;
			RECT	82.967 38.008 82.999 38.072 ;
			RECT	83.303 38.008 83.335 38.072 ;
			RECT	83.639 38.008 83.671 38.072 ;
			RECT	83.975 38.008 84.007 38.072 ;
			RECT	84.311 38.008 84.343 38.072 ;
			RECT	84.647 38.008 84.679 38.072 ;
			RECT	84.983 38.008 85.015 38.072 ;
			RECT	85.319 38.008 85.351 38.072 ;
			RECT	85.655 38.008 85.687 38.072 ;
			RECT	85.991 38.008 86.023 38.072 ;
			RECT	86.327 38.008 86.359 38.072 ;
			RECT	86.663 38.008 86.695 38.072 ;
			RECT	86.999 38.008 87.031 38.072 ;
			RECT	87.335 38.008 87.367 38.072 ;
			RECT	87.671 38.008 87.703 38.072 ;
			RECT	88.007 38.008 88.039 38.072 ;
			RECT	88.343 38.008 88.375 38.072 ;
			RECT	88.679 38.008 88.711 38.072 ;
			RECT	89.015 38.008 89.047 38.072 ;
			RECT	89.351 38.008 89.383 38.072 ;
			RECT	89.687 38.008 89.719 38.072 ;
			RECT	90.023 38.008 90.055 38.072 ;
			RECT	90.359 38.008 90.391 38.072 ;
			RECT	90.695 38.008 90.727 38.072 ;
			RECT	91.031 38.008 91.063 38.072 ;
			RECT	91.367 38.008 91.399 38.072 ;
			RECT	91.703 38.008 91.735 38.072 ;
			RECT	92.039 38.008 92.071 38.072 ;
			RECT	92.375 38.008 92.407 38.072 ;
			RECT	92.711 38.008 92.743 38.072 ;
			RECT	93.047 38.008 93.079 38.072 ;
			RECT	93.383 38.008 93.415 38.072 ;
			RECT	93.719 38.008 93.751 38.072 ;
			RECT	94.055 38.008 94.087 38.072 ;
			RECT	94.391 38.008 94.423 38.072 ;
			RECT	94.727 38.008 94.759 38.072 ;
			RECT	95.063 38.008 95.095 38.072 ;
			RECT	95.399 38.008 95.431 38.072 ;
			RECT	95.735 38.008 95.767 38.072 ;
			RECT	96.071 38.008 96.103 38.072 ;
			RECT	96.407 38.008 96.439 38.072 ;
			RECT	96.743 38.008 96.775 38.072 ;
			RECT	97.079 38.008 97.111 38.072 ;
			RECT	97.415 38.008 97.447 38.072 ;
			RECT	97.751 38.008 97.783 38.072 ;
			RECT	98.087 38.008 98.119 38.072 ;
			RECT	98.423 38.008 98.455 38.072 ;
			RECT	98.759 38.008 98.791 38.072 ;
			RECT	99.095 38.008 99.127 38.072 ;
			RECT	99.431 38.008 99.463 38.072 ;
			RECT	99.767 38.008 99.799 38.072 ;
			RECT	100.103 38.008 100.135 38.072 ;
			RECT	100.439 38.008 100.471 38.072 ;
			RECT	100.775 38.008 100.807 38.072 ;
			RECT	101.111 38.008 101.143 38.072 ;
			RECT	101.447 38.008 101.479 38.072 ;
			RECT	101.783 38.008 101.815 38.072 ;
			RECT	102.414 38.007 102.446 38.071 ;
			RECT	103.756 38.007 103.788 38.071 ;
			RECT	104.387 38.008 104.419 38.072 ;
			RECT	104.723 38.008 104.755 38.072 ;
			RECT	105.059 38.008 105.091 38.072 ;
			RECT	105.395 38.008 105.427 38.072 ;
			RECT	105.731 38.008 105.763 38.072 ;
			RECT	106.067 38.008 106.099 38.072 ;
			RECT	106.403 38.008 106.435 38.072 ;
			RECT	106.739 38.008 106.771 38.072 ;
			RECT	107.075 38.008 107.107 38.072 ;
			RECT	107.411 38.008 107.443 38.072 ;
			RECT	107.747 38.008 107.779 38.072 ;
			RECT	108.083 38.008 108.115 38.072 ;
			RECT	108.419 38.008 108.451 38.072 ;
			RECT	108.755 38.008 108.787 38.072 ;
			RECT	109.091 38.008 109.123 38.072 ;
			RECT	109.427 38.008 109.459 38.072 ;
			RECT	109.763 38.008 109.795 38.072 ;
			RECT	110.099 38.008 110.131 38.072 ;
			RECT	110.435 38.008 110.467 38.072 ;
			RECT	110.771 38.008 110.803 38.072 ;
			RECT	111.107 38.008 111.139 38.072 ;
			RECT	111.443 38.008 111.475 38.072 ;
			RECT	111.779 38.008 111.811 38.072 ;
			RECT	112.115 38.008 112.147 38.072 ;
			RECT	112.451 38.008 112.483 38.072 ;
			RECT	112.787 38.008 112.819 38.072 ;
			RECT	113.123 38.008 113.155 38.072 ;
			RECT	113.459 38.008 113.491 38.072 ;
			RECT	113.795 38.008 113.827 38.072 ;
			RECT	114.131 38.008 114.163 38.072 ;
			RECT	114.467 38.008 114.499 38.072 ;
			RECT	114.803 38.008 114.835 38.072 ;
			RECT	115.139 38.008 115.171 38.072 ;
			RECT	115.475 38.008 115.507 38.072 ;
			RECT	115.811 38.008 115.843 38.072 ;
			RECT	116.147 38.008 116.179 38.072 ;
			RECT	116.483 38.008 116.515 38.072 ;
			RECT	116.819 38.008 116.851 38.072 ;
			RECT	117.155 38.008 117.187 38.072 ;
			RECT	117.491 38.008 117.523 38.072 ;
			RECT	117.827 38.008 117.859 38.072 ;
			RECT	118.163 38.008 118.195 38.072 ;
			RECT	118.499 38.008 118.531 38.072 ;
			RECT	118.835 38.008 118.867 38.072 ;
			RECT	119.171 38.008 119.203 38.072 ;
			RECT	119.507 38.008 119.539 38.072 ;
			RECT	119.843 38.008 119.875 38.072 ;
			RECT	120.179 38.008 120.211 38.072 ;
			RECT	120.515 38.008 120.547 38.072 ;
			RECT	120.851 38.008 120.883 38.072 ;
			RECT	121.187 38.008 121.219 38.072 ;
			RECT	121.523 38.008 121.555 38.072 ;
			RECT	121.859 38.008 121.891 38.072 ;
			RECT	122.195 38.008 122.227 38.072 ;
			RECT	122.531 38.008 122.563 38.072 ;
			RECT	122.867 38.008 122.899 38.072 ;
			RECT	123.203 38.008 123.235 38.072 ;
			RECT	123.539 38.008 123.571 38.072 ;
			RECT	123.875 38.008 123.907 38.072 ;
			RECT	124.211 38.008 124.243 38.072 ;
			RECT	124.547 38.008 124.579 38.072 ;
			RECT	124.883 38.008 124.915 38.072 ;
			RECT	125.219 38.008 125.251 38.072 ;
			RECT	125.555 38.008 125.587 38.072 ;
			RECT	125.886 38.024 125.918 38.056 ;
			RECT	126.222 38.024 126.254 38.056 ;
			RECT	126.558 38.024 126.59 38.056 ;
			RECT	126.894 38.008 126.926 38.072 ;
			RECT	127.23 38.024 127.262 38.056 ;
			RECT	127.566 38.024 127.598 38.056 ;
			RECT	127.902 38.024 127.934 38.056 ;
			RECT	128.238 38.024 128.27 38.056 ;
			RECT	128.574 38.008 128.606 38.072 ;
			RECT	128.91 38.024 128.942 38.056 ;
			RECT	129.246 38.024 129.278 38.056 ;
			RECT	129.582 38.024 129.614 38.056 ;
			RECT	129.918 38.008 129.95 38.072 ;
			RECT	130.254 38.024 130.286 38.056 ;
			RECT	130.59 38.024 130.622 38.056 ;
			RECT	130.926 38.024 130.958 38.056 ;
			RECT	132.606 38.024 132.638 38.056 ;
			RECT	132.942 38.024 132.974 38.056 ;
			RECT	133.278 38.008 133.31 38.072 ;
			RECT	133.614 38.024 133.646 38.056 ;
			RECT	135.63 38.024 135.662 38.056 ;
			RECT	135.966 38.024 135.998 38.056 ;
			RECT	136.302 38.024 136.334 38.056 ;
			RECT	136.638 38.008 136.67 38.072 ;
			RECT	136.974 38.024 137.006 38.056 ;
			RECT	137.646 38.024 137.678 38.056 ;
			RECT	137.982 38.024 138.014 38.056 ;
			RECT	139.662 38.024 139.694 38.056 ;
			RECT	139.998 38.024 140.03 38.056 ;
			RECT	140.334 38.024 140.366 38.056 ;
			RECT	140.67 38.008 140.702 38.072 ;
			RECT	141.006 38.024 141.038 38.056 ;
			RECT	141.342 38.024 141.374 38.056 ;
			RECT	141.678 38.024 141.71 38.056 ;
			RECT	142.678 38.024 142.71 38.056 ;
			RECT	143.022 38.024 143.054 38.056 ;
			RECT	144.03 38.024 144.062 38.056 ;
			RECT	144.366 38.008 144.398 38.072 ;
			RECT	145.038 38.024 145.07 38.056 ;
			RECT	145.374 38.024 145.406 38.056 ;
			RECT	146.046 38.024 146.078 38.056 ;
			RECT	146.382 38.008 146.414 38.072 ;
			RECT	146.718 38.024 146.75 38.056 ;
			RECT	147.054 38.024 147.086 38.056 ;
			RECT	147.309 38.024 147.373 38.056 ;
			RECT	149.918 38.008 149.95 38.072 ;
			RECT	150.966 38.024 151.03 38.056 ;
			RECT	151.892 38.008 151.924 38.072 ;
			RECT	152.81 38.004 152.842 38.068 ;
			RECT	153.967 38.024 154.031 38.056 ;
			RECT	155.178 38.008 155.21 38.072 ;
			RECT	155.361 38.008 155.393 38.072 ;
			RECT	155.909 38.008 155.941 38.072 ;
			RECT	156.827 38.024 156.891 38.056 ;
			RECT	157.114 38.024 157.146 38.056 ;
			RECT	157.45 38.024 157.482 38.056 ;
			RECT	157.786 38.008 157.818 38.072 ;
			RECT	158.122 38.024 158.154 38.056 ;
			RECT	158.794 38.024 158.826 38.056 ;
			RECT	159.13 38.024 159.162 38.056 ;
			RECT	159.802 38.008 159.834 38.072 ;
			RECT	160.138 38.024 160.17 38.056 ;
			RECT	161.146 38.024 161.178 38.056 ;
			RECT	161.49 38.024 161.522 38.056 ;
			RECT	162.49 38.024 162.522 38.056 ;
			RECT	162.826 38.024 162.858 38.056 ;
			RECT	163.162 38.024 163.194 38.056 ;
			RECT	163.498 38.008 163.53 38.072 ;
			RECT	163.834 38.024 163.866 38.056 ;
			RECT	164.17 38.024 164.202 38.056 ;
			RECT	164.506 38.024 164.538 38.056 ;
			RECT	166.186 38.024 166.218 38.056 ;
			RECT	166.522 38.024 166.554 38.056 ;
			RECT	167.194 38.024 167.226 38.056 ;
			RECT	167.53 38.008 167.562 38.072 ;
			RECT	167.866 38.024 167.898 38.056 ;
			RECT	168.202 38.024 168.234 38.056 ;
			RECT	168.538 38.024 168.57 38.056 ;
			RECT	170.554 38.024 170.586 38.056 ;
			RECT	170.89 38.008 170.922 38.072 ;
			RECT	171.226 38.024 171.258 38.056 ;
			RECT	171.562 38.024 171.594 38.056 ;
			RECT	173.242 38.024 173.274 38.056 ;
			RECT	173.578 38.024 173.61 38.056 ;
			RECT	173.914 38.024 173.946 38.056 ;
			RECT	174.25 38.008 174.282 38.072 ;
			RECT	174.586 38.024 174.618 38.056 ;
			RECT	174.922 38.024 174.954 38.056 ;
			RECT	175.258 38.024 175.29 38.056 ;
			RECT	175.594 38.008 175.626 38.072 ;
			RECT	175.93 38.024 175.962 38.056 ;
			RECT	176.266 38.024 176.298 38.056 ;
			RECT	176.602 38.024 176.634 38.056 ;
			RECT	176.938 38.024 176.97 38.056 ;
			RECT	177.274 38.008 177.306 38.072 ;
			RECT	177.61 38.024 177.642 38.056 ;
			RECT	177.946 38.024 177.978 38.056 ;
			RECT	178.282 38.024 178.314 38.056 ;
			RECT	178.613 38.008 178.645 38.072 ;
			RECT	178.949 38.008 178.981 38.072 ;
			RECT	179.285 38.008 179.317 38.072 ;
			RECT	179.621 38.008 179.653 38.072 ;
			RECT	179.957 38.008 179.989 38.072 ;
			RECT	180.293 38.008 180.325 38.072 ;
			RECT	180.629 38.008 180.661 38.072 ;
			RECT	180.965 38.008 180.997 38.072 ;
			RECT	181.301 38.008 181.333 38.072 ;
			RECT	181.637 38.008 181.669 38.072 ;
			RECT	181.973 38.008 182.005 38.072 ;
			RECT	182.309 38.008 182.341 38.072 ;
			RECT	182.645 38.008 182.677 38.072 ;
			RECT	182.981 38.008 183.013 38.072 ;
			RECT	183.317 38.008 183.349 38.072 ;
			RECT	183.653 38.008 183.685 38.072 ;
			RECT	183.989 38.008 184.021 38.072 ;
			RECT	184.325 38.008 184.357 38.072 ;
			RECT	184.661 38.008 184.693 38.072 ;
			RECT	184.997 38.008 185.029 38.072 ;
			RECT	185.333 38.008 185.365 38.072 ;
			RECT	185.669 38.008 185.701 38.072 ;
			RECT	186.005 38.008 186.037 38.072 ;
			RECT	186.341 38.008 186.373 38.072 ;
			RECT	186.677 38.008 186.709 38.072 ;
			RECT	187.013 38.008 187.045 38.072 ;
			RECT	187.349 38.008 187.381 38.072 ;
			RECT	187.685 38.008 187.717 38.072 ;
			RECT	188.021 38.008 188.053 38.072 ;
			RECT	188.357 38.008 188.389 38.072 ;
			RECT	188.693 38.008 188.725 38.072 ;
			RECT	189.029 38.008 189.061 38.072 ;
			RECT	189.365 38.008 189.397 38.072 ;
			RECT	189.701 38.008 189.733 38.072 ;
			RECT	190.037 38.008 190.069 38.072 ;
			RECT	190.373 38.008 190.405 38.072 ;
			RECT	190.709 38.008 190.741 38.072 ;
			RECT	191.045 38.008 191.077 38.072 ;
			RECT	191.381 38.008 191.413 38.072 ;
			RECT	191.717 38.008 191.749 38.072 ;
			RECT	192.053 38.008 192.085 38.072 ;
			RECT	192.389 38.008 192.421 38.072 ;
			RECT	192.725 38.008 192.757 38.072 ;
			RECT	193.061 38.008 193.093 38.072 ;
			RECT	193.397 38.008 193.429 38.072 ;
			RECT	193.733 38.008 193.765 38.072 ;
			RECT	194.069 38.008 194.101 38.072 ;
			RECT	194.405 38.008 194.437 38.072 ;
			RECT	194.741 38.008 194.773 38.072 ;
			RECT	195.077 38.008 195.109 38.072 ;
			RECT	195.413 38.008 195.445 38.072 ;
			RECT	195.749 38.008 195.781 38.072 ;
			RECT	196.085 38.008 196.117 38.072 ;
			RECT	196.421 38.008 196.453 38.072 ;
			RECT	196.757 38.008 196.789 38.072 ;
			RECT	197.093 38.008 197.125 38.072 ;
			RECT	197.429 38.008 197.461 38.072 ;
			RECT	197.765 38.008 197.797 38.072 ;
			RECT	198.101 38.008 198.133 38.072 ;
			RECT	198.437 38.008 198.469 38.072 ;
			RECT	198.773 38.008 198.805 38.072 ;
			RECT	199.109 38.008 199.141 38.072 ;
			RECT	199.445 38.008 199.477 38.072 ;
			RECT	199.781 38.008 199.813 38.072 ;
			RECT	200.412 38.007 200.444 38.071 ;
			RECT	200.9 38.008 200.932 38.072 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 38.984 201.665 39.074 ;
			LAYER	J3 ;
			RECT	1.661 38.997 1.693 39.061 ;
			RECT	2.323 39.013 2.387 39.045 ;
			RECT	3.305 38.997 3.337 39.061 ;
			RECT	3.438 38.997 3.47 39.061 ;
			RECT	4.354 38.997 4.386 39.061 ;
			RECT	4.536 38.997 4.568 39.061 ;
			RECT	4.805 38.997 4.837 39.061 ;
			RECT	5.252 38.997 5.284 39.061 ;
			RECT	5.758 38.998 5.79 39.062 ;
			RECT	28.56 39.013 28.592 39.045 ;
			RECT	28.896 38.997 28.928 39.061 ;
			RECT	29.232 39.013 29.264 39.045 ;
			RECT	29.904 39.013 29.936 39.045 ;
			RECT	30.24 38.997 30.272 39.061 ;
			RECT	30.576 38.997 30.608 39.061 ;
			RECT	30.912 39.013 30.944 39.045 ;
			RECT	31.248 38.997 31.28 39.061 ;
			RECT	31.584 39.013 31.616 39.045 ;
			RECT	31.92 38.997 31.952 39.061 ;
			RECT	32.592 38.997 32.624 39.061 ;
			RECT	33.264 38.997 33.296 39.061 ;
			RECT	34.272 38.997 34.304 39.061 ;
			RECT	35.28 38.997 35.312 39.061 ;
			RECT	35.952 38.997 35.984 39.061 ;
			RECT	37.632 38.997 37.664 39.061 ;
			RECT	38.64 38.997 38.672 39.061 ;
			RECT	39.648 38.997 39.68 39.061 ;
			RECT	41.328 38.997 41.36 39.061 ;
			RECT	42.336 38.997 42.368 39.061 ;
			RECT	42.672 38.997 42.704 39.061 ;
			RECT	43.344 39.013 43.376 39.045 ;
			RECT	43.68 38.997 43.712 39.061 ;
			RECT	46.368 38.997 46.4 39.061 ;
			RECT	47.04 38.997 47.072 39.061 ;
			RECT	49.091 38.997 49.123 39.061 ;
			RECT	49.311 39.013 49.375 39.045 ;
			RECT	50.417 39.013 50.481 39.045 ;
			RECT	51.92 38.997 51.952 39.061 ;
			RECT	52.15 38.997 52.182 39.061 ;
			RECT	52.454 38.997 52.486 39.061 ;
			RECT	52.968 39.013 53.032 39.045 ;
			RECT	53.91 38.997 53.942 39.061 ;
			RECT	54.379 38.997 54.411 39.061 ;
			RECT	54.812 38.997 54.844 39.061 ;
			RECT	55.224 38.997 55.256 39.061 ;
			RECT	55.578 38.997 55.61 39.061 ;
			RECT	55.985 38.997 56.017 39.061 ;
			RECT	56.144 38.998 56.176 39.062 ;
			RECT	57.363 38.997 57.395 39.061 ;
			RECT	58.829 39.013 58.893 39.045 ;
			RECT	59.081 38.997 59.113 39.061 ;
			RECT	61.132 38.997 61.164 39.061 ;
			RECT	61.804 38.997 61.836 39.061 ;
			RECT	64.492 38.997 64.524 39.061 ;
			RECT	64.828 39.013 64.86 39.045 ;
			RECT	65.5 38.997 65.532 39.061 ;
			RECT	65.836 38.997 65.868 39.061 ;
			RECT	66.844 38.997 66.876 39.061 ;
			RECT	68.524 38.997 68.556 39.061 ;
			RECT	69.532 38.997 69.564 39.061 ;
			RECT	70.54 38.997 70.572 39.061 ;
			RECT	72.22 38.997 72.252 39.061 ;
			RECT	72.892 38.997 72.924 39.061 ;
			RECT	73.9 38.997 73.932 39.061 ;
			RECT	74.908 38.997 74.94 39.061 ;
			RECT	75.58 38.997 75.612 39.061 ;
			RECT	76.252 38.997 76.284 39.061 ;
			RECT	76.588 39.013 76.62 39.045 ;
			RECT	76.924 38.997 76.956 39.061 ;
			RECT	77.26 39.013 77.292 39.045 ;
			RECT	77.596 38.997 77.628 39.061 ;
			RECT	77.932 38.997 77.964 39.061 ;
			RECT	78.268 39.013 78.3 39.045 ;
			RECT	78.94 39.013 78.972 39.045 ;
			RECT	79.276 38.997 79.308 39.061 ;
			RECT	79.612 39.013 79.644 39.045 ;
			RECT	102.414 38.998 102.446 39.062 ;
			RECT	103.756 38.998 103.788 39.062 ;
			RECT	126.558 39.013 126.59 39.045 ;
			RECT	126.894 38.997 126.926 39.061 ;
			RECT	127.23 39.013 127.262 39.045 ;
			RECT	127.902 39.013 127.934 39.045 ;
			RECT	128.238 38.997 128.27 39.061 ;
			RECT	128.574 38.997 128.606 39.061 ;
			RECT	128.91 39.013 128.942 39.045 ;
			RECT	129.246 38.997 129.278 39.061 ;
			RECT	129.582 39.013 129.614 39.045 ;
			RECT	129.918 38.997 129.95 39.061 ;
			RECT	130.59 38.997 130.622 39.061 ;
			RECT	131.262 38.997 131.294 39.061 ;
			RECT	132.27 38.997 132.302 39.061 ;
			RECT	133.278 38.997 133.31 39.061 ;
			RECT	133.95 38.997 133.982 39.061 ;
			RECT	135.63 38.997 135.662 39.061 ;
			RECT	136.638 38.997 136.67 39.061 ;
			RECT	137.646 38.997 137.678 39.061 ;
			RECT	139.326 38.997 139.358 39.061 ;
			RECT	140.334 38.997 140.366 39.061 ;
			RECT	140.67 38.997 140.702 39.061 ;
			RECT	141.342 39.013 141.374 39.045 ;
			RECT	141.678 38.997 141.71 39.061 ;
			RECT	144.366 38.997 144.398 39.061 ;
			RECT	145.038 38.997 145.07 39.061 ;
			RECT	147.089 38.997 147.121 39.061 ;
			RECT	147.309 39.013 147.373 39.045 ;
			RECT	148.415 39.013 148.479 39.045 ;
			RECT	149.918 38.997 149.95 39.061 ;
			RECT	150.148 38.997 150.18 39.061 ;
			RECT	150.452 38.997 150.484 39.061 ;
			RECT	150.966 39.013 151.03 39.045 ;
			RECT	151.908 38.997 151.94 39.061 ;
			RECT	152.377 38.997 152.409 39.061 ;
			RECT	152.81 38.997 152.842 39.061 ;
			RECT	153.222 38.997 153.254 39.061 ;
			RECT	153.576 38.997 153.608 39.061 ;
			RECT	153.983 38.997 154.015 39.061 ;
			RECT	154.142 38.998 154.174 39.062 ;
			RECT	155.361 38.997 155.393 39.061 ;
			RECT	156.827 39.013 156.891 39.045 ;
			RECT	157.079 38.997 157.111 39.061 ;
			RECT	159.13 38.997 159.162 39.061 ;
			RECT	159.802 38.997 159.834 39.061 ;
			RECT	162.49 38.997 162.522 39.061 ;
			RECT	162.826 39.013 162.858 39.045 ;
			RECT	163.498 38.997 163.53 39.061 ;
			RECT	163.834 38.997 163.866 39.061 ;
			RECT	164.842 38.997 164.874 39.061 ;
			RECT	166.522 38.997 166.554 39.061 ;
			RECT	167.53 38.997 167.562 39.061 ;
			RECT	168.538 38.997 168.57 39.061 ;
			RECT	170.218 38.997 170.25 39.061 ;
			RECT	170.89 38.997 170.922 39.061 ;
			RECT	171.898 38.997 171.93 39.061 ;
			RECT	172.906 38.997 172.938 39.061 ;
			RECT	173.578 38.997 173.61 39.061 ;
			RECT	174.25 38.997 174.282 39.061 ;
			RECT	174.586 39.013 174.618 39.045 ;
			RECT	174.922 38.997 174.954 39.061 ;
			RECT	175.258 39.013 175.29 39.045 ;
			RECT	175.594 38.997 175.626 39.061 ;
			RECT	175.93 38.997 175.962 39.061 ;
			RECT	176.266 39.013 176.298 39.045 ;
			RECT	176.938 39.013 176.97 39.045 ;
			RECT	177.274 38.997 177.306 39.061 ;
			RECT	177.61 39.013 177.642 39.045 ;
			RECT	200.412 38.998 200.444 39.062 ;
			RECT	200.9 38.997 200.932 39.061 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 40.149 201.665 40.269 ;
			LAYER	J3 ;
			RECT	1.645 40.177 1.709 40.241 ;
			RECT	2.197 40.177 2.229 40.241 ;
			RECT	2.323 40.177 2.387 40.241 ;
			RECT	3.438 40.177 3.47 40.241 ;
			RECT	4.354 40.177 4.386 40.241 ;
			RECT	4.536 40.177 4.568 40.241 ;
			RECT	5.252 40.177 5.284 40.241 ;
			RECT	5.758 40.177 5.79 40.241 ;
			RECT	27.888 40.177 27.92 40.241 ;
			RECT	28.56 40.177 28.592 40.241 ;
			RECT	29.232 40.177 29.264 40.241 ;
			RECT	29.904 40.177 29.936 40.241 ;
			RECT	30.576 40.177 30.608 40.241 ;
			RECT	31.92 40.177 31.952 40.241 ;
			RECT	33.264 40.177 33.296 40.241 ;
			RECT	34.272 40.177 34.304 40.241 ;
			RECT	34.608 40.177 34.64 40.241 ;
			RECT	37.296 40.177 37.328 40.241 ;
			RECT	38.64 40.177 38.672 40.241 ;
			RECT	39.648 40.177 39.68 40.241 ;
			RECT	39.984 40.177 40.016 40.241 ;
			RECT	40.32 40.177 40.352 40.241 ;
			RECT	40.656 40.177 40.688 40.241 ;
			RECT	43.344 40.177 43.376 40.241 ;
			RECT	44.016 40.177 44.048 40.241 ;
			RECT	44.688 40.177 44.72 40.241 ;
			RECT	46.032 40.177 46.064 40.241 ;
			RECT	46.704 40.177 46.736 40.241 ;
			RECT	47.712 40.177 47.744 40.241 ;
			RECT	49.311 40.177 49.375 40.241 ;
			RECT	49.711 40.177 49.743 40.241 ;
			RECT	50.417 40.177 50.481 40.241 ;
			RECT	50.648 40.177 50.68 40.241 ;
			RECT	51.274 40.177 51.306 40.241 ;
			RECT	51.92 40.177 51.952 40.241 ;
			RECT	52.968 40.177 53.032 40.241 ;
			RECT	53.91 40.177 53.942 40.241 ;
			RECT	54.363 40.177 54.427 40.241 ;
			RECT	54.812 40.177 54.844 40.241 ;
			RECT	55.562 40.177 55.626 40.241 ;
			RECT	55.969 40.177 56.033 40.241 ;
			RECT	56.144 40.177 56.176 40.241 ;
			RECT	56.664 40.177 56.696 40.241 ;
			RECT	57.415 40.177 57.479 40.241 ;
			RECT	57.911 40.177 57.943 40.241 ;
			RECT	58.461 40.177 58.493 40.241 ;
			RECT	58.829 40.177 58.893 40.241 ;
			RECT	60.46 40.177 60.492 40.241 ;
			RECT	61.468 40.177 61.5 40.241 ;
			RECT	62.14 40.177 62.172 40.241 ;
			RECT	63.484 40.177 63.516 40.241 ;
			RECT	64.156 40.177 64.188 40.241 ;
			RECT	64.828 40.177 64.86 40.241 ;
			RECT	67.516 40.177 67.548 40.241 ;
			RECT	67.852 40.177 67.884 40.241 ;
			RECT	68.188 40.177 68.22 40.241 ;
			RECT	68.524 40.177 68.556 40.241 ;
			RECT	69.532 40.177 69.564 40.241 ;
			RECT	70.876 40.177 70.908 40.241 ;
			RECT	73.564 40.177 73.596 40.241 ;
			RECT	73.9 40.177 73.932 40.241 ;
			RECT	74.908 40.177 74.94 40.241 ;
			RECT	76.252 40.177 76.284 40.241 ;
			RECT	77.596 40.177 77.628 40.241 ;
			RECT	78.268 40.177 78.3 40.241 ;
			RECT	78.94 40.177 78.972 40.241 ;
			RECT	79.612 40.177 79.644 40.241 ;
			RECT	80.284 40.177 80.316 40.241 ;
			RECT	102.414 40.177 102.446 40.241 ;
			RECT	103.756 40.177 103.788 40.241 ;
			RECT	125.886 40.177 125.918 40.241 ;
			RECT	126.558 40.177 126.59 40.241 ;
			RECT	127.23 40.177 127.262 40.241 ;
			RECT	127.902 40.177 127.934 40.241 ;
			RECT	128.574 40.177 128.606 40.241 ;
			RECT	129.918 40.177 129.95 40.241 ;
			RECT	131.262 40.177 131.294 40.241 ;
			RECT	132.27 40.177 132.302 40.241 ;
			RECT	132.606 40.177 132.638 40.241 ;
			RECT	135.294 40.177 135.326 40.241 ;
			RECT	136.638 40.177 136.67 40.241 ;
			RECT	137.646 40.177 137.678 40.241 ;
			RECT	137.982 40.177 138.014 40.241 ;
			RECT	138.318 40.177 138.35 40.241 ;
			RECT	138.654 40.177 138.686 40.241 ;
			RECT	141.342 40.177 141.374 40.241 ;
			RECT	142.014 40.177 142.046 40.241 ;
			RECT	142.686 40.177 142.718 40.241 ;
			RECT	144.03 40.177 144.062 40.241 ;
			RECT	144.702 40.177 144.734 40.241 ;
			RECT	145.71 40.177 145.742 40.241 ;
			RECT	147.309 40.177 147.373 40.241 ;
			RECT	147.709 40.177 147.741 40.241 ;
			RECT	148.415 40.177 148.479 40.241 ;
			RECT	148.646 40.177 148.678 40.241 ;
			RECT	149.272 40.177 149.304 40.241 ;
			RECT	149.918 40.177 149.95 40.241 ;
			RECT	150.966 40.177 151.03 40.241 ;
			RECT	151.908 40.177 151.94 40.241 ;
			RECT	152.361 40.177 152.425 40.241 ;
			RECT	152.81 40.177 152.842 40.241 ;
			RECT	153.56 40.177 153.624 40.241 ;
			RECT	153.967 40.177 154.031 40.241 ;
			RECT	154.142 40.177 154.174 40.241 ;
			RECT	154.662 40.177 154.694 40.241 ;
			RECT	155.413 40.177 155.477 40.241 ;
			RECT	155.909 40.177 155.941 40.241 ;
			RECT	156.459 40.177 156.491 40.241 ;
			RECT	156.827 40.177 156.891 40.241 ;
			RECT	158.458 40.177 158.49 40.241 ;
			RECT	159.466 40.177 159.498 40.241 ;
			RECT	160.138 40.177 160.17 40.241 ;
			RECT	161.482 40.177 161.514 40.241 ;
			RECT	162.154 40.177 162.186 40.241 ;
			RECT	162.826 40.177 162.858 40.241 ;
			RECT	165.514 40.177 165.546 40.241 ;
			RECT	165.85 40.177 165.882 40.241 ;
			RECT	166.186 40.177 166.218 40.241 ;
			RECT	166.522 40.177 166.554 40.241 ;
			RECT	167.53 40.177 167.562 40.241 ;
			RECT	168.874 40.177 168.906 40.241 ;
			RECT	171.562 40.177 171.594 40.241 ;
			RECT	171.898 40.177 171.93 40.241 ;
			RECT	172.906 40.177 172.938 40.241 ;
			RECT	174.25 40.177 174.282 40.241 ;
			RECT	175.594 40.177 175.626 40.241 ;
			RECT	176.266 40.177 176.298 40.241 ;
			RECT	176.938 40.177 176.97 40.241 ;
			RECT	177.61 40.177 177.642 40.241 ;
			RECT	178.282 40.177 178.314 40.241 ;
			RECT	200.412 40.177 200.444 40.241 ;
			RECT	200.9 40.177 200.932 40.241 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 41.356 201.665 41.446 ;
			LAYER	J3 ;
			RECT	1.661 41.369 1.693 41.433 ;
			RECT	2.323 41.385 2.387 41.417 ;
			RECT	3.451 41.369 3.483 41.433 ;
			RECT	4.354 41.369 4.386 41.433 ;
			RECT	4.61 41.369 4.642 41.433 ;
			RECT	4.805 41.369 4.837 41.433 ;
			RECT	5.567 41.369 5.599 41.433 ;
			RECT	5.758 41.369 5.79 41.433 ;
			RECT	6.389 41.369 6.421 41.433 ;
			RECT	6.725 41.369 6.757 41.433 ;
			RECT	7.061 41.369 7.093 41.433 ;
			RECT	7.397 41.369 7.429 41.433 ;
			RECT	7.733 41.369 7.765 41.433 ;
			RECT	8.069 41.369 8.101 41.433 ;
			RECT	8.405 41.369 8.437 41.433 ;
			RECT	8.741 41.369 8.773 41.433 ;
			RECT	9.077 41.369 9.109 41.433 ;
			RECT	9.413 41.369 9.445 41.433 ;
			RECT	9.749 41.369 9.781 41.433 ;
			RECT	10.085 41.369 10.117 41.433 ;
			RECT	10.421 41.369 10.453 41.433 ;
			RECT	10.757 41.369 10.789 41.433 ;
			RECT	11.093 41.369 11.125 41.433 ;
			RECT	11.429 41.369 11.461 41.433 ;
			RECT	11.765 41.369 11.797 41.433 ;
			RECT	12.101 41.369 12.133 41.433 ;
			RECT	12.437 41.369 12.469 41.433 ;
			RECT	12.773 41.369 12.805 41.433 ;
			RECT	13.109 41.369 13.141 41.433 ;
			RECT	13.445 41.369 13.477 41.433 ;
			RECT	13.781 41.369 13.813 41.433 ;
			RECT	14.117 41.369 14.149 41.433 ;
			RECT	14.453 41.369 14.485 41.433 ;
			RECT	14.789 41.369 14.821 41.433 ;
			RECT	15.125 41.369 15.157 41.433 ;
			RECT	15.461 41.369 15.493 41.433 ;
			RECT	15.797 41.369 15.829 41.433 ;
			RECT	16.133 41.369 16.165 41.433 ;
			RECT	16.469 41.369 16.501 41.433 ;
			RECT	16.805 41.369 16.837 41.433 ;
			RECT	17.141 41.369 17.173 41.433 ;
			RECT	17.477 41.369 17.509 41.433 ;
			RECT	17.813 41.369 17.845 41.433 ;
			RECT	18.149 41.369 18.181 41.433 ;
			RECT	18.485 41.369 18.517 41.433 ;
			RECT	18.821 41.369 18.853 41.433 ;
			RECT	19.157 41.369 19.189 41.433 ;
			RECT	19.493 41.369 19.525 41.433 ;
			RECT	19.829 41.369 19.861 41.433 ;
			RECT	20.165 41.369 20.197 41.433 ;
			RECT	20.501 41.369 20.533 41.433 ;
			RECT	20.837 41.369 20.869 41.433 ;
			RECT	21.173 41.369 21.205 41.433 ;
			RECT	21.509 41.369 21.541 41.433 ;
			RECT	21.845 41.369 21.877 41.433 ;
			RECT	22.181 41.369 22.213 41.433 ;
			RECT	22.517 41.369 22.549 41.433 ;
			RECT	22.853 41.369 22.885 41.433 ;
			RECT	23.189 41.369 23.221 41.433 ;
			RECT	23.525 41.369 23.557 41.433 ;
			RECT	23.861 41.369 23.893 41.433 ;
			RECT	24.197 41.369 24.229 41.433 ;
			RECT	24.533 41.369 24.565 41.433 ;
			RECT	24.869 41.369 24.901 41.433 ;
			RECT	25.205 41.369 25.237 41.433 ;
			RECT	25.541 41.369 25.573 41.433 ;
			RECT	25.877 41.369 25.909 41.433 ;
			RECT	26.213 41.369 26.245 41.433 ;
			RECT	26.549 41.369 26.581 41.433 ;
			RECT	26.885 41.369 26.917 41.433 ;
			RECT	27.221 41.369 27.253 41.433 ;
			RECT	27.557 41.369 27.589 41.433 ;
			RECT	27.888 41.369 27.92 41.433 ;
			RECT	28.56 41.369 28.592 41.433 ;
			RECT	29.232 41.369 29.264 41.433 ;
			RECT	29.568 41.369 29.6 41.433 ;
			RECT	29.904 41.369 29.936 41.433 ;
			RECT	30.24 41.369 30.272 41.433 ;
			RECT	30.576 41.369 30.608 41.433 ;
			RECT	30.912 41.369 30.944 41.433 ;
			RECT	31.584 41.369 31.616 41.433 ;
			RECT	31.92 41.369 31.952 41.433 ;
			RECT	33.264 41.369 33.296 41.433 ;
			RECT	34.272 41.369 34.304 41.433 ;
			RECT	34.608 41.369 34.64 41.433 ;
			RECT	35.616 41.369 35.648 41.433 ;
			RECT	36.288 41.369 36.32 41.433 ;
			RECT	36.96 41.369 36.992 41.433 ;
			RECT	37.296 41.369 37.328 41.433 ;
			RECT	37.632 41.369 37.664 41.433 ;
			RECT	37.968 41.369 38 41.433 ;
			RECT	39.312 41.369 39.344 41.433 ;
			RECT	39.984 41.369 40.016 41.433 ;
			RECT	40.32 41.369 40.352 41.433 ;
			RECT	41.328 41.369 41.36 41.433 ;
			RECT	41.664 41.369 41.696 41.433 ;
			RECT	42.672 41.369 42.704 41.433 ;
			RECT	44.016 41.369 44.048 41.433 ;
			RECT	44.688 41.369 44.72 41.433 ;
			RECT	45.694 41.369 45.726 41.433 ;
			RECT	46.032 41.369 46.064 41.433 ;
			RECT	46.704 41.369 46.736 41.433 ;
			RECT	47.376 41.369 47.408 41.433 ;
			RECT	47.712 41.369 47.744 41.433 ;
			RECT	48.52 41.385 48.584 41.417 ;
			RECT	49.091 41.369 49.123 41.433 ;
			RECT	49.311 41.385 49.375 41.417 ;
			RECT	50.33 41.369 50.362 41.433 ;
			RECT	50.648 41.369 50.68 41.433 ;
			RECT	51.92 41.369 51.952 41.433 ;
			RECT	52.968 41.385 53.032 41.417 ;
			RECT	53.91 41.385 53.942 41.417 ;
			RECT	54.379 41.369 54.411 41.433 ;
			RECT	54.812 41.369 54.844 41.433 ;
			RECT	55.562 41.385 55.626 41.417 ;
			RECT	55.985 41.369 56.017 41.433 ;
			RECT	57.363 41.369 57.395 41.433 ;
			RECT	57.911 41.369 57.943 41.433 ;
			RECT	58.829 41.385 58.893 41.417 ;
			RECT	59.081 41.369 59.113 41.433 ;
			RECT	59.62 41.385 59.684 41.417 ;
			RECT	60.46 41.369 60.492 41.433 ;
			RECT	60.796 41.369 60.828 41.433 ;
			RECT	61.468 41.369 61.5 41.433 ;
			RECT	62.14 41.369 62.172 41.433 ;
			RECT	62.478 41.369 62.51 41.433 ;
			RECT	63.484 41.369 63.516 41.433 ;
			RECT	64.156 41.369 64.188 41.433 ;
			RECT	65.5 41.369 65.532 41.433 ;
			RECT	66.508 41.369 66.54 41.433 ;
			RECT	66.844 41.369 66.876 41.433 ;
			RECT	67.852 41.369 67.884 41.433 ;
			RECT	68.188 41.369 68.22 41.433 ;
			RECT	68.86 41.369 68.892 41.433 ;
			RECT	70.204 41.369 70.236 41.433 ;
			RECT	70.54 41.369 70.572 41.433 ;
			RECT	70.876 41.369 70.908 41.433 ;
			RECT	71.212 41.369 71.244 41.433 ;
			RECT	71.884 41.369 71.916 41.433 ;
			RECT	72.556 41.369 72.588 41.433 ;
			RECT	73.564 41.369 73.596 41.433 ;
			RECT	73.9 41.369 73.932 41.433 ;
			RECT	74.908 41.369 74.94 41.433 ;
			RECT	76.252 41.369 76.284 41.433 ;
			RECT	76.588 41.369 76.62 41.433 ;
			RECT	77.26 41.369 77.292 41.433 ;
			RECT	77.596 41.369 77.628 41.433 ;
			RECT	77.932 41.369 77.964 41.433 ;
			RECT	78.268 41.369 78.3 41.433 ;
			RECT	78.604 41.369 78.636 41.433 ;
			RECT	78.94 41.369 78.972 41.433 ;
			RECT	79.612 41.369 79.644 41.433 ;
			RECT	80.284 41.369 80.316 41.433 ;
			RECT	80.615 41.369 80.647 41.433 ;
			RECT	80.951 41.369 80.983 41.433 ;
			RECT	81.287 41.369 81.319 41.433 ;
			RECT	81.623 41.369 81.655 41.433 ;
			RECT	81.959 41.369 81.991 41.433 ;
			RECT	82.295 41.369 82.327 41.433 ;
			RECT	82.631 41.369 82.663 41.433 ;
			RECT	82.967 41.369 82.999 41.433 ;
			RECT	83.303 41.369 83.335 41.433 ;
			RECT	83.639 41.369 83.671 41.433 ;
			RECT	83.975 41.369 84.007 41.433 ;
			RECT	84.311 41.369 84.343 41.433 ;
			RECT	84.647 41.369 84.679 41.433 ;
			RECT	84.983 41.369 85.015 41.433 ;
			RECT	85.319 41.369 85.351 41.433 ;
			RECT	85.655 41.369 85.687 41.433 ;
			RECT	85.991 41.369 86.023 41.433 ;
			RECT	86.327 41.369 86.359 41.433 ;
			RECT	86.663 41.369 86.695 41.433 ;
			RECT	86.999 41.369 87.031 41.433 ;
			RECT	87.335 41.369 87.367 41.433 ;
			RECT	87.671 41.369 87.703 41.433 ;
			RECT	88.007 41.369 88.039 41.433 ;
			RECT	88.343 41.369 88.375 41.433 ;
			RECT	88.679 41.369 88.711 41.433 ;
			RECT	89.015 41.369 89.047 41.433 ;
			RECT	89.351 41.369 89.383 41.433 ;
			RECT	89.687 41.369 89.719 41.433 ;
			RECT	90.023 41.369 90.055 41.433 ;
			RECT	90.359 41.369 90.391 41.433 ;
			RECT	90.695 41.369 90.727 41.433 ;
			RECT	91.031 41.369 91.063 41.433 ;
			RECT	91.367 41.369 91.399 41.433 ;
			RECT	91.703 41.369 91.735 41.433 ;
			RECT	92.039 41.369 92.071 41.433 ;
			RECT	92.375 41.369 92.407 41.433 ;
			RECT	92.711 41.369 92.743 41.433 ;
			RECT	93.047 41.369 93.079 41.433 ;
			RECT	93.383 41.369 93.415 41.433 ;
			RECT	93.719 41.369 93.751 41.433 ;
			RECT	94.055 41.369 94.087 41.433 ;
			RECT	94.391 41.369 94.423 41.433 ;
			RECT	94.727 41.369 94.759 41.433 ;
			RECT	95.063 41.369 95.095 41.433 ;
			RECT	95.399 41.369 95.431 41.433 ;
			RECT	95.735 41.369 95.767 41.433 ;
			RECT	96.071 41.369 96.103 41.433 ;
			RECT	96.407 41.369 96.439 41.433 ;
			RECT	96.743 41.369 96.775 41.433 ;
			RECT	97.079 41.369 97.111 41.433 ;
			RECT	97.415 41.369 97.447 41.433 ;
			RECT	97.751 41.369 97.783 41.433 ;
			RECT	98.087 41.369 98.119 41.433 ;
			RECT	98.423 41.369 98.455 41.433 ;
			RECT	98.759 41.369 98.791 41.433 ;
			RECT	99.095 41.369 99.127 41.433 ;
			RECT	99.431 41.369 99.463 41.433 ;
			RECT	99.767 41.369 99.799 41.433 ;
			RECT	100.103 41.369 100.135 41.433 ;
			RECT	100.439 41.369 100.471 41.433 ;
			RECT	100.775 41.369 100.807 41.433 ;
			RECT	101.111 41.369 101.143 41.433 ;
			RECT	101.447 41.369 101.479 41.433 ;
			RECT	101.783 41.369 101.815 41.433 ;
			RECT	102.414 41.369 102.446 41.433 ;
			RECT	102.605 41.369 102.637 41.433 ;
			RECT	103.565 41.369 103.597 41.433 ;
			RECT	103.756 41.369 103.788 41.433 ;
			RECT	104.387 41.369 104.419 41.433 ;
			RECT	104.723 41.369 104.755 41.433 ;
			RECT	105.059 41.369 105.091 41.433 ;
			RECT	105.395 41.369 105.427 41.433 ;
			RECT	105.731 41.369 105.763 41.433 ;
			RECT	106.067 41.369 106.099 41.433 ;
			RECT	106.403 41.369 106.435 41.433 ;
			RECT	106.739 41.369 106.771 41.433 ;
			RECT	107.075 41.369 107.107 41.433 ;
			RECT	107.411 41.369 107.443 41.433 ;
			RECT	107.747 41.369 107.779 41.433 ;
			RECT	108.083 41.369 108.115 41.433 ;
			RECT	108.419 41.369 108.451 41.433 ;
			RECT	108.755 41.369 108.787 41.433 ;
			RECT	109.091 41.369 109.123 41.433 ;
			RECT	109.427 41.369 109.459 41.433 ;
			RECT	109.763 41.369 109.795 41.433 ;
			RECT	110.099 41.369 110.131 41.433 ;
			RECT	110.435 41.369 110.467 41.433 ;
			RECT	110.771 41.369 110.803 41.433 ;
			RECT	111.107 41.369 111.139 41.433 ;
			RECT	111.443 41.369 111.475 41.433 ;
			RECT	111.779 41.369 111.811 41.433 ;
			RECT	112.115 41.369 112.147 41.433 ;
			RECT	112.451 41.369 112.483 41.433 ;
			RECT	112.787 41.369 112.819 41.433 ;
			RECT	113.123 41.369 113.155 41.433 ;
			RECT	113.459 41.369 113.491 41.433 ;
			RECT	113.795 41.369 113.827 41.433 ;
			RECT	114.131 41.369 114.163 41.433 ;
			RECT	114.467 41.369 114.499 41.433 ;
			RECT	114.803 41.369 114.835 41.433 ;
			RECT	115.139 41.369 115.171 41.433 ;
			RECT	115.475 41.369 115.507 41.433 ;
			RECT	115.811 41.369 115.843 41.433 ;
			RECT	116.147 41.369 116.179 41.433 ;
			RECT	116.483 41.369 116.515 41.433 ;
			RECT	116.819 41.369 116.851 41.433 ;
			RECT	117.155 41.369 117.187 41.433 ;
			RECT	117.491 41.369 117.523 41.433 ;
			RECT	117.827 41.369 117.859 41.433 ;
			RECT	118.163 41.369 118.195 41.433 ;
			RECT	118.499 41.369 118.531 41.433 ;
			RECT	118.835 41.369 118.867 41.433 ;
			RECT	119.171 41.369 119.203 41.433 ;
			RECT	119.507 41.369 119.539 41.433 ;
			RECT	119.843 41.369 119.875 41.433 ;
			RECT	120.179 41.369 120.211 41.433 ;
			RECT	120.515 41.369 120.547 41.433 ;
			RECT	120.851 41.369 120.883 41.433 ;
			RECT	121.187 41.369 121.219 41.433 ;
			RECT	121.523 41.369 121.555 41.433 ;
			RECT	121.859 41.369 121.891 41.433 ;
			RECT	122.195 41.369 122.227 41.433 ;
			RECT	122.531 41.369 122.563 41.433 ;
			RECT	122.867 41.369 122.899 41.433 ;
			RECT	123.203 41.369 123.235 41.433 ;
			RECT	123.539 41.369 123.571 41.433 ;
			RECT	123.875 41.369 123.907 41.433 ;
			RECT	124.211 41.369 124.243 41.433 ;
			RECT	124.547 41.369 124.579 41.433 ;
			RECT	124.883 41.369 124.915 41.433 ;
			RECT	125.219 41.369 125.251 41.433 ;
			RECT	125.555 41.369 125.587 41.433 ;
			RECT	125.886 41.369 125.918 41.433 ;
			RECT	126.558 41.369 126.59 41.433 ;
			RECT	127.23 41.369 127.262 41.433 ;
			RECT	127.566 41.369 127.598 41.433 ;
			RECT	127.902 41.369 127.934 41.433 ;
			RECT	128.238 41.369 128.27 41.433 ;
			RECT	128.574 41.369 128.606 41.433 ;
			RECT	128.91 41.369 128.942 41.433 ;
			RECT	129.582 41.369 129.614 41.433 ;
			RECT	129.918 41.369 129.95 41.433 ;
			RECT	131.262 41.369 131.294 41.433 ;
			RECT	132.27 41.369 132.302 41.433 ;
			RECT	132.606 41.369 132.638 41.433 ;
			RECT	133.614 41.369 133.646 41.433 ;
			RECT	134.286 41.369 134.318 41.433 ;
			RECT	134.958 41.369 134.99 41.433 ;
			RECT	135.294 41.369 135.326 41.433 ;
			RECT	135.63 41.369 135.662 41.433 ;
			RECT	135.966 41.369 135.998 41.433 ;
			RECT	137.31 41.369 137.342 41.433 ;
			RECT	137.982 41.369 138.014 41.433 ;
			RECT	138.318 41.369 138.35 41.433 ;
			RECT	139.326 41.369 139.358 41.433 ;
			RECT	139.662 41.369 139.694 41.433 ;
			RECT	140.67 41.369 140.702 41.433 ;
			RECT	142.014 41.369 142.046 41.433 ;
			RECT	142.686 41.369 142.718 41.433 ;
			RECT	143.692 41.369 143.724 41.433 ;
			RECT	144.03 41.369 144.062 41.433 ;
			RECT	144.702 41.369 144.734 41.433 ;
			RECT	145.374 41.369 145.406 41.433 ;
			RECT	145.71 41.369 145.742 41.433 ;
			RECT	146.518 41.385 146.582 41.417 ;
			RECT	147.089 41.369 147.121 41.433 ;
			RECT	147.309 41.385 147.373 41.417 ;
			RECT	148.328 41.369 148.36 41.433 ;
			RECT	148.646 41.369 148.678 41.433 ;
			RECT	149.918 41.369 149.95 41.433 ;
			RECT	150.966 41.385 151.03 41.417 ;
			RECT	151.908 41.385 151.94 41.417 ;
			RECT	152.377 41.369 152.409 41.433 ;
			RECT	152.81 41.369 152.842 41.433 ;
			RECT	153.56 41.385 153.624 41.417 ;
			RECT	153.983 41.369 154.015 41.433 ;
			RECT	155.361 41.369 155.393 41.433 ;
			RECT	155.909 41.369 155.941 41.433 ;
			RECT	156.827 41.385 156.891 41.417 ;
			RECT	157.079 41.369 157.111 41.433 ;
			RECT	157.618 41.385 157.682 41.417 ;
			RECT	158.458 41.369 158.49 41.433 ;
			RECT	158.794 41.369 158.826 41.433 ;
			RECT	159.466 41.369 159.498 41.433 ;
			RECT	160.138 41.369 160.17 41.433 ;
			RECT	160.476 41.369 160.508 41.433 ;
			RECT	161.482 41.369 161.514 41.433 ;
			RECT	162.154 41.369 162.186 41.433 ;
			RECT	163.498 41.369 163.53 41.433 ;
			RECT	164.506 41.369 164.538 41.433 ;
			RECT	164.842 41.369 164.874 41.433 ;
			RECT	165.85 41.369 165.882 41.433 ;
			RECT	166.186 41.369 166.218 41.433 ;
			RECT	166.858 41.369 166.89 41.433 ;
			RECT	168.202 41.369 168.234 41.433 ;
			RECT	168.538 41.369 168.57 41.433 ;
			RECT	168.874 41.369 168.906 41.433 ;
			RECT	169.21 41.369 169.242 41.433 ;
			RECT	169.882 41.369 169.914 41.433 ;
			RECT	170.554 41.369 170.586 41.433 ;
			RECT	171.562 41.369 171.594 41.433 ;
			RECT	171.898 41.369 171.93 41.433 ;
			RECT	172.906 41.369 172.938 41.433 ;
			RECT	174.25 41.369 174.282 41.433 ;
			RECT	174.586 41.369 174.618 41.433 ;
			RECT	175.258 41.369 175.29 41.433 ;
			RECT	175.594 41.369 175.626 41.433 ;
			RECT	175.93 41.369 175.962 41.433 ;
			RECT	176.266 41.369 176.298 41.433 ;
			RECT	176.602 41.369 176.634 41.433 ;
			RECT	176.938 41.369 176.97 41.433 ;
			RECT	177.61 41.369 177.642 41.433 ;
			RECT	178.282 41.369 178.314 41.433 ;
			RECT	178.613 41.369 178.645 41.433 ;
			RECT	178.949 41.369 178.981 41.433 ;
			RECT	179.285 41.369 179.317 41.433 ;
			RECT	179.621 41.369 179.653 41.433 ;
			RECT	179.957 41.369 179.989 41.433 ;
			RECT	180.293 41.369 180.325 41.433 ;
			RECT	180.629 41.369 180.661 41.433 ;
			RECT	180.965 41.369 180.997 41.433 ;
			RECT	181.301 41.369 181.333 41.433 ;
			RECT	181.637 41.369 181.669 41.433 ;
			RECT	181.973 41.369 182.005 41.433 ;
			RECT	182.309 41.369 182.341 41.433 ;
			RECT	182.645 41.369 182.677 41.433 ;
			RECT	182.981 41.369 183.013 41.433 ;
			RECT	183.317 41.369 183.349 41.433 ;
			RECT	183.653 41.369 183.685 41.433 ;
			RECT	183.989 41.369 184.021 41.433 ;
			RECT	184.325 41.369 184.357 41.433 ;
			RECT	184.661 41.369 184.693 41.433 ;
			RECT	184.997 41.369 185.029 41.433 ;
			RECT	185.333 41.369 185.365 41.433 ;
			RECT	185.669 41.369 185.701 41.433 ;
			RECT	186.005 41.369 186.037 41.433 ;
			RECT	186.341 41.369 186.373 41.433 ;
			RECT	186.677 41.369 186.709 41.433 ;
			RECT	187.013 41.369 187.045 41.433 ;
			RECT	187.349 41.369 187.381 41.433 ;
			RECT	187.685 41.369 187.717 41.433 ;
			RECT	188.021 41.369 188.053 41.433 ;
			RECT	188.357 41.369 188.389 41.433 ;
			RECT	188.693 41.369 188.725 41.433 ;
			RECT	189.029 41.369 189.061 41.433 ;
			RECT	189.365 41.369 189.397 41.433 ;
			RECT	189.701 41.369 189.733 41.433 ;
			RECT	190.037 41.369 190.069 41.433 ;
			RECT	190.373 41.369 190.405 41.433 ;
			RECT	190.709 41.369 190.741 41.433 ;
			RECT	191.045 41.369 191.077 41.433 ;
			RECT	191.381 41.369 191.413 41.433 ;
			RECT	191.717 41.369 191.749 41.433 ;
			RECT	192.053 41.369 192.085 41.433 ;
			RECT	192.389 41.369 192.421 41.433 ;
			RECT	192.725 41.369 192.757 41.433 ;
			RECT	193.061 41.369 193.093 41.433 ;
			RECT	193.397 41.369 193.429 41.433 ;
			RECT	193.733 41.369 193.765 41.433 ;
			RECT	194.069 41.369 194.101 41.433 ;
			RECT	194.405 41.369 194.437 41.433 ;
			RECT	194.741 41.369 194.773 41.433 ;
			RECT	195.077 41.369 195.109 41.433 ;
			RECT	195.413 41.369 195.445 41.433 ;
			RECT	195.749 41.369 195.781 41.433 ;
			RECT	196.085 41.369 196.117 41.433 ;
			RECT	196.421 41.369 196.453 41.433 ;
			RECT	196.757 41.369 196.789 41.433 ;
			RECT	197.093 41.369 197.125 41.433 ;
			RECT	197.429 41.369 197.461 41.433 ;
			RECT	197.765 41.369 197.797 41.433 ;
			RECT	198.101 41.369 198.133 41.433 ;
			RECT	198.437 41.369 198.469 41.433 ;
			RECT	198.773 41.369 198.805 41.433 ;
			RECT	199.109 41.369 199.141 41.433 ;
			RECT	199.445 41.369 199.477 41.433 ;
			RECT	199.781 41.369 199.813 41.433 ;
			RECT	200.412 41.369 200.444 41.433 ;
			RECT	200.603 41.369 200.635 41.433 ;
			RECT	200.9 41.369 200.932 41.433 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 42.251 201.665 42.341 ;
			LAYER	J3 ;
			RECT	1.661 42.264 1.693 42.328 ;
			RECT	2.323 42.28 2.387 42.312 ;
			RECT	3.451 42.264 3.483 42.328 ;
			RECT	4.354 42.264 4.386 42.328 ;
			RECT	4.61 42.264 4.642 42.328 ;
			RECT	4.805 42.264 4.837 42.328 ;
			RECT	5.758 42.264 5.79 42.328 ;
			RECT	27.888 42.264 27.92 42.328 ;
			RECT	28.56 42.264 28.592 42.328 ;
			RECT	29.232 42.264 29.264 42.328 ;
			RECT	29.568 42.264 29.6 42.328 ;
			RECT	29.904 42.264 29.936 42.328 ;
			RECT	30.24 42.264 30.272 42.328 ;
			RECT	30.576 42.264 30.608 42.328 ;
			RECT	30.912 42.264 30.944 42.328 ;
			RECT	31.584 42.264 31.616 42.328 ;
			RECT	31.92 42.264 31.952 42.328 ;
			RECT	33.264 42.264 33.296 42.328 ;
			RECT	34.272 42.264 34.304 42.328 ;
			RECT	34.608 42.264 34.64 42.328 ;
			RECT	35.616 42.264 35.648 42.328 ;
			RECT	35.952 42.264 35.984 42.328 ;
			RECT	36.284 42.264 36.316 42.328 ;
			RECT	36.96 42.264 36.992 42.328 ;
			RECT	37.296 42.264 37.328 42.328 ;
			RECT	37.628 42.264 37.66 42.328 ;
			RECT	37.968 42.264 38 42.328 ;
			RECT	38.304 42.264 38.336 42.328 ;
			RECT	38.64 42.264 38.672 42.328 ;
			RECT	39.312 42.264 39.344 42.328 ;
			RECT	39.984 42.264 40.016 42.328 ;
			RECT	40.32 42.264 40.352 42.328 ;
			RECT	41.328 42.264 41.36 42.328 ;
			RECT	42.672 42.264 42.704 42.328 ;
			RECT	44.016 42.264 44.048 42.328 ;
			RECT	44.688 42.264 44.72 42.328 ;
			RECT	45.36 42.264 45.392 42.328 ;
			RECT	46.032 42.264 46.064 42.328 ;
			RECT	48.52 42.28 48.584 42.312 ;
			RECT	49.091 42.264 49.123 42.328 ;
			RECT	49.311 42.28 49.375 42.312 ;
			RECT	49.711 42.264 49.743 42.328 ;
			RECT	50.33 42.264 50.362 42.328 ;
			RECT	51.92 42.264 51.952 42.328 ;
			RECT	52.968 42.28 53.032 42.312 ;
			RECT	53.91 42.264 53.942 42.328 ;
			RECT	54.812 42.264 54.844 42.328 ;
			RECT	55.562 42.28 55.626 42.312 ;
			RECT	55.969 42.28 56.033 42.312 ;
			RECT	58.461 42.264 58.493 42.328 ;
			RECT	58.829 42.28 58.893 42.312 ;
			RECT	59.081 42.264 59.113 42.328 ;
			RECT	59.62 42.28 59.684 42.312 ;
			RECT	62.14 42.264 62.172 42.328 ;
			RECT	62.812 42.264 62.844 42.328 ;
			RECT	63.484 42.264 63.516 42.328 ;
			RECT	64.156 42.264 64.188 42.328 ;
			RECT	65.5 42.264 65.532 42.328 ;
			RECT	66.844 42.264 66.876 42.328 ;
			RECT	67.852 42.264 67.884 42.328 ;
			RECT	68.188 42.264 68.22 42.328 ;
			RECT	68.86 42.264 68.892 42.328 ;
			RECT	69.532 42.264 69.564 42.328 ;
			RECT	69.868 42.264 69.9 42.328 ;
			RECT	70.204 42.264 70.236 42.328 ;
			RECT	70.544 42.264 70.576 42.328 ;
			RECT	70.876 42.264 70.908 42.328 ;
			RECT	71.212 42.264 71.244 42.328 ;
			RECT	71.888 42.264 71.92 42.328 ;
			RECT	72.22 42.264 72.252 42.328 ;
			RECT	72.556 42.264 72.588 42.328 ;
			RECT	73.564 42.264 73.596 42.328 ;
			RECT	73.9 42.264 73.932 42.328 ;
			RECT	74.908 42.264 74.94 42.328 ;
			RECT	76.252 42.264 76.284 42.328 ;
			RECT	76.588 42.264 76.62 42.328 ;
			RECT	77.26 42.264 77.292 42.328 ;
			RECT	77.596 42.264 77.628 42.328 ;
			RECT	77.932 42.264 77.964 42.328 ;
			RECT	78.268 42.264 78.3 42.328 ;
			RECT	78.604 42.264 78.636 42.328 ;
			RECT	78.94 42.264 78.972 42.328 ;
			RECT	79.612 42.264 79.644 42.328 ;
			RECT	80.284 42.264 80.316 42.328 ;
			RECT	102.414 42.264 102.446 42.328 ;
			RECT	103.756 42.264 103.788 42.328 ;
			RECT	125.886 42.264 125.918 42.328 ;
			RECT	126.558 42.264 126.59 42.328 ;
			RECT	127.23 42.264 127.262 42.328 ;
			RECT	127.566 42.264 127.598 42.328 ;
			RECT	127.902 42.264 127.934 42.328 ;
			RECT	128.238 42.264 128.27 42.328 ;
			RECT	128.574 42.264 128.606 42.328 ;
			RECT	128.91 42.264 128.942 42.328 ;
			RECT	129.582 42.264 129.614 42.328 ;
			RECT	129.918 42.264 129.95 42.328 ;
			RECT	131.262 42.264 131.294 42.328 ;
			RECT	132.27 42.264 132.302 42.328 ;
			RECT	132.606 42.264 132.638 42.328 ;
			RECT	133.614 42.264 133.646 42.328 ;
			RECT	133.95 42.264 133.982 42.328 ;
			RECT	134.282 42.264 134.314 42.328 ;
			RECT	134.958 42.264 134.99 42.328 ;
			RECT	135.294 42.264 135.326 42.328 ;
			RECT	135.626 42.264 135.658 42.328 ;
			RECT	135.966 42.264 135.998 42.328 ;
			RECT	136.302 42.264 136.334 42.328 ;
			RECT	136.638 42.264 136.67 42.328 ;
			RECT	137.31 42.264 137.342 42.328 ;
			RECT	137.982 42.264 138.014 42.328 ;
			RECT	138.318 42.264 138.35 42.328 ;
			RECT	139.326 42.264 139.358 42.328 ;
			RECT	140.67 42.264 140.702 42.328 ;
			RECT	142.014 42.264 142.046 42.328 ;
			RECT	142.686 42.264 142.718 42.328 ;
			RECT	143.358 42.264 143.39 42.328 ;
			RECT	144.03 42.264 144.062 42.328 ;
			RECT	146.518 42.28 146.582 42.312 ;
			RECT	147.089 42.264 147.121 42.328 ;
			RECT	147.309 42.28 147.373 42.312 ;
			RECT	147.709 42.264 147.741 42.328 ;
			RECT	148.328 42.264 148.36 42.328 ;
			RECT	149.918 42.264 149.95 42.328 ;
			RECT	150.966 42.28 151.03 42.312 ;
			RECT	151.908 42.264 151.94 42.328 ;
			RECT	152.81 42.264 152.842 42.328 ;
			RECT	153.56 42.28 153.624 42.312 ;
			RECT	153.967 42.28 154.031 42.312 ;
			RECT	156.459 42.264 156.491 42.328 ;
			RECT	156.827 42.28 156.891 42.312 ;
			RECT	157.079 42.264 157.111 42.328 ;
			RECT	157.618 42.28 157.682 42.312 ;
			RECT	160.138 42.264 160.17 42.328 ;
			RECT	160.81 42.264 160.842 42.328 ;
			RECT	161.482 42.264 161.514 42.328 ;
			RECT	162.154 42.264 162.186 42.328 ;
			RECT	163.498 42.264 163.53 42.328 ;
			RECT	164.842 42.264 164.874 42.328 ;
			RECT	165.85 42.264 165.882 42.328 ;
			RECT	166.186 42.264 166.218 42.328 ;
			RECT	166.858 42.264 166.89 42.328 ;
			RECT	167.53 42.264 167.562 42.328 ;
			RECT	167.866 42.264 167.898 42.328 ;
			RECT	168.202 42.264 168.234 42.328 ;
			RECT	168.542 42.264 168.574 42.328 ;
			RECT	168.874 42.264 168.906 42.328 ;
			RECT	169.21 42.264 169.242 42.328 ;
			RECT	169.886 42.264 169.918 42.328 ;
			RECT	170.218 42.264 170.25 42.328 ;
			RECT	170.554 42.264 170.586 42.328 ;
			RECT	171.562 42.264 171.594 42.328 ;
			RECT	171.898 42.264 171.93 42.328 ;
			RECT	172.906 42.264 172.938 42.328 ;
			RECT	174.25 42.264 174.282 42.328 ;
			RECT	174.586 42.264 174.618 42.328 ;
			RECT	175.258 42.264 175.29 42.328 ;
			RECT	175.594 42.264 175.626 42.328 ;
			RECT	175.93 42.264 175.962 42.328 ;
			RECT	176.266 42.264 176.298 42.328 ;
			RECT	176.602 42.264 176.634 42.328 ;
			RECT	176.938 42.264 176.97 42.328 ;
			RECT	177.61 42.264 177.642 42.328 ;
			RECT	178.282 42.264 178.314 42.328 ;
			RECT	200.412 42.264 200.444 42.328 ;
			RECT	200.9 42.264 200.932 42.328 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 43.803 201.665 43.923 ;
			LAYER	J3 ;
			RECT	1.645 43.831 1.709 43.895 ;
			RECT	1.981 43.831 2.013 43.895 ;
			RECT	2.323 43.831 2.387 43.895 ;
			RECT	3.451 43.831 3.483 43.895 ;
			RECT	4.61 43.831 4.642 43.895 ;
			RECT	4.805 43.831 4.837 43.895 ;
			RECT	5.252 43.831 5.284 43.895 ;
			RECT	5.567 43.831 5.599 43.895 ;
			RECT	5.793 43.831 5.825 43.895 ;
			RECT	6.389 43.831 6.421 43.895 ;
			RECT	6.725 43.831 6.757 43.895 ;
			RECT	7.061 43.831 7.093 43.895 ;
			RECT	7.397 43.831 7.429 43.895 ;
			RECT	7.733 43.831 7.765 43.895 ;
			RECT	8.069 43.831 8.101 43.895 ;
			RECT	8.405 43.831 8.437 43.895 ;
			RECT	8.741 43.831 8.773 43.895 ;
			RECT	9.077 43.831 9.109 43.895 ;
			RECT	9.413 43.831 9.445 43.895 ;
			RECT	9.749 43.831 9.781 43.895 ;
			RECT	10.085 43.831 10.117 43.895 ;
			RECT	10.421 43.831 10.453 43.895 ;
			RECT	10.757 43.831 10.789 43.895 ;
			RECT	11.093 43.831 11.125 43.895 ;
			RECT	11.429 43.831 11.461 43.895 ;
			RECT	11.765 43.831 11.797 43.895 ;
			RECT	12.101 43.831 12.133 43.895 ;
			RECT	12.437 43.831 12.469 43.895 ;
			RECT	12.773 43.831 12.805 43.895 ;
			RECT	13.109 43.831 13.141 43.895 ;
			RECT	13.445 43.831 13.477 43.895 ;
			RECT	13.781 43.831 13.813 43.895 ;
			RECT	14.117 43.831 14.149 43.895 ;
			RECT	14.453 43.831 14.485 43.895 ;
			RECT	14.789 43.831 14.821 43.895 ;
			RECT	15.125 43.831 15.157 43.895 ;
			RECT	15.461 43.831 15.493 43.895 ;
			RECT	15.797 43.831 15.829 43.895 ;
			RECT	16.133 43.831 16.165 43.895 ;
			RECT	16.469 43.831 16.501 43.895 ;
			RECT	16.805 43.831 16.837 43.895 ;
			RECT	17.141 43.831 17.173 43.895 ;
			RECT	17.477 43.831 17.509 43.895 ;
			RECT	17.813 43.831 17.845 43.895 ;
			RECT	18.149 43.831 18.181 43.895 ;
			RECT	18.485 43.831 18.517 43.895 ;
			RECT	18.821 43.831 18.853 43.895 ;
			RECT	19.157 43.831 19.189 43.895 ;
			RECT	19.493 43.831 19.525 43.895 ;
			RECT	19.829 43.831 19.861 43.895 ;
			RECT	20.165 43.831 20.197 43.895 ;
			RECT	20.501 43.831 20.533 43.895 ;
			RECT	20.837 43.831 20.869 43.895 ;
			RECT	21.173 43.831 21.205 43.895 ;
			RECT	21.509 43.831 21.541 43.895 ;
			RECT	21.845 43.831 21.877 43.895 ;
			RECT	22.181 43.831 22.213 43.895 ;
			RECT	22.517 43.831 22.549 43.895 ;
			RECT	22.853 43.831 22.885 43.895 ;
			RECT	23.189 43.831 23.221 43.895 ;
			RECT	23.525 43.831 23.557 43.895 ;
			RECT	23.861 43.831 23.893 43.895 ;
			RECT	24.197 43.831 24.229 43.895 ;
			RECT	24.533 43.831 24.565 43.895 ;
			RECT	24.869 43.831 24.901 43.895 ;
			RECT	25.205 43.831 25.237 43.895 ;
			RECT	25.541 43.831 25.573 43.895 ;
			RECT	25.877 43.831 25.909 43.895 ;
			RECT	26.213 43.831 26.245 43.895 ;
			RECT	26.549 43.831 26.581 43.895 ;
			RECT	26.885 43.831 26.917 43.895 ;
			RECT	27.221 43.831 27.253 43.895 ;
			RECT	27.557 43.831 27.589 43.895 ;
			RECT	27.888 43.831 27.92 43.895 ;
			RECT	28.56 43.831 28.592 43.895 ;
			RECT	29.232 43.831 29.264 43.895 ;
			RECT	29.568 43.831 29.6 43.895 ;
			RECT	29.904 43.831 29.936 43.895 ;
			RECT	30.24 43.831 30.272 43.895 ;
			RECT	30.576 43.831 30.608 43.895 ;
			RECT	30.912 43.831 30.944 43.895 ;
			RECT	31.584 43.831 31.616 43.895 ;
			RECT	31.92 43.831 31.952 43.895 ;
			RECT	32.592 43.831 32.624 43.895 ;
			RECT	34.272 43.831 34.304 43.895 ;
			RECT	34.608 43.831 34.64 43.895 ;
			RECT	35.616 43.831 35.648 43.895 ;
			RECT	35.952 43.831 35.984 43.895 ;
			RECT	36.96 43.831 36.992 43.895 ;
			RECT	37.296 43.831 37.328 43.895 ;
			RECT	38.304 43.831 38.336 43.895 ;
			RECT	38.64 43.831 38.672 43.895 ;
			RECT	39.648 43.831 39.68 43.895 ;
			RECT	40.32 43.831 40.352 43.895 ;
			RECT	41.328 43.831 41.36 43.895 ;
			RECT	42.672 43.831 42.704 43.895 ;
			RECT	43.68 43.831 43.712 43.895 ;
			RECT	44.201 43.831 44.233 43.895 ;
			RECT	45.36 43.831 45.392 43.895 ;
			RECT	46.032 43.831 46.064 43.895 ;
			RECT	47.04 43.831 47.072 43.895 ;
			RECT	48.52 43.831 48.584 43.895 ;
			RECT	49.056 43.831 49.088 43.895 ;
			RECT	49.311 43.831 49.375 43.895 ;
			RECT	49.675 43.831 49.707 43.895 ;
			RECT	50.33 43.831 50.362 43.895 ;
			RECT	51.92 43.831 51.952 43.895 ;
			RECT	52.968 43.831 53.032 43.895 ;
			RECT	53.91 43.831 53.942 43.895 ;
			RECT	54.251 43.831 54.283 43.895 ;
			RECT	54.657 43.831 54.689 43.895 ;
			RECT	54.812 43.831 54.844 43.895 ;
			RECT	55.208 43.831 55.272 43.895 ;
			RECT	55.562 43.831 55.626 43.895 ;
			RECT	55.842 43.831 55.874 43.895 ;
			RECT	55.969 43.831 56.033 43.895 ;
			RECT	58.497 43.831 58.529 43.895 ;
			RECT	58.829 43.831 58.893 43.895 ;
			RECT	59.116 43.831 59.148 43.895 ;
			RECT	59.62 43.831 59.684 43.895 ;
			RECT	61.132 43.831 61.164 43.895 ;
			RECT	62.14 43.831 62.172 43.895 ;
			RECT	62.812 43.831 62.844 43.895 ;
			RECT	63.971 43.831 64.003 43.895 ;
			RECT	64.492 43.831 64.524 43.895 ;
			RECT	65.5 43.831 65.532 43.895 ;
			RECT	66.844 43.831 66.876 43.895 ;
			RECT	67.852 43.831 67.884 43.895 ;
			RECT	68.524 43.831 68.556 43.895 ;
			RECT	69.532 43.831 69.564 43.895 ;
			RECT	69.868 43.831 69.9 43.895 ;
			RECT	70.876 43.831 70.908 43.895 ;
			RECT	71.212 43.831 71.244 43.895 ;
			RECT	72.22 43.831 72.252 43.895 ;
			RECT	72.556 43.831 72.588 43.895 ;
			RECT	73.564 43.831 73.596 43.895 ;
			RECT	73.9 43.831 73.932 43.895 ;
			RECT	75.58 43.831 75.612 43.895 ;
			RECT	76.252 43.831 76.284 43.895 ;
			RECT	76.588 43.831 76.62 43.895 ;
			RECT	77.26 43.831 77.292 43.895 ;
			RECT	77.596 43.831 77.628 43.895 ;
			RECT	77.932 43.831 77.964 43.895 ;
			RECT	78.268 43.831 78.3 43.895 ;
			RECT	78.604 43.831 78.636 43.895 ;
			RECT	78.94 43.831 78.972 43.895 ;
			RECT	79.612 43.831 79.644 43.895 ;
			RECT	80.284 43.831 80.316 43.895 ;
			RECT	80.615 43.831 80.647 43.895 ;
			RECT	80.951 43.831 80.983 43.895 ;
			RECT	81.287 43.831 81.319 43.895 ;
			RECT	81.623 43.831 81.655 43.895 ;
			RECT	81.959 43.831 81.991 43.895 ;
			RECT	82.295 43.831 82.327 43.895 ;
			RECT	82.631 43.831 82.663 43.895 ;
			RECT	82.967 43.831 82.999 43.895 ;
			RECT	83.303 43.831 83.335 43.895 ;
			RECT	83.639 43.831 83.671 43.895 ;
			RECT	83.975 43.831 84.007 43.895 ;
			RECT	84.311 43.831 84.343 43.895 ;
			RECT	84.647 43.831 84.679 43.895 ;
			RECT	84.983 43.831 85.015 43.895 ;
			RECT	85.319 43.831 85.351 43.895 ;
			RECT	85.655 43.831 85.687 43.895 ;
			RECT	85.991 43.831 86.023 43.895 ;
			RECT	86.327 43.831 86.359 43.895 ;
			RECT	86.663 43.831 86.695 43.895 ;
			RECT	86.999 43.831 87.031 43.895 ;
			RECT	87.335 43.831 87.367 43.895 ;
			RECT	87.671 43.831 87.703 43.895 ;
			RECT	88.007 43.831 88.039 43.895 ;
			RECT	88.343 43.831 88.375 43.895 ;
			RECT	88.679 43.831 88.711 43.895 ;
			RECT	89.015 43.831 89.047 43.895 ;
			RECT	89.351 43.831 89.383 43.895 ;
			RECT	89.687 43.831 89.719 43.895 ;
			RECT	90.023 43.831 90.055 43.895 ;
			RECT	90.359 43.831 90.391 43.895 ;
			RECT	90.695 43.831 90.727 43.895 ;
			RECT	91.031 43.831 91.063 43.895 ;
			RECT	91.367 43.831 91.399 43.895 ;
			RECT	91.703 43.831 91.735 43.895 ;
			RECT	92.039 43.831 92.071 43.895 ;
			RECT	92.375 43.831 92.407 43.895 ;
			RECT	92.711 43.831 92.743 43.895 ;
			RECT	93.047 43.831 93.079 43.895 ;
			RECT	93.383 43.831 93.415 43.895 ;
			RECT	93.719 43.831 93.751 43.895 ;
			RECT	94.055 43.831 94.087 43.895 ;
			RECT	94.391 43.831 94.423 43.895 ;
			RECT	94.727 43.831 94.759 43.895 ;
			RECT	95.063 43.831 95.095 43.895 ;
			RECT	95.399 43.831 95.431 43.895 ;
			RECT	95.735 43.831 95.767 43.895 ;
			RECT	96.071 43.831 96.103 43.895 ;
			RECT	96.407 43.831 96.439 43.895 ;
			RECT	96.743 43.831 96.775 43.895 ;
			RECT	97.079 43.831 97.111 43.895 ;
			RECT	97.415 43.831 97.447 43.895 ;
			RECT	97.751 43.831 97.783 43.895 ;
			RECT	98.087 43.831 98.119 43.895 ;
			RECT	98.423 43.831 98.455 43.895 ;
			RECT	98.759 43.831 98.791 43.895 ;
			RECT	99.095 43.831 99.127 43.895 ;
			RECT	99.431 43.831 99.463 43.895 ;
			RECT	99.767 43.831 99.799 43.895 ;
			RECT	100.103 43.831 100.135 43.895 ;
			RECT	100.439 43.831 100.471 43.895 ;
			RECT	100.775 43.831 100.807 43.895 ;
			RECT	101.111 43.831 101.143 43.895 ;
			RECT	101.447 43.831 101.479 43.895 ;
			RECT	101.783 43.831 101.815 43.895 ;
			RECT	102.379 43.831 102.411 43.895 ;
			RECT	102.605 43.831 102.637 43.895 ;
			RECT	103.565 43.831 103.597 43.895 ;
			RECT	103.791 43.831 103.823 43.895 ;
			RECT	104.387 43.831 104.419 43.895 ;
			RECT	104.723 43.831 104.755 43.895 ;
			RECT	105.059 43.831 105.091 43.895 ;
			RECT	105.395 43.831 105.427 43.895 ;
			RECT	105.731 43.831 105.763 43.895 ;
			RECT	106.067 43.831 106.099 43.895 ;
			RECT	106.403 43.831 106.435 43.895 ;
			RECT	106.739 43.831 106.771 43.895 ;
			RECT	107.075 43.831 107.107 43.895 ;
			RECT	107.411 43.831 107.443 43.895 ;
			RECT	107.747 43.831 107.779 43.895 ;
			RECT	108.083 43.831 108.115 43.895 ;
			RECT	108.419 43.831 108.451 43.895 ;
			RECT	108.755 43.831 108.787 43.895 ;
			RECT	109.091 43.831 109.123 43.895 ;
			RECT	109.427 43.831 109.459 43.895 ;
			RECT	109.763 43.831 109.795 43.895 ;
			RECT	110.099 43.831 110.131 43.895 ;
			RECT	110.435 43.831 110.467 43.895 ;
			RECT	110.771 43.831 110.803 43.895 ;
			RECT	111.107 43.831 111.139 43.895 ;
			RECT	111.443 43.831 111.475 43.895 ;
			RECT	111.779 43.831 111.811 43.895 ;
			RECT	112.115 43.831 112.147 43.895 ;
			RECT	112.451 43.831 112.483 43.895 ;
			RECT	112.787 43.831 112.819 43.895 ;
			RECT	113.123 43.831 113.155 43.895 ;
			RECT	113.459 43.831 113.491 43.895 ;
			RECT	113.795 43.831 113.827 43.895 ;
			RECT	114.131 43.831 114.163 43.895 ;
			RECT	114.467 43.831 114.499 43.895 ;
			RECT	114.803 43.831 114.835 43.895 ;
			RECT	115.139 43.831 115.171 43.895 ;
			RECT	115.475 43.831 115.507 43.895 ;
			RECT	115.811 43.831 115.843 43.895 ;
			RECT	116.147 43.831 116.179 43.895 ;
			RECT	116.483 43.831 116.515 43.895 ;
			RECT	116.819 43.831 116.851 43.895 ;
			RECT	117.155 43.831 117.187 43.895 ;
			RECT	117.491 43.831 117.523 43.895 ;
			RECT	117.827 43.831 117.859 43.895 ;
			RECT	118.163 43.831 118.195 43.895 ;
			RECT	118.499 43.831 118.531 43.895 ;
			RECT	118.835 43.831 118.867 43.895 ;
			RECT	119.171 43.831 119.203 43.895 ;
			RECT	119.507 43.831 119.539 43.895 ;
			RECT	119.843 43.831 119.875 43.895 ;
			RECT	120.179 43.831 120.211 43.895 ;
			RECT	120.515 43.831 120.547 43.895 ;
			RECT	120.851 43.831 120.883 43.895 ;
			RECT	121.187 43.831 121.219 43.895 ;
			RECT	121.523 43.831 121.555 43.895 ;
			RECT	121.859 43.831 121.891 43.895 ;
			RECT	122.195 43.831 122.227 43.895 ;
			RECT	122.531 43.831 122.563 43.895 ;
			RECT	122.867 43.831 122.899 43.895 ;
			RECT	123.203 43.831 123.235 43.895 ;
			RECT	123.539 43.831 123.571 43.895 ;
			RECT	123.875 43.831 123.907 43.895 ;
			RECT	124.211 43.831 124.243 43.895 ;
			RECT	124.547 43.831 124.579 43.895 ;
			RECT	124.883 43.831 124.915 43.895 ;
			RECT	125.219 43.831 125.251 43.895 ;
			RECT	125.555 43.831 125.587 43.895 ;
			RECT	125.886 43.831 125.918 43.895 ;
			RECT	126.558 43.831 126.59 43.895 ;
			RECT	127.23 43.831 127.262 43.895 ;
			RECT	127.566 43.831 127.598 43.895 ;
			RECT	127.902 43.831 127.934 43.895 ;
			RECT	128.238 43.831 128.27 43.895 ;
			RECT	128.574 43.831 128.606 43.895 ;
			RECT	128.91 43.831 128.942 43.895 ;
			RECT	129.582 43.831 129.614 43.895 ;
			RECT	129.918 43.831 129.95 43.895 ;
			RECT	130.59 43.831 130.622 43.895 ;
			RECT	132.27 43.831 132.302 43.895 ;
			RECT	132.606 43.831 132.638 43.895 ;
			RECT	133.614 43.831 133.646 43.895 ;
			RECT	133.95 43.831 133.982 43.895 ;
			RECT	134.958 43.831 134.99 43.895 ;
			RECT	135.294 43.831 135.326 43.895 ;
			RECT	136.302 43.831 136.334 43.895 ;
			RECT	136.638 43.831 136.67 43.895 ;
			RECT	137.646 43.831 137.678 43.895 ;
			RECT	138.318 43.831 138.35 43.895 ;
			RECT	139.326 43.831 139.358 43.895 ;
			RECT	140.67 43.831 140.702 43.895 ;
			RECT	141.678 43.831 141.71 43.895 ;
			RECT	142.199 43.831 142.231 43.895 ;
			RECT	143.358 43.831 143.39 43.895 ;
			RECT	144.03 43.831 144.062 43.895 ;
			RECT	145.038 43.831 145.07 43.895 ;
			RECT	146.518 43.831 146.582 43.895 ;
			RECT	147.054 43.831 147.086 43.895 ;
			RECT	147.309 43.831 147.373 43.895 ;
			RECT	147.673 43.831 147.705 43.895 ;
			RECT	148.328 43.831 148.36 43.895 ;
			RECT	149.918 43.831 149.95 43.895 ;
			RECT	150.966 43.831 151.03 43.895 ;
			RECT	151.908 43.831 151.94 43.895 ;
			RECT	152.249 43.831 152.281 43.895 ;
			RECT	152.655 43.831 152.687 43.895 ;
			RECT	152.81 43.831 152.842 43.895 ;
			RECT	153.206 43.831 153.27 43.895 ;
			RECT	153.56 43.831 153.624 43.895 ;
			RECT	153.84 43.831 153.872 43.895 ;
			RECT	153.967 43.831 154.031 43.895 ;
			RECT	156.495 43.831 156.527 43.895 ;
			RECT	156.827 43.831 156.891 43.895 ;
			RECT	157.114 43.831 157.146 43.895 ;
			RECT	157.618 43.831 157.682 43.895 ;
			RECT	159.13 43.831 159.162 43.895 ;
			RECT	160.138 43.831 160.17 43.895 ;
			RECT	160.81 43.831 160.842 43.895 ;
			RECT	161.969 43.831 162.001 43.895 ;
			RECT	162.49 43.831 162.522 43.895 ;
			RECT	163.498 43.831 163.53 43.895 ;
			RECT	164.842 43.831 164.874 43.895 ;
			RECT	165.85 43.831 165.882 43.895 ;
			RECT	166.522 43.831 166.554 43.895 ;
			RECT	167.53 43.831 167.562 43.895 ;
			RECT	167.866 43.831 167.898 43.895 ;
			RECT	168.874 43.831 168.906 43.895 ;
			RECT	169.21 43.831 169.242 43.895 ;
			RECT	170.218 43.831 170.25 43.895 ;
			RECT	170.554 43.831 170.586 43.895 ;
			RECT	171.562 43.831 171.594 43.895 ;
			RECT	171.898 43.831 171.93 43.895 ;
			RECT	173.578 43.831 173.61 43.895 ;
			RECT	174.25 43.831 174.282 43.895 ;
			RECT	174.586 43.831 174.618 43.895 ;
			RECT	175.258 43.831 175.29 43.895 ;
			RECT	175.594 43.831 175.626 43.895 ;
			RECT	175.93 43.831 175.962 43.895 ;
			RECT	176.266 43.831 176.298 43.895 ;
			RECT	176.602 43.831 176.634 43.895 ;
			RECT	176.938 43.831 176.97 43.895 ;
			RECT	177.61 43.831 177.642 43.895 ;
			RECT	178.282 43.831 178.314 43.895 ;
			RECT	178.613 43.831 178.645 43.895 ;
			RECT	178.949 43.831 178.981 43.895 ;
			RECT	179.285 43.831 179.317 43.895 ;
			RECT	179.621 43.831 179.653 43.895 ;
			RECT	179.957 43.831 179.989 43.895 ;
			RECT	180.293 43.831 180.325 43.895 ;
			RECT	180.629 43.831 180.661 43.895 ;
			RECT	180.965 43.831 180.997 43.895 ;
			RECT	181.301 43.831 181.333 43.895 ;
			RECT	181.637 43.831 181.669 43.895 ;
			RECT	181.973 43.831 182.005 43.895 ;
			RECT	182.309 43.831 182.341 43.895 ;
			RECT	182.645 43.831 182.677 43.895 ;
			RECT	182.981 43.831 183.013 43.895 ;
			RECT	183.317 43.831 183.349 43.895 ;
			RECT	183.653 43.831 183.685 43.895 ;
			RECT	183.989 43.831 184.021 43.895 ;
			RECT	184.325 43.831 184.357 43.895 ;
			RECT	184.661 43.831 184.693 43.895 ;
			RECT	184.997 43.831 185.029 43.895 ;
			RECT	185.333 43.831 185.365 43.895 ;
			RECT	185.669 43.831 185.701 43.895 ;
			RECT	186.005 43.831 186.037 43.895 ;
			RECT	186.341 43.831 186.373 43.895 ;
			RECT	186.677 43.831 186.709 43.895 ;
			RECT	187.013 43.831 187.045 43.895 ;
			RECT	187.349 43.831 187.381 43.895 ;
			RECT	187.685 43.831 187.717 43.895 ;
			RECT	188.021 43.831 188.053 43.895 ;
			RECT	188.357 43.831 188.389 43.895 ;
			RECT	188.693 43.831 188.725 43.895 ;
			RECT	189.029 43.831 189.061 43.895 ;
			RECT	189.365 43.831 189.397 43.895 ;
			RECT	189.701 43.831 189.733 43.895 ;
			RECT	190.037 43.831 190.069 43.895 ;
			RECT	190.373 43.831 190.405 43.895 ;
			RECT	190.709 43.831 190.741 43.895 ;
			RECT	191.045 43.831 191.077 43.895 ;
			RECT	191.381 43.831 191.413 43.895 ;
			RECT	191.717 43.831 191.749 43.895 ;
			RECT	192.053 43.831 192.085 43.895 ;
			RECT	192.389 43.831 192.421 43.895 ;
			RECT	192.725 43.831 192.757 43.895 ;
			RECT	193.061 43.831 193.093 43.895 ;
			RECT	193.397 43.831 193.429 43.895 ;
			RECT	193.733 43.831 193.765 43.895 ;
			RECT	194.069 43.831 194.101 43.895 ;
			RECT	194.405 43.831 194.437 43.895 ;
			RECT	194.741 43.831 194.773 43.895 ;
			RECT	195.077 43.831 195.109 43.895 ;
			RECT	195.413 43.831 195.445 43.895 ;
			RECT	195.749 43.831 195.781 43.895 ;
			RECT	196.085 43.831 196.117 43.895 ;
			RECT	196.421 43.831 196.453 43.895 ;
			RECT	196.757 43.831 196.789 43.895 ;
			RECT	197.093 43.831 197.125 43.895 ;
			RECT	197.429 43.831 197.461 43.895 ;
			RECT	197.765 43.831 197.797 43.895 ;
			RECT	198.101 43.831 198.133 43.895 ;
			RECT	198.437 43.831 198.469 43.895 ;
			RECT	198.773 43.831 198.805 43.895 ;
			RECT	199.109 43.831 199.141 43.895 ;
			RECT	199.445 43.831 199.477 43.895 ;
			RECT	199.781 43.831 199.813 43.895 ;
			RECT	200.377 43.831 200.409 43.895 ;
			RECT	200.603 43.831 200.635 43.895 ;
			RECT	200.9 43.831 200.932 43.895 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 44.979 201.665 45.069 ;
			LAYER	J3 ;
			RECT	1.661 44.992 1.693 45.056 ;
			RECT	1.981 44.992 2.013 45.056 ;
			RECT	2.323 45.008 2.387 45.04 ;
			RECT	3.451 44.992 3.483 45.056 ;
			RECT	4.347 44.992 4.379 45.056 ;
			RECT	4.568 45.008 4.632 45.04 ;
			RECT	4.805 44.991 4.837 45.055 ;
			RECT	5.252 44.992 5.284 45.056 ;
			RECT	5.567 44.992 5.599 45.056 ;
			RECT	5.793 44.992 5.825 45.056 ;
			RECT	6.389 44.992 6.421 45.056 ;
			RECT	6.725 44.992 6.757 45.056 ;
			RECT	7.061 44.992 7.093 45.056 ;
			RECT	7.397 44.992 7.429 45.056 ;
			RECT	7.733 44.992 7.765 45.056 ;
			RECT	8.069 44.992 8.101 45.056 ;
			RECT	8.405 44.992 8.437 45.056 ;
			RECT	8.741 44.992 8.773 45.056 ;
			RECT	9.077 44.992 9.109 45.056 ;
			RECT	9.413 44.992 9.445 45.056 ;
			RECT	9.749 44.992 9.781 45.056 ;
			RECT	10.085 44.992 10.117 45.056 ;
			RECT	10.421 44.992 10.453 45.056 ;
			RECT	10.757 44.992 10.789 45.056 ;
			RECT	11.093 44.992 11.125 45.056 ;
			RECT	11.429 44.992 11.461 45.056 ;
			RECT	11.765 44.992 11.797 45.056 ;
			RECT	12.101 44.992 12.133 45.056 ;
			RECT	12.437 44.992 12.469 45.056 ;
			RECT	12.773 44.992 12.805 45.056 ;
			RECT	13.109 44.992 13.141 45.056 ;
			RECT	13.445 44.992 13.477 45.056 ;
			RECT	13.781 44.992 13.813 45.056 ;
			RECT	14.117 44.992 14.149 45.056 ;
			RECT	14.453 44.992 14.485 45.056 ;
			RECT	14.789 44.992 14.821 45.056 ;
			RECT	15.125 44.992 15.157 45.056 ;
			RECT	15.461 44.992 15.493 45.056 ;
			RECT	15.797 44.992 15.829 45.056 ;
			RECT	16.133 44.992 16.165 45.056 ;
			RECT	16.469 44.992 16.501 45.056 ;
			RECT	16.805 44.992 16.837 45.056 ;
			RECT	17.141 44.992 17.173 45.056 ;
			RECT	17.477 44.992 17.509 45.056 ;
			RECT	17.813 44.992 17.845 45.056 ;
			RECT	18.149 44.992 18.181 45.056 ;
			RECT	18.485 44.992 18.517 45.056 ;
			RECT	18.821 44.992 18.853 45.056 ;
			RECT	19.157 44.992 19.189 45.056 ;
			RECT	19.493 44.992 19.525 45.056 ;
			RECT	19.829 44.992 19.861 45.056 ;
			RECT	20.165 44.992 20.197 45.056 ;
			RECT	20.501 44.992 20.533 45.056 ;
			RECT	20.837 44.992 20.869 45.056 ;
			RECT	21.173 44.992 21.205 45.056 ;
			RECT	21.509 44.992 21.541 45.056 ;
			RECT	21.845 44.992 21.877 45.056 ;
			RECT	22.181 44.992 22.213 45.056 ;
			RECT	22.517 44.992 22.549 45.056 ;
			RECT	22.853 44.992 22.885 45.056 ;
			RECT	23.189 44.992 23.221 45.056 ;
			RECT	23.525 44.992 23.557 45.056 ;
			RECT	23.861 44.992 23.893 45.056 ;
			RECT	24.197 44.992 24.229 45.056 ;
			RECT	24.533 44.992 24.565 45.056 ;
			RECT	24.869 44.992 24.901 45.056 ;
			RECT	25.205 44.992 25.237 45.056 ;
			RECT	25.541 44.992 25.573 45.056 ;
			RECT	25.877 44.992 25.909 45.056 ;
			RECT	26.213 44.992 26.245 45.056 ;
			RECT	26.549 44.992 26.581 45.056 ;
			RECT	26.885 44.992 26.917 45.056 ;
			RECT	27.221 44.992 27.253 45.056 ;
			RECT	27.557 44.992 27.589 45.056 ;
			RECT	27.878 44.992 27.91 45.056 ;
			RECT	28.214 44.992 28.246 45.056 ;
			RECT	28.55 44.992 28.582 45.056 ;
			RECT	28.886 44.992 28.918 45.056 ;
			RECT	29.222 44.992 29.254 45.056 ;
			RECT	29.558 44.992 29.59 45.056 ;
			RECT	29.894 44.992 29.926 45.056 ;
			RECT	30.23 44.992 30.262 45.056 ;
			RECT	30.566 44.992 30.598 45.056 ;
			RECT	30.902 44.992 30.934 45.056 ;
			RECT	31.238 44.992 31.27 45.056 ;
			RECT	31.574 44.992 31.606 45.056 ;
			RECT	31.91 44.992 31.942 45.056 ;
			RECT	32.246 44.992 32.278 45.056 ;
			RECT	32.582 44.992 32.614 45.056 ;
			RECT	33.254 44.992 33.286 45.056 ;
			RECT	33.59 44.992 33.622 45.056 ;
			RECT	33.926 44.992 33.958 45.056 ;
			RECT	34.262 44.992 34.294 45.056 ;
			RECT	34.598 44.992 34.63 45.056 ;
			RECT	34.934 44.992 34.966 45.056 ;
			RECT	35.27 44.992 35.302 45.056 ;
			RECT	35.606 44.992 35.638 45.056 ;
			RECT	35.942 44.992 35.974 45.056 ;
			RECT	36.278 44.992 36.31 45.056 ;
			RECT	36.614 44.992 36.646 45.056 ;
			RECT	36.95 44.992 36.982 45.056 ;
			RECT	37.286 44.992 37.318 45.056 ;
			RECT	37.622 44.992 37.654 45.056 ;
			RECT	37.958 44.992 37.99 45.056 ;
			RECT	38.294 44.992 38.326 45.056 ;
			RECT	38.63 44.992 38.662 45.056 ;
			RECT	38.966 44.992 38.998 45.056 ;
			RECT	39.302 44.992 39.334 45.056 ;
			RECT	39.638 44.992 39.67 45.056 ;
			RECT	39.974 44.992 40.006 45.056 ;
			RECT	40.31 44.992 40.342 45.056 ;
			RECT	40.646 44.992 40.678 45.056 ;
			RECT	40.982 44.992 41.014 45.056 ;
			RECT	41.318 44.992 41.35 45.056 ;
			RECT	41.654 44.992 41.686 45.056 ;
			RECT	41.99 44.992 42.022 45.056 ;
			RECT	42.326 44.992 42.358 45.056 ;
			RECT	42.662 44.992 42.694 45.056 ;
			RECT	42.998 44.992 43.03 45.056 ;
			RECT	43.334 44.992 43.366 45.056 ;
			RECT	43.67 44.992 43.702 45.056 ;
			RECT	44.342 44.992 44.374 45.056 ;
			RECT	44.678 44.992 44.71 45.056 ;
			RECT	45.014 44.992 45.046 45.056 ;
			RECT	45.35 44.992 45.382 45.056 ;
			RECT	46.022 44.992 46.054 45.056 ;
			RECT	46.358 44.992 46.39 45.056 ;
			RECT	47.03 44.992 47.062 45.056 ;
			RECT	47.366 44.992 47.398 45.056 ;
			RECT	47.702 44.992 47.734 45.056 ;
			RECT	48.038 44.992 48.07 45.056 ;
			RECT	48.374 44.992 48.406 45.056 ;
			RECT	48.71 44.992 48.742 45.056 ;
			RECT	49.046 44.992 49.078 45.056 ;
			RECT	49.311 45.008 49.375 45.04 ;
			RECT	49.566 44.992 49.598 45.056 ;
			RECT	51.92 44.992 51.952 45.056 ;
			RECT	53.91 44.992 53.942 45.056 ;
			RECT	54.251 44.992 54.283 45.056 ;
			RECT	54.657 44.994 54.689 45.058 ;
			RECT	54.812 44.994 54.844 45.058 ;
			RECT	55.224 44.992 55.256 45.056 ;
			RECT	55.706 44.993 55.738 45.057 ;
			RECT	55.842 44.992 55.874 45.056 ;
			RECT	55.985 44.992 56.017 45.056 ;
			RECT	58.606 44.992 58.638 45.056 ;
			RECT	58.829 45.008 58.893 45.04 ;
			RECT	59.126 44.992 59.158 45.056 ;
			RECT	59.462 44.992 59.494 45.056 ;
			RECT	59.798 44.992 59.83 45.056 ;
			RECT	60.134 44.992 60.166 45.056 ;
			RECT	60.47 44.992 60.502 45.056 ;
			RECT	60.806 44.992 60.838 45.056 ;
			RECT	61.142 44.992 61.174 45.056 ;
			RECT	61.814 44.992 61.846 45.056 ;
			RECT	62.15 44.992 62.182 45.056 ;
			RECT	62.822 44.992 62.854 45.056 ;
			RECT	63.158 44.992 63.19 45.056 ;
			RECT	63.494 44.992 63.526 45.056 ;
			RECT	63.83 44.992 63.862 45.056 ;
			RECT	64.502 44.992 64.534 45.056 ;
			RECT	64.838 44.992 64.87 45.056 ;
			RECT	65.174 44.992 65.206 45.056 ;
			RECT	65.51 44.992 65.542 45.056 ;
			RECT	65.846 44.992 65.878 45.056 ;
			RECT	66.182 44.992 66.214 45.056 ;
			RECT	66.518 44.992 66.55 45.056 ;
			RECT	66.854 44.992 66.886 45.056 ;
			RECT	67.19 44.992 67.222 45.056 ;
			RECT	67.526 44.992 67.558 45.056 ;
			RECT	67.862 44.992 67.894 45.056 ;
			RECT	68.198 44.992 68.23 45.056 ;
			RECT	68.534 44.992 68.566 45.056 ;
			RECT	68.87 44.992 68.902 45.056 ;
			RECT	69.206 44.992 69.238 45.056 ;
			RECT	69.542 44.992 69.574 45.056 ;
			RECT	69.878 44.992 69.91 45.056 ;
			RECT	70.214 44.992 70.246 45.056 ;
			RECT	70.55 44.992 70.582 45.056 ;
			RECT	70.886 44.992 70.918 45.056 ;
			RECT	71.222 44.992 71.254 45.056 ;
			RECT	71.558 44.992 71.59 45.056 ;
			RECT	71.894 44.992 71.926 45.056 ;
			RECT	72.23 44.992 72.262 45.056 ;
			RECT	72.566 44.992 72.598 45.056 ;
			RECT	72.902 44.992 72.934 45.056 ;
			RECT	73.238 44.992 73.27 45.056 ;
			RECT	73.574 44.992 73.606 45.056 ;
			RECT	73.91 44.992 73.942 45.056 ;
			RECT	74.246 44.992 74.278 45.056 ;
			RECT	74.582 44.992 74.614 45.056 ;
			RECT	74.918 44.992 74.95 45.056 ;
			RECT	75.59 44.992 75.622 45.056 ;
			RECT	75.926 44.992 75.958 45.056 ;
			RECT	76.262 44.992 76.294 45.056 ;
			RECT	76.598 44.992 76.63 45.056 ;
			RECT	76.934 44.992 76.966 45.056 ;
			RECT	77.27 44.992 77.302 45.056 ;
			RECT	77.606 44.992 77.638 45.056 ;
			RECT	77.942 44.992 77.974 45.056 ;
			RECT	78.278 44.992 78.31 45.056 ;
			RECT	78.614 44.992 78.646 45.056 ;
			RECT	78.95 44.992 78.982 45.056 ;
			RECT	79.286 44.992 79.318 45.056 ;
			RECT	79.622 44.992 79.654 45.056 ;
			RECT	79.958 44.992 79.99 45.056 ;
			RECT	80.294 44.992 80.326 45.056 ;
			RECT	80.615 44.992 80.647 45.056 ;
			RECT	80.951 44.992 80.983 45.056 ;
			RECT	81.287 44.992 81.319 45.056 ;
			RECT	81.623 44.992 81.655 45.056 ;
			RECT	81.959 44.992 81.991 45.056 ;
			RECT	82.295 44.992 82.327 45.056 ;
			RECT	82.631 44.992 82.663 45.056 ;
			RECT	82.967 44.992 82.999 45.056 ;
			RECT	83.303 44.992 83.335 45.056 ;
			RECT	83.639 44.992 83.671 45.056 ;
			RECT	83.975 44.992 84.007 45.056 ;
			RECT	84.311 44.992 84.343 45.056 ;
			RECT	84.647 44.992 84.679 45.056 ;
			RECT	84.983 44.992 85.015 45.056 ;
			RECT	85.319 44.992 85.351 45.056 ;
			RECT	85.655 44.992 85.687 45.056 ;
			RECT	85.991 44.992 86.023 45.056 ;
			RECT	86.327 44.992 86.359 45.056 ;
			RECT	86.663 44.992 86.695 45.056 ;
			RECT	86.999 44.992 87.031 45.056 ;
			RECT	87.335 44.992 87.367 45.056 ;
			RECT	87.671 44.992 87.703 45.056 ;
			RECT	88.007 44.992 88.039 45.056 ;
			RECT	88.343 44.992 88.375 45.056 ;
			RECT	88.679 44.992 88.711 45.056 ;
			RECT	89.015 44.992 89.047 45.056 ;
			RECT	89.351 44.992 89.383 45.056 ;
			RECT	89.687 44.992 89.719 45.056 ;
			RECT	90.023 44.992 90.055 45.056 ;
			RECT	90.359 44.992 90.391 45.056 ;
			RECT	90.695 44.992 90.727 45.056 ;
			RECT	91.031 44.992 91.063 45.056 ;
			RECT	91.367 44.992 91.399 45.056 ;
			RECT	91.703 44.992 91.735 45.056 ;
			RECT	92.039 44.992 92.071 45.056 ;
			RECT	92.375 44.992 92.407 45.056 ;
			RECT	92.711 44.992 92.743 45.056 ;
			RECT	93.047 44.992 93.079 45.056 ;
			RECT	93.383 44.992 93.415 45.056 ;
			RECT	93.719 44.992 93.751 45.056 ;
			RECT	94.055 44.992 94.087 45.056 ;
			RECT	94.391 44.992 94.423 45.056 ;
			RECT	94.727 44.992 94.759 45.056 ;
			RECT	95.063 44.992 95.095 45.056 ;
			RECT	95.399 44.992 95.431 45.056 ;
			RECT	95.735 44.992 95.767 45.056 ;
			RECT	96.071 44.992 96.103 45.056 ;
			RECT	96.407 44.992 96.439 45.056 ;
			RECT	96.743 44.992 96.775 45.056 ;
			RECT	97.079 44.992 97.111 45.056 ;
			RECT	97.415 44.992 97.447 45.056 ;
			RECT	97.751 44.992 97.783 45.056 ;
			RECT	98.087 44.992 98.119 45.056 ;
			RECT	98.423 44.992 98.455 45.056 ;
			RECT	98.759 44.992 98.791 45.056 ;
			RECT	99.095 44.992 99.127 45.056 ;
			RECT	99.431 44.992 99.463 45.056 ;
			RECT	99.767 44.992 99.799 45.056 ;
			RECT	100.103 44.992 100.135 45.056 ;
			RECT	100.439 44.992 100.471 45.056 ;
			RECT	100.775 44.992 100.807 45.056 ;
			RECT	101.111 44.992 101.143 45.056 ;
			RECT	101.447 44.992 101.479 45.056 ;
			RECT	101.783 44.992 101.815 45.056 ;
			RECT	102.379 44.992 102.411 45.056 ;
			RECT	102.605 44.992 102.637 45.056 ;
			RECT	103.565 44.992 103.597 45.056 ;
			RECT	103.791 44.992 103.823 45.056 ;
			RECT	104.387 44.992 104.419 45.056 ;
			RECT	104.723 44.992 104.755 45.056 ;
			RECT	105.059 44.992 105.091 45.056 ;
			RECT	105.395 44.992 105.427 45.056 ;
			RECT	105.731 44.992 105.763 45.056 ;
			RECT	106.067 44.992 106.099 45.056 ;
			RECT	106.403 44.992 106.435 45.056 ;
			RECT	106.739 44.992 106.771 45.056 ;
			RECT	107.075 44.992 107.107 45.056 ;
			RECT	107.411 44.992 107.443 45.056 ;
			RECT	107.747 44.992 107.779 45.056 ;
			RECT	108.083 44.992 108.115 45.056 ;
			RECT	108.419 44.992 108.451 45.056 ;
			RECT	108.755 44.992 108.787 45.056 ;
			RECT	109.091 44.992 109.123 45.056 ;
			RECT	109.427 44.992 109.459 45.056 ;
			RECT	109.763 44.992 109.795 45.056 ;
			RECT	110.099 44.992 110.131 45.056 ;
			RECT	110.435 44.992 110.467 45.056 ;
			RECT	110.771 44.992 110.803 45.056 ;
			RECT	111.107 44.992 111.139 45.056 ;
			RECT	111.443 44.992 111.475 45.056 ;
			RECT	111.779 44.992 111.811 45.056 ;
			RECT	112.115 44.992 112.147 45.056 ;
			RECT	112.451 44.992 112.483 45.056 ;
			RECT	112.787 44.992 112.819 45.056 ;
			RECT	113.123 44.992 113.155 45.056 ;
			RECT	113.459 44.992 113.491 45.056 ;
			RECT	113.795 44.992 113.827 45.056 ;
			RECT	114.131 44.992 114.163 45.056 ;
			RECT	114.467 44.992 114.499 45.056 ;
			RECT	114.803 44.992 114.835 45.056 ;
			RECT	115.139 44.992 115.171 45.056 ;
			RECT	115.475 44.992 115.507 45.056 ;
			RECT	115.811 44.992 115.843 45.056 ;
			RECT	116.147 44.992 116.179 45.056 ;
			RECT	116.483 44.992 116.515 45.056 ;
			RECT	116.819 44.992 116.851 45.056 ;
			RECT	117.155 44.992 117.187 45.056 ;
			RECT	117.491 44.992 117.523 45.056 ;
			RECT	117.827 44.992 117.859 45.056 ;
			RECT	118.163 44.992 118.195 45.056 ;
			RECT	118.499 44.992 118.531 45.056 ;
			RECT	118.835 44.992 118.867 45.056 ;
			RECT	119.171 44.992 119.203 45.056 ;
			RECT	119.507 44.992 119.539 45.056 ;
			RECT	119.843 44.992 119.875 45.056 ;
			RECT	120.179 44.992 120.211 45.056 ;
			RECT	120.515 44.992 120.547 45.056 ;
			RECT	120.851 44.992 120.883 45.056 ;
			RECT	121.187 44.992 121.219 45.056 ;
			RECT	121.523 44.992 121.555 45.056 ;
			RECT	121.859 44.992 121.891 45.056 ;
			RECT	122.195 44.992 122.227 45.056 ;
			RECT	122.531 44.992 122.563 45.056 ;
			RECT	122.867 44.992 122.899 45.056 ;
			RECT	123.203 44.992 123.235 45.056 ;
			RECT	123.539 44.992 123.571 45.056 ;
			RECT	123.875 44.992 123.907 45.056 ;
			RECT	124.211 44.992 124.243 45.056 ;
			RECT	124.547 44.992 124.579 45.056 ;
			RECT	124.883 44.992 124.915 45.056 ;
			RECT	125.219 44.992 125.251 45.056 ;
			RECT	125.555 44.992 125.587 45.056 ;
			RECT	125.876 44.992 125.908 45.056 ;
			RECT	126.212 44.992 126.244 45.056 ;
			RECT	126.548 44.992 126.58 45.056 ;
			RECT	126.884 44.992 126.916 45.056 ;
			RECT	127.22 44.992 127.252 45.056 ;
			RECT	127.556 44.992 127.588 45.056 ;
			RECT	127.892 44.992 127.924 45.056 ;
			RECT	128.228 44.992 128.26 45.056 ;
			RECT	128.564 44.992 128.596 45.056 ;
			RECT	128.9 44.992 128.932 45.056 ;
			RECT	129.236 44.992 129.268 45.056 ;
			RECT	129.572 44.992 129.604 45.056 ;
			RECT	129.908 44.992 129.94 45.056 ;
			RECT	130.244 44.992 130.276 45.056 ;
			RECT	130.58 44.992 130.612 45.056 ;
			RECT	131.252 44.992 131.284 45.056 ;
			RECT	131.588 44.992 131.62 45.056 ;
			RECT	131.924 44.992 131.956 45.056 ;
			RECT	132.26 44.992 132.292 45.056 ;
			RECT	132.596 44.992 132.628 45.056 ;
			RECT	132.932 44.992 132.964 45.056 ;
			RECT	133.268 44.992 133.3 45.056 ;
			RECT	133.604 44.992 133.636 45.056 ;
			RECT	133.94 44.992 133.972 45.056 ;
			RECT	134.276 44.992 134.308 45.056 ;
			RECT	134.612 44.992 134.644 45.056 ;
			RECT	134.948 44.992 134.98 45.056 ;
			RECT	135.284 44.992 135.316 45.056 ;
			RECT	135.62 44.992 135.652 45.056 ;
			RECT	135.956 44.992 135.988 45.056 ;
			RECT	136.292 44.992 136.324 45.056 ;
			RECT	136.628 44.992 136.66 45.056 ;
			RECT	136.964 44.992 136.996 45.056 ;
			RECT	137.3 44.992 137.332 45.056 ;
			RECT	137.636 44.992 137.668 45.056 ;
			RECT	137.972 44.992 138.004 45.056 ;
			RECT	138.308 44.992 138.34 45.056 ;
			RECT	138.644 44.992 138.676 45.056 ;
			RECT	138.98 44.992 139.012 45.056 ;
			RECT	139.316 44.992 139.348 45.056 ;
			RECT	139.652 44.992 139.684 45.056 ;
			RECT	139.988 44.992 140.02 45.056 ;
			RECT	140.324 44.992 140.356 45.056 ;
			RECT	140.66 44.992 140.692 45.056 ;
			RECT	140.996 44.992 141.028 45.056 ;
			RECT	141.332 44.992 141.364 45.056 ;
			RECT	141.668 44.992 141.7 45.056 ;
			RECT	142.34 44.992 142.372 45.056 ;
			RECT	142.676 44.992 142.708 45.056 ;
			RECT	143.012 44.992 143.044 45.056 ;
			RECT	143.348 44.992 143.38 45.056 ;
			RECT	144.02 44.992 144.052 45.056 ;
			RECT	144.356 44.992 144.388 45.056 ;
			RECT	145.028 44.992 145.06 45.056 ;
			RECT	145.364 44.992 145.396 45.056 ;
			RECT	145.7 44.992 145.732 45.056 ;
			RECT	146.036 44.992 146.068 45.056 ;
			RECT	146.372 44.992 146.404 45.056 ;
			RECT	146.708 44.992 146.74 45.056 ;
			RECT	147.044 44.992 147.076 45.056 ;
			RECT	147.309 45.008 147.373 45.04 ;
			RECT	147.564 44.992 147.596 45.056 ;
			RECT	149.918 44.992 149.95 45.056 ;
			RECT	151.908 44.992 151.94 45.056 ;
			RECT	152.249 44.992 152.281 45.056 ;
			RECT	152.655 44.994 152.687 45.058 ;
			RECT	152.81 44.994 152.842 45.058 ;
			RECT	153.222 44.992 153.254 45.056 ;
			RECT	153.704 44.993 153.736 45.057 ;
			RECT	153.84 44.992 153.872 45.056 ;
			RECT	153.983 44.992 154.015 45.056 ;
			RECT	156.604 44.992 156.636 45.056 ;
			RECT	156.827 45.008 156.891 45.04 ;
			RECT	157.124 44.992 157.156 45.056 ;
			RECT	157.46 44.992 157.492 45.056 ;
			RECT	157.796 44.992 157.828 45.056 ;
			RECT	158.132 44.992 158.164 45.056 ;
			RECT	158.468 44.992 158.5 45.056 ;
			RECT	158.804 44.992 158.836 45.056 ;
			RECT	159.14 44.992 159.172 45.056 ;
			RECT	159.812 44.992 159.844 45.056 ;
			RECT	160.148 44.992 160.18 45.056 ;
			RECT	160.82 44.992 160.852 45.056 ;
			RECT	161.156 44.992 161.188 45.056 ;
			RECT	161.492 44.992 161.524 45.056 ;
			RECT	161.828 44.992 161.86 45.056 ;
			RECT	162.5 44.992 162.532 45.056 ;
			RECT	162.836 44.992 162.868 45.056 ;
			RECT	163.172 44.992 163.204 45.056 ;
			RECT	163.508 44.992 163.54 45.056 ;
			RECT	163.844 44.992 163.876 45.056 ;
			RECT	164.18 44.992 164.212 45.056 ;
			RECT	164.516 44.992 164.548 45.056 ;
			RECT	164.852 44.992 164.884 45.056 ;
			RECT	165.188 44.992 165.22 45.056 ;
			RECT	165.524 44.992 165.556 45.056 ;
			RECT	165.86 44.992 165.892 45.056 ;
			RECT	166.196 44.992 166.228 45.056 ;
			RECT	166.532 44.992 166.564 45.056 ;
			RECT	166.868 44.992 166.9 45.056 ;
			RECT	167.204 44.992 167.236 45.056 ;
			RECT	167.54 44.992 167.572 45.056 ;
			RECT	167.876 44.992 167.908 45.056 ;
			RECT	168.212 44.992 168.244 45.056 ;
			RECT	168.548 44.992 168.58 45.056 ;
			RECT	168.884 44.992 168.916 45.056 ;
			RECT	169.22 44.992 169.252 45.056 ;
			RECT	169.556 44.992 169.588 45.056 ;
			RECT	169.892 44.992 169.924 45.056 ;
			RECT	170.228 44.992 170.26 45.056 ;
			RECT	170.564 44.992 170.596 45.056 ;
			RECT	170.9 44.992 170.932 45.056 ;
			RECT	171.236 44.992 171.268 45.056 ;
			RECT	171.572 44.992 171.604 45.056 ;
			RECT	171.908 44.992 171.94 45.056 ;
			RECT	172.244 44.992 172.276 45.056 ;
			RECT	172.58 44.992 172.612 45.056 ;
			RECT	172.916 44.992 172.948 45.056 ;
			RECT	173.588 44.992 173.62 45.056 ;
			RECT	173.924 44.992 173.956 45.056 ;
			RECT	174.26 44.992 174.292 45.056 ;
			RECT	174.596 44.992 174.628 45.056 ;
			RECT	174.932 44.992 174.964 45.056 ;
			RECT	175.268 44.992 175.3 45.056 ;
			RECT	175.604 44.992 175.636 45.056 ;
			RECT	175.94 44.992 175.972 45.056 ;
			RECT	176.276 44.992 176.308 45.056 ;
			RECT	176.612 44.992 176.644 45.056 ;
			RECT	176.948 44.992 176.98 45.056 ;
			RECT	177.284 44.992 177.316 45.056 ;
			RECT	177.62 44.992 177.652 45.056 ;
			RECT	177.956 44.992 177.988 45.056 ;
			RECT	178.292 44.992 178.324 45.056 ;
			RECT	178.613 44.992 178.645 45.056 ;
			RECT	178.949 44.992 178.981 45.056 ;
			RECT	179.285 44.992 179.317 45.056 ;
			RECT	179.621 44.992 179.653 45.056 ;
			RECT	179.957 44.992 179.989 45.056 ;
			RECT	180.293 44.992 180.325 45.056 ;
			RECT	180.629 44.992 180.661 45.056 ;
			RECT	180.965 44.992 180.997 45.056 ;
			RECT	181.301 44.992 181.333 45.056 ;
			RECT	181.637 44.992 181.669 45.056 ;
			RECT	181.973 44.992 182.005 45.056 ;
			RECT	182.309 44.992 182.341 45.056 ;
			RECT	182.645 44.992 182.677 45.056 ;
			RECT	182.981 44.992 183.013 45.056 ;
			RECT	183.317 44.992 183.349 45.056 ;
			RECT	183.653 44.992 183.685 45.056 ;
			RECT	183.989 44.992 184.021 45.056 ;
			RECT	184.325 44.992 184.357 45.056 ;
			RECT	184.661 44.992 184.693 45.056 ;
			RECT	184.997 44.992 185.029 45.056 ;
			RECT	185.333 44.992 185.365 45.056 ;
			RECT	185.669 44.992 185.701 45.056 ;
			RECT	186.005 44.992 186.037 45.056 ;
			RECT	186.341 44.992 186.373 45.056 ;
			RECT	186.677 44.992 186.709 45.056 ;
			RECT	187.013 44.992 187.045 45.056 ;
			RECT	187.349 44.992 187.381 45.056 ;
			RECT	187.685 44.992 187.717 45.056 ;
			RECT	188.021 44.992 188.053 45.056 ;
			RECT	188.357 44.992 188.389 45.056 ;
			RECT	188.693 44.992 188.725 45.056 ;
			RECT	189.029 44.992 189.061 45.056 ;
			RECT	189.365 44.992 189.397 45.056 ;
			RECT	189.701 44.992 189.733 45.056 ;
			RECT	190.037 44.992 190.069 45.056 ;
			RECT	190.373 44.992 190.405 45.056 ;
			RECT	190.709 44.992 190.741 45.056 ;
			RECT	191.045 44.992 191.077 45.056 ;
			RECT	191.381 44.992 191.413 45.056 ;
			RECT	191.717 44.992 191.749 45.056 ;
			RECT	192.053 44.992 192.085 45.056 ;
			RECT	192.389 44.992 192.421 45.056 ;
			RECT	192.725 44.992 192.757 45.056 ;
			RECT	193.061 44.992 193.093 45.056 ;
			RECT	193.397 44.992 193.429 45.056 ;
			RECT	193.733 44.992 193.765 45.056 ;
			RECT	194.069 44.992 194.101 45.056 ;
			RECT	194.405 44.992 194.437 45.056 ;
			RECT	194.741 44.992 194.773 45.056 ;
			RECT	195.077 44.992 195.109 45.056 ;
			RECT	195.413 44.992 195.445 45.056 ;
			RECT	195.749 44.992 195.781 45.056 ;
			RECT	196.085 44.992 196.117 45.056 ;
			RECT	196.421 44.992 196.453 45.056 ;
			RECT	196.757 44.992 196.789 45.056 ;
			RECT	197.093 44.992 197.125 45.056 ;
			RECT	197.429 44.992 197.461 45.056 ;
			RECT	197.765 44.992 197.797 45.056 ;
			RECT	198.101 44.992 198.133 45.056 ;
			RECT	198.437 44.992 198.469 45.056 ;
			RECT	198.773 44.992 198.805 45.056 ;
			RECT	199.109 44.992 199.141 45.056 ;
			RECT	199.445 44.992 199.477 45.056 ;
			RECT	199.781 44.992 199.813 45.056 ;
			RECT	200.377 44.992 200.409 45.056 ;
			RECT	200.603 44.992 200.635 45.056 ;
			RECT	200.9 44.992 200.932 45.056 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 45.843 201.665 45.963 ;
			LAYER	J3 ;
			RECT	1.661 45.871 1.693 45.935 ;
			RECT	2.323 45.871 2.387 45.935 ;
			RECT	3.451 45.871 3.483 45.935 ;
			RECT	4.568 45.887 4.632 45.919 ;
			RECT	4.805 45.871 4.837 45.935 ;
			RECT	5.252 45.871 5.284 45.935 ;
			RECT	5.793 45.887 5.825 45.919 ;
			RECT	49.311 45.871 49.375 45.935 ;
			RECT	49.566 45.871 49.598 45.935 ;
			RECT	51.92 45.871 51.952 45.935 ;
			RECT	52.968 45.871 53.032 45.935 ;
			RECT	53.91 45.871 53.942 45.935 ;
			RECT	54.251 45.871 54.283 45.935 ;
			RECT	54.812 45.871 54.844 45.935 ;
			RECT	55.706 45.871 55.738 45.935 ;
			RECT	55.842 45.871 55.874 45.935 ;
			RECT	55.985 45.871 56.017 45.935 ;
			RECT	57.372 45.871 57.404 45.935 ;
			RECT	58.606 45.871 58.638 45.935 ;
			RECT	58.829 45.871 58.893 45.935 ;
			RECT	102.379 45.887 102.411 45.919 ;
			RECT	103.791 45.887 103.823 45.919 ;
			RECT	147.309 45.871 147.373 45.935 ;
			RECT	147.564 45.871 147.596 45.935 ;
			RECT	149.918 45.871 149.95 45.935 ;
			RECT	150.966 45.871 151.03 45.935 ;
			RECT	151.908 45.871 151.94 45.935 ;
			RECT	152.249 45.871 152.281 45.935 ;
			RECT	152.81 45.871 152.842 45.935 ;
			RECT	153.704 45.871 153.736 45.935 ;
			RECT	153.84 45.871 153.872 45.935 ;
			RECT	153.983 45.871 154.015 45.935 ;
			RECT	155.37 45.871 155.402 45.935 ;
			RECT	156.604 45.871 156.636 45.935 ;
			RECT	156.827 45.871 156.891 45.935 ;
			RECT	200.377 45.887 200.409 45.919 ;
			RECT	200.9 45.871 200.932 45.935 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 46.743 201.665 46.833 ;
			LAYER	J3 ;
			RECT	1.661 46.756 1.693 46.82 ;
			RECT	2.323 46.772 2.387 46.804 ;
			RECT	3.451 46.756 3.483 46.82 ;
			RECT	4.354 46.756 4.386 46.82 ;
			RECT	4.568 46.772 4.632 46.804 ;
			RECT	4.805 46.756 4.837 46.82 ;
			RECT	5.252 46.756 5.284 46.82 ;
			RECT	5.793 46.756 5.825 46.82 ;
			RECT	49.311 46.772 49.375 46.804 ;
			RECT	49.566 46.756 49.598 46.82 ;
			RECT	51.92 46.756 51.952 46.82 ;
			RECT	52.968 46.772 53.032 46.804 ;
			RECT	53.219 46.756 53.251 46.82 ;
			RECT	53.91 46.756 53.942 46.82 ;
			RECT	54.251 46.756 54.283 46.82 ;
			RECT	54.812 46.772 54.844 46.804 ;
			RECT	55.706 46.756 55.738 46.82 ;
			RECT	55.842 46.756 55.874 46.82 ;
			RECT	55.985 46.756 56.017 46.82 ;
			RECT	57.372 46.756 57.404 46.82 ;
			RECT	58.606 46.756 58.638 46.82 ;
			RECT	58.829 46.772 58.893 46.804 ;
			RECT	102.379 46.756 102.411 46.82 ;
			RECT	103.791 46.756 103.823 46.82 ;
			RECT	147.309 46.772 147.373 46.804 ;
			RECT	147.564 46.756 147.596 46.82 ;
			RECT	149.918 46.756 149.95 46.82 ;
			RECT	150.966 46.772 151.03 46.804 ;
			RECT	151.217 46.756 151.249 46.82 ;
			RECT	151.908 46.756 151.94 46.82 ;
			RECT	152.249 46.756 152.281 46.82 ;
			RECT	152.81 46.772 152.842 46.804 ;
			RECT	153.704 46.756 153.736 46.82 ;
			RECT	153.84 46.756 153.872 46.82 ;
			RECT	153.983 46.756 154.015 46.82 ;
			RECT	155.37 46.756 155.402 46.82 ;
			RECT	156.604 46.756 156.636 46.82 ;
			RECT	156.827 46.772 156.891 46.804 ;
			RECT	200.377 46.756 200.409 46.82 ;
			RECT	200.9 46.756 200.932 46.82 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 47.593 201.665 47.713 ;
			LAYER	J3 ;
			RECT	1.645 47.621 1.709 47.685 ;
			RECT	2.323 47.621 2.387 47.685 ;
			RECT	3.451 47.621 3.483 47.685 ;
			RECT	4.179 47.621 4.211 47.685 ;
			RECT	4.568 47.637 4.632 47.669 ;
			RECT	4.805 47.621 4.837 47.685 ;
			RECT	4.96 47.621 4.992 47.685 ;
			RECT	5.252 47.621 5.284 47.685 ;
			RECT	5.808 47.621 5.84 47.685 ;
			RECT	6.179 47.621 6.211 47.685 ;
			RECT	6.347 47.621 6.379 47.685 ;
			RECT	6.515 47.621 6.547 47.685 ;
			RECT	6.683 47.621 6.715 47.685 ;
			RECT	6.851 47.621 6.883 47.685 ;
			RECT	7.019 47.621 7.051 47.685 ;
			RECT	7.187 47.621 7.219 47.685 ;
			RECT	7.355 47.621 7.387 47.685 ;
			RECT	7.523 47.621 7.555 47.685 ;
			RECT	7.691 47.621 7.723 47.685 ;
			RECT	7.859 47.621 7.891 47.685 ;
			RECT	8.027 47.621 8.059 47.685 ;
			RECT	8.195 47.621 8.227 47.685 ;
			RECT	8.363 47.621 8.395 47.685 ;
			RECT	8.531 47.621 8.563 47.685 ;
			RECT	8.699 47.621 8.731 47.685 ;
			RECT	8.867 47.621 8.899 47.685 ;
			RECT	9.035 47.621 9.067 47.685 ;
			RECT	9.203 47.621 9.235 47.685 ;
			RECT	9.371 47.621 9.403 47.685 ;
			RECT	9.539 47.621 9.571 47.685 ;
			RECT	9.707 47.621 9.739 47.685 ;
			RECT	9.875 47.621 9.907 47.685 ;
			RECT	10.043 47.621 10.075 47.685 ;
			RECT	10.211 47.621 10.243 47.685 ;
			RECT	10.379 47.621 10.411 47.685 ;
			RECT	10.547 47.621 10.579 47.685 ;
			RECT	10.715 47.621 10.747 47.685 ;
			RECT	10.883 47.621 10.915 47.685 ;
			RECT	11.051 47.621 11.083 47.685 ;
			RECT	11.219 47.621 11.251 47.685 ;
			RECT	11.387 47.621 11.419 47.685 ;
			RECT	11.555 47.621 11.587 47.685 ;
			RECT	11.723 47.621 11.755 47.685 ;
			RECT	11.891 47.621 11.923 47.685 ;
			RECT	12.059 47.621 12.091 47.685 ;
			RECT	12.227 47.621 12.259 47.685 ;
			RECT	12.395 47.621 12.427 47.685 ;
			RECT	12.563 47.621 12.595 47.685 ;
			RECT	12.731 47.621 12.763 47.685 ;
			RECT	12.899 47.621 12.931 47.685 ;
			RECT	13.067 47.621 13.099 47.685 ;
			RECT	13.235 47.621 13.267 47.685 ;
			RECT	13.403 47.621 13.435 47.685 ;
			RECT	13.571 47.621 13.603 47.685 ;
			RECT	13.739 47.621 13.771 47.685 ;
			RECT	13.907 47.621 13.939 47.685 ;
			RECT	14.075 47.621 14.107 47.685 ;
			RECT	14.243 47.621 14.275 47.685 ;
			RECT	14.411 47.621 14.443 47.685 ;
			RECT	14.579 47.621 14.611 47.685 ;
			RECT	14.747 47.621 14.779 47.685 ;
			RECT	14.915 47.621 14.947 47.685 ;
			RECT	15.083 47.621 15.115 47.685 ;
			RECT	15.251 47.621 15.283 47.685 ;
			RECT	15.419 47.621 15.451 47.685 ;
			RECT	15.587 47.621 15.619 47.685 ;
			RECT	15.755 47.621 15.787 47.685 ;
			RECT	15.923 47.621 15.955 47.685 ;
			RECT	16.091 47.621 16.123 47.685 ;
			RECT	16.259 47.621 16.291 47.685 ;
			RECT	16.427 47.621 16.459 47.685 ;
			RECT	16.595 47.621 16.627 47.685 ;
			RECT	16.763 47.621 16.795 47.685 ;
			RECT	16.931 47.621 16.963 47.685 ;
			RECT	17.099 47.621 17.131 47.685 ;
			RECT	17.267 47.621 17.299 47.685 ;
			RECT	17.435 47.621 17.467 47.685 ;
			RECT	17.603 47.621 17.635 47.685 ;
			RECT	17.771 47.621 17.803 47.685 ;
			RECT	17.939 47.621 17.971 47.685 ;
			RECT	18.107 47.621 18.139 47.685 ;
			RECT	18.275 47.621 18.307 47.685 ;
			RECT	18.443 47.621 18.475 47.685 ;
			RECT	18.611 47.621 18.643 47.685 ;
			RECT	18.779 47.621 18.811 47.685 ;
			RECT	18.947 47.621 18.979 47.685 ;
			RECT	19.115 47.621 19.147 47.685 ;
			RECT	19.283 47.621 19.315 47.685 ;
			RECT	19.451 47.621 19.483 47.685 ;
			RECT	19.619 47.621 19.651 47.685 ;
			RECT	19.787 47.621 19.819 47.685 ;
			RECT	19.955 47.621 19.987 47.685 ;
			RECT	20.123 47.621 20.155 47.685 ;
			RECT	20.291 47.621 20.323 47.685 ;
			RECT	20.459 47.621 20.491 47.685 ;
			RECT	20.627 47.621 20.659 47.685 ;
			RECT	20.795 47.621 20.827 47.685 ;
			RECT	20.963 47.621 20.995 47.685 ;
			RECT	21.131 47.621 21.163 47.685 ;
			RECT	21.299 47.621 21.331 47.685 ;
			RECT	21.467 47.621 21.499 47.685 ;
			RECT	21.635 47.621 21.667 47.685 ;
			RECT	21.803 47.621 21.835 47.685 ;
			RECT	21.971 47.621 22.003 47.685 ;
			RECT	22.139 47.621 22.171 47.685 ;
			RECT	22.307 47.621 22.339 47.685 ;
			RECT	22.475 47.621 22.507 47.685 ;
			RECT	22.643 47.621 22.675 47.685 ;
			RECT	22.811 47.621 22.843 47.685 ;
			RECT	22.979 47.621 23.011 47.685 ;
			RECT	23.147 47.621 23.179 47.685 ;
			RECT	23.315 47.621 23.347 47.685 ;
			RECT	23.483 47.621 23.515 47.685 ;
			RECT	23.651 47.621 23.683 47.685 ;
			RECT	23.819 47.621 23.851 47.685 ;
			RECT	23.987 47.621 24.019 47.685 ;
			RECT	24.155 47.621 24.187 47.685 ;
			RECT	24.323 47.621 24.355 47.685 ;
			RECT	24.491 47.621 24.523 47.685 ;
			RECT	24.659 47.621 24.691 47.685 ;
			RECT	24.827 47.621 24.859 47.685 ;
			RECT	24.995 47.621 25.027 47.685 ;
			RECT	25.163 47.621 25.195 47.685 ;
			RECT	25.331 47.621 25.363 47.685 ;
			RECT	25.499 47.621 25.531 47.685 ;
			RECT	25.667 47.621 25.699 47.685 ;
			RECT	25.835 47.621 25.867 47.685 ;
			RECT	26.003 47.621 26.035 47.685 ;
			RECT	26.171 47.621 26.203 47.685 ;
			RECT	26.339 47.621 26.371 47.685 ;
			RECT	26.507 47.621 26.539 47.685 ;
			RECT	26.675 47.621 26.707 47.685 ;
			RECT	26.843 47.621 26.875 47.685 ;
			RECT	27.011 47.621 27.043 47.685 ;
			RECT	27.179 47.621 27.211 47.685 ;
			RECT	27.347 47.621 27.379 47.685 ;
			RECT	27.515 47.621 27.547 47.685 ;
			RECT	27.683 47.621 27.715 47.685 ;
			RECT	27.851 47.621 27.883 47.685 ;
			RECT	28.019 47.621 28.051 47.685 ;
			RECT	28.187 47.621 28.219 47.685 ;
			RECT	28.355 47.621 28.387 47.685 ;
			RECT	28.523 47.621 28.555 47.685 ;
			RECT	28.691 47.621 28.723 47.685 ;
			RECT	28.859 47.621 28.891 47.685 ;
			RECT	29.027 47.621 29.059 47.685 ;
			RECT	29.195 47.621 29.227 47.685 ;
			RECT	29.363 47.621 29.395 47.685 ;
			RECT	29.531 47.621 29.563 47.685 ;
			RECT	29.699 47.621 29.731 47.685 ;
			RECT	29.867 47.621 29.899 47.685 ;
			RECT	30.035 47.621 30.067 47.685 ;
			RECT	30.203 47.621 30.235 47.685 ;
			RECT	30.371 47.621 30.403 47.685 ;
			RECT	30.539 47.621 30.571 47.685 ;
			RECT	30.707 47.621 30.739 47.685 ;
			RECT	30.875 47.621 30.907 47.685 ;
			RECT	31.043 47.621 31.075 47.685 ;
			RECT	31.211 47.621 31.243 47.685 ;
			RECT	31.379 47.621 31.411 47.685 ;
			RECT	31.547 47.621 31.579 47.685 ;
			RECT	31.715 47.621 31.747 47.685 ;
			RECT	31.883 47.621 31.915 47.685 ;
			RECT	32.051 47.621 32.083 47.685 ;
			RECT	32.219 47.621 32.251 47.685 ;
			RECT	32.387 47.621 32.419 47.685 ;
			RECT	32.555 47.621 32.587 47.685 ;
			RECT	32.723 47.621 32.755 47.685 ;
			RECT	32.891 47.621 32.923 47.685 ;
			RECT	33.059 47.621 33.091 47.685 ;
			RECT	33.227 47.621 33.259 47.685 ;
			RECT	33.395 47.621 33.427 47.685 ;
			RECT	33.563 47.621 33.595 47.685 ;
			RECT	33.731 47.621 33.763 47.685 ;
			RECT	33.899 47.621 33.931 47.685 ;
			RECT	34.067 47.621 34.099 47.685 ;
			RECT	34.235 47.621 34.267 47.685 ;
			RECT	34.403 47.621 34.435 47.685 ;
			RECT	34.571 47.621 34.603 47.685 ;
			RECT	34.739 47.621 34.771 47.685 ;
			RECT	34.907 47.621 34.939 47.685 ;
			RECT	35.075 47.621 35.107 47.685 ;
			RECT	35.243 47.621 35.275 47.685 ;
			RECT	35.411 47.621 35.443 47.685 ;
			RECT	35.579 47.621 35.611 47.685 ;
			RECT	35.747 47.621 35.779 47.685 ;
			RECT	35.915 47.621 35.947 47.685 ;
			RECT	36.083 47.621 36.115 47.685 ;
			RECT	36.251 47.621 36.283 47.685 ;
			RECT	36.419 47.621 36.451 47.685 ;
			RECT	36.587 47.621 36.619 47.685 ;
			RECT	36.755 47.621 36.787 47.685 ;
			RECT	36.923 47.621 36.955 47.685 ;
			RECT	37.091 47.621 37.123 47.685 ;
			RECT	37.259 47.621 37.291 47.685 ;
			RECT	37.427 47.621 37.459 47.685 ;
			RECT	37.595 47.621 37.627 47.685 ;
			RECT	37.763 47.621 37.795 47.685 ;
			RECT	37.931 47.621 37.963 47.685 ;
			RECT	38.099 47.621 38.131 47.685 ;
			RECT	38.267 47.621 38.299 47.685 ;
			RECT	38.435 47.621 38.467 47.685 ;
			RECT	38.603 47.621 38.635 47.685 ;
			RECT	38.771 47.621 38.803 47.685 ;
			RECT	38.939 47.621 38.971 47.685 ;
			RECT	39.107 47.621 39.139 47.685 ;
			RECT	39.275 47.621 39.307 47.685 ;
			RECT	39.443 47.621 39.475 47.685 ;
			RECT	39.611 47.621 39.643 47.685 ;
			RECT	39.779 47.621 39.811 47.685 ;
			RECT	39.947 47.621 39.979 47.685 ;
			RECT	40.115 47.621 40.147 47.685 ;
			RECT	40.283 47.621 40.315 47.685 ;
			RECT	40.451 47.621 40.483 47.685 ;
			RECT	40.619 47.621 40.651 47.685 ;
			RECT	40.787 47.621 40.819 47.685 ;
			RECT	40.955 47.621 40.987 47.685 ;
			RECT	41.123 47.621 41.155 47.685 ;
			RECT	41.291 47.621 41.323 47.685 ;
			RECT	41.459 47.621 41.491 47.685 ;
			RECT	41.627 47.621 41.659 47.685 ;
			RECT	41.795 47.621 41.827 47.685 ;
			RECT	41.963 47.621 41.995 47.685 ;
			RECT	42.131 47.621 42.163 47.685 ;
			RECT	42.299 47.621 42.331 47.685 ;
			RECT	42.467 47.621 42.499 47.685 ;
			RECT	42.635 47.621 42.667 47.685 ;
			RECT	42.803 47.621 42.835 47.685 ;
			RECT	42.971 47.621 43.003 47.685 ;
			RECT	43.139 47.621 43.171 47.685 ;
			RECT	43.307 47.621 43.339 47.685 ;
			RECT	43.475 47.621 43.507 47.685 ;
			RECT	43.643 47.621 43.675 47.685 ;
			RECT	43.811 47.621 43.843 47.685 ;
			RECT	43.979 47.621 44.011 47.685 ;
			RECT	44.147 47.621 44.179 47.685 ;
			RECT	44.315 47.621 44.347 47.685 ;
			RECT	44.483 47.621 44.515 47.685 ;
			RECT	44.651 47.621 44.683 47.685 ;
			RECT	44.819 47.621 44.851 47.685 ;
			RECT	44.987 47.621 45.019 47.685 ;
			RECT	45.155 47.621 45.187 47.685 ;
			RECT	45.323 47.621 45.355 47.685 ;
			RECT	45.491 47.621 45.523 47.685 ;
			RECT	45.659 47.621 45.691 47.685 ;
			RECT	45.827 47.621 45.859 47.685 ;
			RECT	45.995 47.621 46.027 47.685 ;
			RECT	46.163 47.621 46.195 47.685 ;
			RECT	46.331 47.621 46.363 47.685 ;
			RECT	46.499 47.621 46.531 47.685 ;
			RECT	46.667 47.621 46.699 47.685 ;
			RECT	46.835 47.621 46.867 47.685 ;
			RECT	47.003 47.621 47.035 47.685 ;
			RECT	47.171 47.621 47.203 47.685 ;
			RECT	47.339 47.621 47.371 47.685 ;
			RECT	47.507 47.621 47.539 47.685 ;
			RECT	47.675 47.621 47.707 47.685 ;
			RECT	47.843 47.621 47.875 47.685 ;
			RECT	48.011 47.621 48.043 47.685 ;
			RECT	48.179 47.621 48.211 47.685 ;
			RECT	48.347 47.621 48.379 47.685 ;
			RECT	48.515 47.621 48.547 47.685 ;
			RECT	48.683 47.621 48.715 47.685 ;
			RECT	48.851 47.621 48.883 47.685 ;
			RECT	49.019 47.621 49.051 47.685 ;
			RECT	49.187 47.621 49.219 47.685 ;
			RECT	49.311 47.621 49.375 47.685 ;
			RECT	49.557 47.621 49.589 47.685 ;
			RECT	51.92 47.621 51.952 47.685 ;
			RECT	53.079 47.621 53.111 47.685 ;
			RECT	53.219 47.621 53.251 47.685 ;
			RECT	53.91 47.621 53.942 47.685 ;
			RECT	54.251 47.621 54.283 47.685 ;
			RECT	54.812 47.621 54.844 47.685 ;
			RECT	55.466 47.621 55.498 47.685 ;
			RECT	55.706 47.621 55.738 47.685 ;
			RECT	55.842 47.621 55.874 47.685 ;
			RECT	55.969 47.621 56.033 47.685 ;
			RECT	57.372 47.621 57.404 47.685 ;
			RECT	58.615 47.621 58.647 47.685 ;
			RECT	58.829 47.621 58.893 47.685 ;
			RECT	58.985 47.621 59.017 47.685 ;
			RECT	59.153 47.621 59.185 47.685 ;
			RECT	59.321 47.621 59.353 47.685 ;
			RECT	59.489 47.621 59.521 47.685 ;
			RECT	59.657 47.621 59.689 47.685 ;
			RECT	59.825 47.621 59.857 47.685 ;
			RECT	59.993 47.621 60.025 47.685 ;
			RECT	60.161 47.621 60.193 47.685 ;
			RECT	60.329 47.621 60.361 47.685 ;
			RECT	60.497 47.621 60.529 47.685 ;
			RECT	60.665 47.621 60.697 47.685 ;
			RECT	60.833 47.621 60.865 47.685 ;
			RECT	61.001 47.621 61.033 47.685 ;
			RECT	61.169 47.621 61.201 47.685 ;
			RECT	61.337 47.621 61.369 47.685 ;
			RECT	61.505 47.621 61.537 47.685 ;
			RECT	61.673 47.621 61.705 47.685 ;
			RECT	61.841 47.621 61.873 47.685 ;
			RECT	62.009 47.621 62.041 47.685 ;
			RECT	62.177 47.621 62.209 47.685 ;
			RECT	62.345 47.621 62.377 47.685 ;
			RECT	62.513 47.621 62.545 47.685 ;
			RECT	62.681 47.621 62.713 47.685 ;
			RECT	62.849 47.621 62.881 47.685 ;
			RECT	63.017 47.621 63.049 47.685 ;
			RECT	63.185 47.621 63.217 47.685 ;
			RECT	63.353 47.621 63.385 47.685 ;
			RECT	63.521 47.621 63.553 47.685 ;
			RECT	63.689 47.621 63.721 47.685 ;
			RECT	63.857 47.621 63.889 47.685 ;
			RECT	64.025 47.621 64.057 47.685 ;
			RECT	64.193 47.621 64.225 47.685 ;
			RECT	64.361 47.621 64.393 47.685 ;
			RECT	64.529 47.621 64.561 47.685 ;
			RECT	64.697 47.621 64.729 47.685 ;
			RECT	64.865 47.621 64.897 47.685 ;
			RECT	65.033 47.621 65.065 47.685 ;
			RECT	65.201 47.621 65.233 47.685 ;
			RECT	65.369 47.621 65.401 47.685 ;
			RECT	65.537 47.621 65.569 47.685 ;
			RECT	65.705 47.621 65.737 47.685 ;
			RECT	65.873 47.621 65.905 47.685 ;
			RECT	66.041 47.621 66.073 47.685 ;
			RECT	66.209 47.621 66.241 47.685 ;
			RECT	66.377 47.621 66.409 47.685 ;
			RECT	66.545 47.621 66.577 47.685 ;
			RECT	66.713 47.621 66.745 47.685 ;
			RECT	66.881 47.621 66.913 47.685 ;
			RECT	67.049 47.621 67.081 47.685 ;
			RECT	67.217 47.621 67.249 47.685 ;
			RECT	67.385 47.621 67.417 47.685 ;
			RECT	67.553 47.621 67.585 47.685 ;
			RECT	67.721 47.621 67.753 47.685 ;
			RECT	67.889 47.621 67.921 47.685 ;
			RECT	68.057 47.621 68.089 47.685 ;
			RECT	68.225 47.621 68.257 47.685 ;
			RECT	68.393 47.621 68.425 47.685 ;
			RECT	68.561 47.621 68.593 47.685 ;
			RECT	68.729 47.621 68.761 47.685 ;
			RECT	68.897 47.621 68.929 47.685 ;
			RECT	69.065 47.621 69.097 47.685 ;
			RECT	69.233 47.621 69.265 47.685 ;
			RECT	69.401 47.621 69.433 47.685 ;
			RECT	69.569 47.621 69.601 47.685 ;
			RECT	69.737 47.621 69.769 47.685 ;
			RECT	69.905 47.621 69.937 47.685 ;
			RECT	70.073 47.621 70.105 47.685 ;
			RECT	70.241 47.621 70.273 47.685 ;
			RECT	70.409 47.621 70.441 47.685 ;
			RECT	70.577 47.621 70.609 47.685 ;
			RECT	70.745 47.621 70.777 47.685 ;
			RECT	70.913 47.621 70.945 47.685 ;
			RECT	71.081 47.621 71.113 47.685 ;
			RECT	71.249 47.621 71.281 47.685 ;
			RECT	71.417 47.621 71.449 47.685 ;
			RECT	71.585 47.621 71.617 47.685 ;
			RECT	71.753 47.621 71.785 47.685 ;
			RECT	71.921 47.621 71.953 47.685 ;
			RECT	72.089 47.621 72.121 47.685 ;
			RECT	72.257 47.621 72.289 47.685 ;
			RECT	72.425 47.621 72.457 47.685 ;
			RECT	72.593 47.621 72.625 47.685 ;
			RECT	72.761 47.621 72.793 47.685 ;
			RECT	72.929 47.621 72.961 47.685 ;
			RECT	73.097 47.621 73.129 47.685 ;
			RECT	73.265 47.621 73.297 47.685 ;
			RECT	73.433 47.621 73.465 47.685 ;
			RECT	73.601 47.621 73.633 47.685 ;
			RECT	73.769 47.621 73.801 47.685 ;
			RECT	73.937 47.621 73.969 47.685 ;
			RECT	74.105 47.621 74.137 47.685 ;
			RECT	74.273 47.621 74.305 47.685 ;
			RECT	74.441 47.621 74.473 47.685 ;
			RECT	74.609 47.621 74.641 47.685 ;
			RECT	74.777 47.621 74.809 47.685 ;
			RECT	74.945 47.621 74.977 47.685 ;
			RECT	75.113 47.621 75.145 47.685 ;
			RECT	75.281 47.621 75.313 47.685 ;
			RECT	75.449 47.621 75.481 47.685 ;
			RECT	75.617 47.621 75.649 47.685 ;
			RECT	75.785 47.621 75.817 47.685 ;
			RECT	75.953 47.621 75.985 47.685 ;
			RECT	76.121 47.621 76.153 47.685 ;
			RECT	76.289 47.621 76.321 47.685 ;
			RECT	76.457 47.621 76.489 47.685 ;
			RECT	76.625 47.621 76.657 47.685 ;
			RECT	76.793 47.621 76.825 47.685 ;
			RECT	76.961 47.621 76.993 47.685 ;
			RECT	77.129 47.621 77.161 47.685 ;
			RECT	77.297 47.621 77.329 47.685 ;
			RECT	77.465 47.621 77.497 47.685 ;
			RECT	77.633 47.621 77.665 47.685 ;
			RECT	77.801 47.621 77.833 47.685 ;
			RECT	77.969 47.621 78.001 47.685 ;
			RECT	78.137 47.621 78.169 47.685 ;
			RECT	78.305 47.621 78.337 47.685 ;
			RECT	78.473 47.621 78.505 47.685 ;
			RECT	78.641 47.621 78.673 47.685 ;
			RECT	78.809 47.621 78.841 47.685 ;
			RECT	78.977 47.621 79.009 47.685 ;
			RECT	79.145 47.621 79.177 47.685 ;
			RECT	79.313 47.621 79.345 47.685 ;
			RECT	79.481 47.621 79.513 47.685 ;
			RECT	79.649 47.621 79.681 47.685 ;
			RECT	79.817 47.621 79.849 47.685 ;
			RECT	79.985 47.621 80.017 47.685 ;
			RECT	80.153 47.621 80.185 47.685 ;
			RECT	80.321 47.621 80.353 47.685 ;
			RECT	80.489 47.621 80.521 47.685 ;
			RECT	80.657 47.621 80.689 47.685 ;
			RECT	80.825 47.621 80.857 47.685 ;
			RECT	80.993 47.621 81.025 47.685 ;
			RECT	81.161 47.621 81.193 47.685 ;
			RECT	81.329 47.621 81.361 47.685 ;
			RECT	81.497 47.621 81.529 47.685 ;
			RECT	81.665 47.621 81.697 47.685 ;
			RECT	81.833 47.621 81.865 47.685 ;
			RECT	82.001 47.621 82.033 47.685 ;
			RECT	82.169 47.621 82.201 47.685 ;
			RECT	82.337 47.621 82.369 47.685 ;
			RECT	82.505 47.621 82.537 47.685 ;
			RECT	82.673 47.621 82.705 47.685 ;
			RECT	82.841 47.621 82.873 47.685 ;
			RECT	83.009 47.621 83.041 47.685 ;
			RECT	83.177 47.621 83.209 47.685 ;
			RECT	83.345 47.621 83.377 47.685 ;
			RECT	83.513 47.621 83.545 47.685 ;
			RECT	83.681 47.621 83.713 47.685 ;
			RECT	83.849 47.621 83.881 47.685 ;
			RECT	84.017 47.621 84.049 47.685 ;
			RECT	84.185 47.621 84.217 47.685 ;
			RECT	84.353 47.621 84.385 47.685 ;
			RECT	84.521 47.621 84.553 47.685 ;
			RECT	84.689 47.621 84.721 47.685 ;
			RECT	84.857 47.621 84.889 47.685 ;
			RECT	85.025 47.621 85.057 47.685 ;
			RECT	85.193 47.621 85.225 47.685 ;
			RECT	85.361 47.621 85.393 47.685 ;
			RECT	85.529 47.621 85.561 47.685 ;
			RECT	85.697 47.621 85.729 47.685 ;
			RECT	85.865 47.621 85.897 47.685 ;
			RECT	86.033 47.621 86.065 47.685 ;
			RECT	86.201 47.621 86.233 47.685 ;
			RECT	86.369 47.621 86.401 47.685 ;
			RECT	86.537 47.621 86.569 47.685 ;
			RECT	86.705 47.621 86.737 47.685 ;
			RECT	86.873 47.621 86.905 47.685 ;
			RECT	87.041 47.621 87.073 47.685 ;
			RECT	87.209 47.621 87.241 47.685 ;
			RECT	87.377 47.621 87.409 47.685 ;
			RECT	87.545 47.621 87.577 47.685 ;
			RECT	87.713 47.621 87.745 47.685 ;
			RECT	87.881 47.621 87.913 47.685 ;
			RECT	88.049 47.621 88.081 47.685 ;
			RECT	88.217 47.621 88.249 47.685 ;
			RECT	88.385 47.621 88.417 47.685 ;
			RECT	88.553 47.621 88.585 47.685 ;
			RECT	88.721 47.621 88.753 47.685 ;
			RECT	88.889 47.621 88.921 47.685 ;
			RECT	89.057 47.621 89.089 47.685 ;
			RECT	89.225 47.621 89.257 47.685 ;
			RECT	89.393 47.621 89.425 47.685 ;
			RECT	89.561 47.621 89.593 47.685 ;
			RECT	89.729 47.621 89.761 47.685 ;
			RECT	89.897 47.621 89.929 47.685 ;
			RECT	90.065 47.621 90.097 47.685 ;
			RECT	90.233 47.621 90.265 47.685 ;
			RECT	90.401 47.621 90.433 47.685 ;
			RECT	90.569 47.621 90.601 47.685 ;
			RECT	90.737 47.621 90.769 47.685 ;
			RECT	90.905 47.621 90.937 47.685 ;
			RECT	91.073 47.621 91.105 47.685 ;
			RECT	91.241 47.621 91.273 47.685 ;
			RECT	91.409 47.621 91.441 47.685 ;
			RECT	91.577 47.621 91.609 47.685 ;
			RECT	91.745 47.621 91.777 47.685 ;
			RECT	91.913 47.621 91.945 47.685 ;
			RECT	92.081 47.621 92.113 47.685 ;
			RECT	92.249 47.621 92.281 47.685 ;
			RECT	92.417 47.621 92.449 47.685 ;
			RECT	92.585 47.621 92.617 47.685 ;
			RECT	92.753 47.621 92.785 47.685 ;
			RECT	92.921 47.621 92.953 47.685 ;
			RECT	93.089 47.621 93.121 47.685 ;
			RECT	93.257 47.621 93.289 47.685 ;
			RECT	93.425 47.621 93.457 47.685 ;
			RECT	93.593 47.621 93.625 47.685 ;
			RECT	93.761 47.621 93.793 47.685 ;
			RECT	93.929 47.621 93.961 47.685 ;
			RECT	94.097 47.621 94.129 47.685 ;
			RECT	94.265 47.621 94.297 47.685 ;
			RECT	94.433 47.621 94.465 47.685 ;
			RECT	94.601 47.621 94.633 47.685 ;
			RECT	94.769 47.621 94.801 47.685 ;
			RECT	94.937 47.621 94.969 47.685 ;
			RECT	95.105 47.621 95.137 47.685 ;
			RECT	95.273 47.621 95.305 47.685 ;
			RECT	95.441 47.621 95.473 47.685 ;
			RECT	95.609 47.621 95.641 47.685 ;
			RECT	95.777 47.621 95.809 47.685 ;
			RECT	95.945 47.621 95.977 47.685 ;
			RECT	96.113 47.621 96.145 47.685 ;
			RECT	96.281 47.621 96.313 47.685 ;
			RECT	96.449 47.621 96.481 47.685 ;
			RECT	96.617 47.621 96.649 47.685 ;
			RECT	96.785 47.621 96.817 47.685 ;
			RECT	96.953 47.621 96.985 47.685 ;
			RECT	97.121 47.621 97.153 47.685 ;
			RECT	97.289 47.621 97.321 47.685 ;
			RECT	97.457 47.621 97.489 47.685 ;
			RECT	97.625 47.621 97.657 47.685 ;
			RECT	97.793 47.621 97.825 47.685 ;
			RECT	97.961 47.621 97.993 47.685 ;
			RECT	98.129 47.621 98.161 47.685 ;
			RECT	98.297 47.621 98.329 47.685 ;
			RECT	98.465 47.621 98.497 47.685 ;
			RECT	98.633 47.621 98.665 47.685 ;
			RECT	98.801 47.621 98.833 47.685 ;
			RECT	98.969 47.621 99.001 47.685 ;
			RECT	99.137 47.621 99.169 47.685 ;
			RECT	99.305 47.621 99.337 47.685 ;
			RECT	99.473 47.621 99.505 47.685 ;
			RECT	99.641 47.621 99.673 47.685 ;
			RECT	99.809 47.621 99.841 47.685 ;
			RECT	99.977 47.621 100.009 47.685 ;
			RECT	100.145 47.621 100.177 47.685 ;
			RECT	100.313 47.621 100.345 47.685 ;
			RECT	100.481 47.621 100.513 47.685 ;
			RECT	100.649 47.621 100.681 47.685 ;
			RECT	100.817 47.621 100.849 47.685 ;
			RECT	100.985 47.621 101.017 47.685 ;
			RECT	101.153 47.621 101.185 47.685 ;
			RECT	101.321 47.621 101.353 47.685 ;
			RECT	101.489 47.621 101.521 47.685 ;
			RECT	101.657 47.621 101.689 47.685 ;
			RECT	101.825 47.621 101.857 47.685 ;
			RECT	101.993 47.621 102.025 47.685 ;
			RECT	102.364 47.621 102.396 47.685 ;
			RECT	103.806 47.621 103.838 47.685 ;
			RECT	104.177 47.621 104.209 47.685 ;
			RECT	104.345 47.621 104.377 47.685 ;
			RECT	104.513 47.621 104.545 47.685 ;
			RECT	104.681 47.621 104.713 47.685 ;
			RECT	104.849 47.621 104.881 47.685 ;
			RECT	105.017 47.621 105.049 47.685 ;
			RECT	105.185 47.621 105.217 47.685 ;
			RECT	105.353 47.621 105.385 47.685 ;
			RECT	105.521 47.621 105.553 47.685 ;
			RECT	105.689 47.621 105.721 47.685 ;
			RECT	105.857 47.621 105.889 47.685 ;
			RECT	106.025 47.621 106.057 47.685 ;
			RECT	106.193 47.621 106.225 47.685 ;
			RECT	106.361 47.621 106.393 47.685 ;
			RECT	106.529 47.621 106.561 47.685 ;
			RECT	106.697 47.621 106.729 47.685 ;
			RECT	106.865 47.621 106.897 47.685 ;
			RECT	107.033 47.621 107.065 47.685 ;
			RECT	107.201 47.621 107.233 47.685 ;
			RECT	107.369 47.621 107.401 47.685 ;
			RECT	107.537 47.621 107.569 47.685 ;
			RECT	107.705 47.621 107.737 47.685 ;
			RECT	107.873 47.621 107.905 47.685 ;
			RECT	108.041 47.621 108.073 47.685 ;
			RECT	108.209 47.621 108.241 47.685 ;
			RECT	108.377 47.621 108.409 47.685 ;
			RECT	108.545 47.621 108.577 47.685 ;
			RECT	108.713 47.621 108.745 47.685 ;
			RECT	108.881 47.621 108.913 47.685 ;
			RECT	109.049 47.621 109.081 47.685 ;
			RECT	109.217 47.621 109.249 47.685 ;
			RECT	109.385 47.621 109.417 47.685 ;
			RECT	109.553 47.621 109.585 47.685 ;
			RECT	109.721 47.621 109.753 47.685 ;
			RECT	109.889 47.621 109.921 47.685 ;
			RECT	110.057 47.621 110.089 47.685 ;
			RECT	110.225 47.621 110.257 47.685 ;
			RECT	110.393 47.621 110.425 47.685 ;
			RECT	110.561 47.621 110.593 47.685 ;
			RECT	110.729 47.621 110.761 47.685 ;
			RECT	110.897 47.621 110.929 47.685 ;
			RECT	111.065 47.621 111.097 47.685 ;
			RECT	111.233 47.621 111.265 47.685 ;
			RECT	111.401 47.621 111.433 47.685 ;
			RECT	111.569 47.621 111.601 47.685 ;
			RECT	111.737 47.621 111.769 47.685 ;
			RECT	111.905 47.621 111.937 47.685 ;
			RECT	112.073 47.621 112.105 47.685 ;
			RECT	112.241 47.621 112.273 47.685 ;
			RECT	112.409 47.621 112.441 47.685 ;
			RECT	112.577 47.621 112.609 47.685 ;
			RECT	112.745 47.621 112.777 47.685 ;
			RECT	112.913 47.621 112.945 47.685 ;
			RECT	113.081 47.621 113.113 47.685 ;
			RECT	113.249 47.621 113.281 47.685 ;
			RECT	113.417 47.621 113.449 47.685 ;
			RECT	113.585 47.621 113.617 47.685 ;
			RECT	113.753 47.621 113.785 47.685 ;
			RECT	113.921 47.621 113.953 47.685 ;
			RECT	114.089 47.621 114.121 47.685 ;
			RECT	114.257 47.621 114.289 47.685 ;
			RECT	114.425 47.621 114.457 47.685 ;
			RECT	114.593 47.621 114.625 47.685 ;
			RECT	114.761 47.621 114.793 47.685 ;
			RECT	114.929 47.621 114.961 47.685 ;
			RECT	115.097 47.621 115.129 47.685 ;
			RECT	115.265 47.621 115.297 47.685 ;
			RECT	115.433 47.621 115.465 47.685 ;
			RECT	115.601 47.621 115.633 47.685 ;
			RECT	115.769 47.621 115.801 47.685 ;
			RECT	115.937 47.621 115.969 47.685 ;
			RECT	116.105 47.621 116.137 47.685 ;
			RECT	116.273 47.621 116.305 47.685 ;
			RECT	116.441 47.621 116.473 47.685 ;
			RECT	116.609 47.621 116.641 47.685 ;
			RECT	116.777 47.621 116.809 47.685 ;
			RECT	116.945 47.621 116.977 47.685 ;
			RECT	117.113 47.621 117.145 47.685 ;
			RECT	117.281 47.621 117.313 47.685 ;
			RECT	117.449 47.621 117.481 47.685 ;
			RECT	117.617 47.621 117.649 47.685 ;
			RECT	117.785 47.621 117.817 47.685 ;
			RECT	117.953 47.621 117.985 47.685 ;
			RECT	118.121 47.621 118.153 47.685 ;
			RECT	118.289 47.621 118.321 47.685 ;
			RECT	118.457 47.621 118.489 47.685 ;
			RECT	118.625 47.621 118.657 47.685 ;
			RECT	118.793 47.621 118.825 47.685 ;
			RECT	118.961 47.621 118.993 47.685 ;
			RECT	119.129 47.621 119.161 47.685 ;
			RECT	119.297 47.621 119.329 47.685 ;
			RECT	119.465 47.621 119.497 47.685 ;
			RECT	119.633 47.621 119.665 47.685 ;
			RECT	119.801 47.621 119.833 47.685 ;
			RECT	119.969 47.621 120.001 47.685 ;
			RECT	120.137 47.621 120.169 47.685 ;
			RECT	120.305 47.621 120.337 47.685 ;
			RECT	120.473 47.621 120.505 47.685 ;
			RECT	120.641 47.621 120.673 47.685 ;
			RECT	120.809 47.621 120.841 47.685 ;
			RECT	120.977 47.621 121.009 47.685 ;
			RECT	121.145 47.621 121.177 47.685 ;
			RECT	121.313 47.621 121.345 47.685 ;
			RECT	121.481 47.621 121.513 47.685 ;
			RECT	121.649 47.621 121.681 47.685 ;
			RECT	121.817 47.621 121.849 47.685 ;
			RECT	121.985 47.621 122.017 47.685 ;
			RECT	122.153 47.621 122.185 47.685 ;
			RECT	122.321 47.621 122.353 47.685 ;
			RECT	122.489 47.621 122.521 47.685 ;
			RECT	122.657 47.621 122.689 47.685 ;
			RECT	122.825 47.621 122.857 47.685 ;
			RECT	122.993 47.621 123.025 47.685 ;
			RECT	123.161 47.621 123.193 47.685 ;
			RECT	123.329 47.621 123.361 47.685 ;
			RECT	123.497 47.621 123.529 47.685 ;
			RECT	123.665 47.621 123.697 47.685 ;
			RECT	123.833 47.621 123.865 47.685 ;
			RECT	124.001 47.621 124.033 47.685 ;
			RECT	124.169 47.621 124.201 47.685 ;
			RECT	124.337 47.621 124.369 47.685 ;
			RECT	124.505 47.621 124.537 47.685 ;
			RECT	124.673 47.621 124.705 47.685 ;
			RECT	124.841 47.621 124.873 47.685 ;
			RECT	125.009 47.621 125.041 47.685 ;
			RECT	125.177 47.621 125.209 47.685 ;
			RECT	125.345 47.621 125.377 47.685 ;
			RECT	125.513 47.621 125.545 47.685 ;
			RECT	125.681 47.621 125.713 47.685 ;
			RECT	125.849 47.621 125.881 47.685 ;
			RECT	126.017 47.621 126.049 47.685 ;
			RECT	126.185 47.621 126.217 47.685 ;
			RECT	126.353 47.621 126.385 47.685 ;
			RECT	126.521 47.621 126.553 47.685 ;
			RECT	126.689 47.621 126.721 47.685 ;
			RECT	126.857 47.621 126.889 47.685 ;
			RECT	127.025 47.621 127.057 47.685 ;
			RECT	127.193 47.621 127.225 47.685 ;
			RECT	127.361 47.621 127.393 47.685 ;
			RECT	127.529 47.621 127.561 47.685 ;
			RECT	127.697 47.621 127.729 47.685 ;
			RECT	127.865 47.621 127.897 47.685 ;
			RECT	128.033 47.621 128.065 47.685 ;
			RECT	128.201 47.621 128.233 47.685 ;
			RECT	128.369 47.621 128.401 47.685 ;
			RECT	128.537 47.621 128.569 47.685 ;
			RECT	128.705 47.621 128.737 47.685 ;
			RECT	128.873 47.621 128.905 47.685 ;
			RECT	129.041 47.621 129.073 47.685 ;
			RECT	129.209 47.621 129.241 47.685 ;
			RECT	129.377 47.621 129.409 47.685 ;
			RECT	129.545 47.621 129.577 47.685 ;
			RECT	129.713 47.621 129.745 47.685 ;
			RECT	129.881 47.621 129.913 47.685 ;
			RECT	130.049 47.621 130.081 47.685 ;
			RECT	130.217 47.621 130.249 47.685 ;
			RECT	130.385 47.621 130.417 47.685 ;
			RECT	130.553 47.621 130.585 47.685 ;
			RECT	130.721 47.621 130.753 47.685 ;
			RECT	130.889 47.621 130.921 47.685 ;
			RECT	131.057 47.621 131.089 47.685 ;
			RECT	131.225 47.621 131.257 47.685 ;
			RECT	131.393 47.621 131.425 47.685 ;
			RECT	131.561 47.621 131.593 47.685 ;
			RECT	131.729 47.621 131.761 47.685 ;
			RECT	131.897 47.621 131.929 47.685 ;
			RECT	132.065 47.621 132.097 47.685 ;
			RECT	132.233 47.621 132.265 47.685 ;
			RECT	132.401 47.621 132.433 47.685 ;
			RECT	132.569 47.621 132.601 47.685 ;
			RECT	132.737 47.621 132.769 47.685 ;
			RECT	132.905 47.621 132.937 47.685 ;
			RECT	133.073 47.621 133.105 47.685 ;
			RECT	133.241 47.621 133.273 47.685 ;
			RECT	133.409 47.621 133.441 47.685 ;
			RECT	133.577 47.621 133.609 47.685 ;
			RECT	133.745 47.621 133.777 47.685 ;
			RECT	133.913 47.621 133.945 47.685 ;
			RECT	134.081 47.621 134.113 47.685 ;
			RECT	134.249 47.621 134.281 47.685 ;
			RECT	134.417 47.621 134.449 47.685 ;
			RECT	134.585 47.621 134.617 47.685 ;
			RECT	134.753 47.621 134.785 47.685 ;
			RECT	134.921 47.621 134.953 47.685 ;
			RECT	135.089 47.621 135.121 47.685 ;
			RECT	135.257 47.621 135.289 47.685 ;
			RECT	135.425 47.621 135.457 47.685 ;
			RECT	135.593 47.621 135.625 47.685 ;
			RECT	135.761 47.621 135.793 47.685 ;
			RECT	135.929 47.621 135.961 47.685 ;
			RECT	136.097 47.621 136.129 47.685 ;
			RECT	136.265 47.621 136.297 47.685 ;
			RECT	136.433 47.621 136.465 47.685 ;
			RECT	136.601 47.621 136.633 47.685 ;
			RECT	136.769 47.621 136.801 47.685 ;
			RECT	136.937 47.621 136.969 47.685 ;
			RECT	137.105 47.621 137.137 47.685 ;
			RECT	137.273 47.621 137.305 47.685 ;
			RECT	137.441 47.621 137.473 47.685 ;
			RECT	137.609 47.621 137.641 47.685 ;
			RECT	137.777 47.621 137.809 47.685 ;
			RECT	137.945 47.621 137.977 47.685 ;
			RECT	138.113 47.621 138.145 47.685 ;
			RECT	138.281 47.621 138.313 47.685 ;
			RECT	138.449 47.621 138.481 47.685 ;
			RECT	138.617 47.621 138.649 47.685 ;
			RECT	138.785 47.621 138.817 47.685 ;
			RECT	138.953 47.621 138.985 47.685 ;
			RECT	139.121 47.621 139.153 47.685 ;
			RECT	139.289 47.621 139.321 47.685 ;
			RECT	139.457 47.621 139.489 47.685 ;
			RECT	139.625 47.621 139.657 47.685 ;
			RECT	139.793 47.621 139.825 47.685 ;
			RECT	139.961 47.621 139.993 47.685 ;
			RECT	140.129 47.621 140.161 47.685 ;
			RECT	140.297 47.621 140.329 47.685 ;
			RECT	140.465 47.621 140.497 47.685 ;
			RECT	140.633 47.621 140.665 47.685 ;
			RECT	140.801 47.621 140.833 47.685 ;
			RECT	140.969 47.621 141.001 47.685 ;
			RECT	141.137 47.621 141.169 47.685 ;
			RECT	141.305 47.621 141.337 47.685 ;
			RECT	141.473 47.621 141.505 47.685 ;
			RECT	141.641 47.621 141.673 47.685 ;
			RECT	141.809 47.621 141.841 47.685 ;
			RECT	141.977 47.621 142.009 47.685 ;
			RECT	142.145 47.621 142.177 47.685 ;
			RECT	142.313 47.621 142.345 47.685 ;
			RECT	142.481 47.621 142.513 47.685 ;
			RECT	142.649 47.621 142.681 47.685 ;
			RECT	142.817 47.621 142.849 47.685 ;
			RECT	142.985 47.621 143.017 47.685 ;
			RECT	143.153 47.621 143.185 47.685 ;
			RECT	143.321 47.621 143.353 47.685 ;
			RECT	143.489 47.621 143.521 47.685 ;
			RECT	143.657 47.621 143.689 47.685 ;
			RECT	143.825 47.621 143.857 47.685 ;
			RECT	143.993 47.621 144.025 47.685 ;
			RECT	144.161 47.621 144.193 47.685 ;
			RECT	144.329 47.621 144.361 47.685 ;
			RECT	144.497 47.621 144.529 47.685 ;
			RECT	144.665 47.621 144.697 47.685 ;
			RECT	144.833 47.621 144.865 47.685 ;
			RECT	145.001 47.621 145.033 47.685 ;
			RECT	145.169 47.621 145.201 47.685 ;
			RECT	145.337 47.621 145.369 47.685 ;
			RECT	145.505 47.621 145.537 47.685 ;
			RECT	145.673 47.621 145.705 47.685 ;
			RECT	145.841 47.621 145.873 47.685 ;
			RECT	146.009 47.621 146.041 47.685 ;
			RECT	146.177 47.621 146.209 47.685 ;
			RECT	146.345 47.621 146.377 47.685 ;
			RECT	146.513 47.621 146.545 47.685 ;
			RECT	146.681 47.621 146.713 47.685 ;
			RECT	146.849 47.621 146.881 47.685 ;
			RECT	147.017 47.621 147.049 47.685 ;
			RECT	147.185 47.621 147.217 47.685 ;
			RECT	147.309 47.621 147.373 47.685 ;
			RECT	147.555 47.621 147.587 47.685 ;
			RECT	149.918 47.621 149.95 47.685 ;
			RECT	151.077 47.621 151.109 47.685 ;
			RECT	151.217 47.621 151.249 47.685 ;
			RECT	151.908 47.621 151.94 47.685 ;
			RECT	152.249 47.621 152.281 47.685 ;
			RECT	152.81 47.621 152.842 47.685 ;
			RECT	153.464 47.621 153.496 47.685 ;
			RECT	153.704 47.621 153.736 47.685 ;
			RECT	153.84 47.621 153.872 47.685 ;
			RECT	153.967 47.621 154.031 47.685 ;
			RECT	155.37 47.621 155.402 47.685 ;
			RECT	156.613 47.621 156.645 47.685 ;
			RECT	156.827 47.621 156.891 47.685 ;
			RECT	156.983 47.621 157.015 47.685 ;
			RECT	157.151 47.621 157.183 47.685 ;
			RECT	157.319 47.621 157.351 47.685 ;
			RECT	157.487 47.621 157.519 47.685 ;
			RECT	157.655 47.621 157.687 47.685 ;
			RECT	157.823 47.621 157.855 47.685 ;
			RECT	157.991 47.621 158.023 47.685 ;
			RECT	158.159 47.621 158.191 47.685 ;
			RECT	158.327 47.621 158.359 47.685 ;
			RECT	158.495 47.621 158.527 47.685 ;
			RECT	158.663 47.621 158.695 47.685 ;
			RECT	158.831 47.621 158.863 47.685 ;
			RECT	158.999 47.621 159.031 47.685 ;
			RECT	159.167 47.621 159.199 47.685 ;
			RECT	159.335 47.621 159.367 47.685 ;
			RECT	159.503 47.621 159.535 47.685 ;
			RECT	159.671 47.621 159.703 47.685 ;
			RECT	159.839 47.621 159.871 47.685 ;
			RECT	160.007 47.621 160.039 47.685 ;
			RECT	160.175 47.621 160.207 47.685 ;
			RECT	160.343 47.621 160.375 47.685 ;
			RECT	160.511 47.621 160.543 47.685 ;
			RECT	160.679 47.621 160.711 47.685 ;
			RECT	160.847 47.621 160.879 47.685 ;
			RECT	161.015 47.621 161.047 47.685 ;
			RECT	161.183 47.621 161.215 47.685 ;
			RECT	161.351 47.621 161.383 47.685 ;
			RECT	161.519 47.621 161.551 47.685 ;
			RECT	161.687 47.621 161.719 47.685 ;
			RECT	161.855 47.621 161.887 47.685 ;
			RECT	162.023 47.621 162.055 47.685 ;
			RECT	162.191 47.621 162.223 47.685 ;
			RECT	162.359 47.621 162.391 47.685 ;
			RECT	162.527 47.621 162.559 47.685 ;
			RECT	162.695 47.621 162.727 47.685 ;
			RECT	162.863 47.621 162.895 47.685 ;
			RECT	163.031 47.621 163.063 47.685 ;
			RECT	163.199 47.621 163.231 47.685 ;
			RECT	163.367 47.621 163.399 47.685 ;
			RECT	163.535 47.621 163.567 47.685 ;
			RECT	163.703 47.621 163.735 47.685 ;
			RECT	163.871 47.621 163.903 47.685 ;
			RECT	164.039 47.621 164.071 47.685 ;
			RECT	164.207 47.621 164.239 47.685 ;
			RECT	164.375 47.621 164.407 47.685 ;
			RECT	164.543 47.621 164.575 47.685 ;
			RECT	164.711 47.621 164.743 47.685 ;
			RECT	164.879 47.621 164.911 47.685 ;
			RECT	165.047 47.621 165.079 47.685 ;
			RECT	165.215 47.621 165.247 47.685 ;
			RECT	165.383 47.621 165.415 47.685 ;
			RECT	165.551 47.621 165.583 47.685 ;
			RECT	165.719 47.621 165.751 47.685 ;
			RECT	165.887 47.621 165.919 47.685 ;
			RECT	166.055 47.621 166.087 47.685 ;
			RECT	166.223 47.621 166.255 47.685 ;
			RECT	166.391 47.621 166.423 47.685 ;
			RECT	166.559 47.621 166.591 47.685 ;
			RECT	166.727 47.621 166.759 47.685 ;
			RECT	166.895 47.621 166.927 47.685 ;
			RECT	167.063 47.621 167.095 47.685 ;
			RECT	167.231 47.621 167.263 47.685 ;
			RECT	167.399 47.621 167.431 47.685 ;
			RECT	167.567 47.621 167.599 47.685 ;
			RECT	167.735 47.621 167.767 47.685 ;
			RECT	167.903 47.621 167.935 47.685 ;
			RECT	168.071 47.621 168.103 47.685 ;
			RECT	168.239 47.621 168.271 47.685 ;
			RECT	168.407 47.621 168.439 47.685 ;
			RECT	168.575 47.621 168.607 47.685 ;
			RECT	168.743 47.621 168.775 47.685 ;
			RECT	168.911 47.621 168.943 47.685 ;
			RECT	169.079 47.621 169.111 47.685 ;
			RECT	169.247 47.621 169.279 47.685 ;
			RECT	169.415 47.621 169.447 47.685 ;
			RECT	169.583 47.621 169.615 47.685 ;
			RECT	169.751 47.621 169.783 47.685 ;
			RECT	169.919 47.621 169.951 47.685 ;
			RECT	170.087 47.621 170.119 47.685 ;
			RECT	170.255 47.621 170.287 47.685 ;
			RECT	170.423 47.621 170.455 47.685 ;
			RECT	170.591 47.621 170.623 47.685 ;
			RECT	170.759 47.621 170.791 47.685 ;
			RECT	170.927 47.621 170.959 47.685 ;
			RECT	171.095 47.621 171.127 47.685 ;
			RECT	171.263 47.621 171.295 47.685 ;
			RECT	171.431 47.621 171.463 47.685 ;
			RECT	171.599 47.621 171.631 47.685 ;
			RECT	171.767 47.621 171.799 47.685 ;
			RECT	171.935 47.621 171.967 47.685 ;
			RECT	172.103 47.621 172.135 47.685 ;
			RECT	172.271 47.621 172.303 47.685 ;
			RECT	172.439 47.621 172.471 47.685 ;
			RECT	172.607 47.621 172.639 47.685 ;
			RECT	172.775 47.621 172.807 47.685 ;
			RECT	172.943 47.621 172.975 47.685 ;
			RECT	173.111 47.621 173.143 47.685 ;
			RECT	173.279 47.621 173.311 47.685 ;
			RECT	173.447 47.621 173.479 47.685 ;
			RECT	173.615 47.621 173.647 47.685 ;
			RECT	173.783 47.621 173.815 47.685 ;
			RECT	173.951 47.621 173.983 47.685 ;
			RECT	174.119 47.621 174.151 47.685 ;
			RECT	174.287 47.621 174.319 47.685 ;
			RECT	174.455 47.621 174.487 47.685 ;
			RECT	174.623 47.621 174.655 47.685 ;
			RECT	174.791 47.621 174.823 47.685 ;
			RECT	174.959 47.621 174.991 47.685 ;
			RECT	175.127 47.621 175.159 47.685 ;
			RECT	175.295 47.621 175.327 47.685 ;
			RECT	175.463 47.621 175.495 47.685 ;
			RECT	175.631 47.621 175.663 47.685 ;
			RECT	175.799 47.621 175.831 47.685 ;
			RECT	175.967 47.621 175.999 47.685 ;
			RECT	176.135 47.621 176.167 47.685 ;
			RECT	176.303 47.621 176.335 47.685 ;
			RECT	176.471 47.621 176.503 47.685 ;
			RECT	176.639 47.621 176.671 47.685 ;
			RECT	176.807 47.621 176.839 47.685 ;
			RECT	176.975 47.621 177.007 47.685 ;
			RECT	177.143 47.621 177.175 47.685 ;
			RECT	177.311 47.621 177.343 47.685 ;
			RECT	177.479 47.621 177.511 47.685 ;
			RECT	177.647 47.621 177.679 47.685 ;
			RECT	177.815 47.621 177.847 47.685 ;
			RECT	177.983 47.621 178.015 47.685 ;
			RECT	178.151 47.621 178.183 47.685 ;
			RECT	178.319 47.621 178.351 47.685 ;
			RECT	178.487 47.621 178.519 47.685 ;
			RECT	178.655 47.621 178.687 47.685 ;
			RECT	178.823 47.621 178.855 47.685 ;
			RECT	178.991 47.621 179.023 47.685 ;
			RECT	179.159 47.621 179.191 47.685 ;
			RECT	179.327 47.621 179.359 47.685 ;
			RECT	179.495 47.621 179.527 47.685 ;
			RECT	179.663 47.621 179.695 47.685 ;
			RECT	179.831 47.621 179.863 47.685 ;
			RECT	179.999 47.621 180.031 47.685 ;
			RECT	180.167 47.621 180.199 47.685 ;
			RECT	180.335 47.621 180.367 47.685 ;
			RECT	180.503 47.621 180.535 47.685 ;
			RECT	180.671 47.621 180.703 47.685 ;
			RECT	180.839 47.621 180.871 47.685 ;
			RECT	181.007 47.621 181.039 47.685 ;
			RECT	181.175 47.621 181.207 47.685 ;
			RECT	181.343 47.621 181.375 47.685 ;
			RECT	181.511 47.621 181.543 47.685 ;
			RECT	181.679 47.621 181.711 47.685 ;
			RECT	181.847 47.621 181.879 47.685 ;
			RECT	182.015 47.621 182.047 47.685 ;
			RECT	182.183 47.621 182.215 47.685 ;
			RECT	182.351 47.621 182.383 47.685 ;
			RECT	182.519 47.621 182.551 47.685 ;
			RECT	182.687 47.621 182.719 47.685 ;
			RECT	182.855 47.621 182.887 47.685 ;
			RECT	183.023 47.621 183.055 47.685 ;
			RECT	183.191 47.621 183.223 47.685 ;
			RECT	183.359 47.621 183.391 47.685 ;
			RECT	183.527 47.621 183.559 47.685 ;
			RECT	183.695 47.621 183.727 47.685 ;
			RECT	183.863 47.621 183.895 47.685 ;
			RECT	184.031 47.621 184.063 47.685 ;
			RECT	184.199 47.621 184.231 47.685 ;
			RECT	184.367 47.621 184.399 47.685 ;
			RECT	184.535 47.621 184.567 47.685 ;
			RECT	184.703 47.621 184.735 47.685 ;
			RECT	184.871 47.621 184.903 47.685 ;
			RECT	185.039 47.621 185.071 47.685 ;
			RECT	185.207 47.621 185.239 47.685 ;
			RECT	185.375 47.621 185.407 47.685 ;
			RECT	185.543 47.621 185.575 47.685 ;
			RECT	185.711 47.621 185.743 47.685 ;
			RECT	185.879 47.621 185.911 47.685 ;
			RECT	186.047 47.621 186.079 47.685 ;
			RECT	186.215 47.621 186.247 47.685 ;
			RECT	186.383 47.621 186.415 47.685 ;
			RECT	186.551 47.621 186.583 47.685 ;
			RECT	186.719 47.621 186.751 47.685 ;
			RECT	186.887 47.621 186.919 47.685 ;
			RECT	187.055 47.621 187.087 47.685 ;
			RECT	187.223 47.621 187.255 47.685 ;
			RECT	187.391 47.621 187.423 47.685 ;
			RECT	187.559 47.621 187.591 47.685 ;
			RECT	187.727 47.621 187.759 47.685 ;
			RECT	187.895 47.621 187.927 47.685 ;
			RECT	188.063 47.621 188.095 47.685 ;
			RECT	188.231 47.621 188.263 47.685 ;
			RECT	188.399 47.621 188.431 47.685 ;
			RECT	188.567 47.621 188.599 47.685 ;
			RECT	188.735 47.621 188.767 47.685 ;
			RECT	188.903 47.621 188.935 47.685 ;
			RECT	189.071 47.621 189.103 47.685 ;
			RECT	189.239 47.621 189.271 47.685 ;
			RECT	189.407 47.621 189.439 47.685 ;
			RECT	189.575 47.621 189.607 47.685 ;
			RECT	189.743 47.621 189.775 47.685 ;
			RECT	189.911 47.621 189.943 47.685 ;
			RECT	190.079 47.621 190.111 47.685 ;
			RECT	190.247 47.621 190.279 47.685 ;
			RECT	190.415 47.621 190.447 47.685 ;
			RECT	190.583 47.621 190.615 47.685 ;
			RECT	190.751 47.621 190.783 47.685 ;
			RECT	190.919 47.621 190.951 47.685 ;
			RECT	191.087 47.621 191.119 47.685 ;
			RECT	191.255 47.621 191.287 47.685 ;
			RECT	191.423 47.621 191.455 47.685 ;
			RECT	191.591 47.621 191.623 47.685 ;
			RECT	191.759 47.621 191.791 47.685 ;
			RECT	191.927 47.621 191.959 47.685 ;
			RECT	192.095 47.621 192.127 47.685 ;
			RECT	192.263 47.621 192.295 47.685 ;
			RECT	192.431 47.621 192.463 47.685 ;
			RECT	192.599 47.621 192.631 47.685 ;
			RECT	192.767 47.621 192.799 47.685 ;
			RECT	192.935 47.621 192.967 47.685 ;
			RECT	193.103 47.621 193.135 47.685 ;
			RECT	193.271 47.621 193.303 47.685 ;
			RECT	193.439 47.621 193.471 47.685 ;
			RECT	193.607 47.621 193.639 47.685 ;
			RECT	193.775 47.621 193.807 47.685 ;
			RECT	193.943 47.621 193.975 47.685 ;
			RECT	194.111 47.621 194.143 47.685 ;
			RECT	194.279 47.621 194.311 47.685 ;
			RECT	194.447 47.621 194.479 47.685 ;
			RECT	194.615 47.621 194.647 47.685 ;
			RECT	194.783 47.621 194.815 47.685 ;
			RECT	194.951 47.621 194.983 47.685 ;
			RECT	195.119 47.621 195.151 47.685 ;
			RECT	195.287 47.621 195.319 47.685 ;
			RECT	195.455 47.621 195.487 47.685 ;
			RECT	195.623 47.621 195.655 47.685 ;
			RECT	195.791 47.621 195.823 47.685 ;
			RECT	195.959 47.621 195.991 47.685 ;
			RECT	196.127 47.621 196.159 47.685 ;
			RECT	196.295 47.621 196.327 47.685 ;
			RECT	196.463 47.621 196.495 47.685 ;
			RECT	196.631 47.621 196.663 47.685 ;
			RECT	196.799 47.621 196.831 47.685 ;
			RECT	196.967 47.621 196.999 47.685 ;
			RECT	197.135 47.621 197.167 47.685 ;
			RECT	197.303 47.621 197.335 47.685 ;
			RECT	197.471 47.621 197.503 47.685 ;
			RECT	197.639 47.621 197.671 47.685 ;
			RECT	197.807 47.621 197.839 47.685 ;
			RECT	197.975 47.621 198.007 47.685 ;
			RECT	198.143 47.621 198.175 47.685 ;
			RECT	198.311 47.621 198.343 47.685 ;
			RECT	198.479 47.621 198.511 47.685 ;
			RECT	198.647 47.621 198.679 47.685 ;
			RECT	198.815 47.621 198.847 47.685 ;
			RECT	198.983 47.621 199.015 47.685 ;
			RECT	199.151 47.621 199.183 47.685 ;
			RECT	199.319 47.621 199.351 47.685 ;
			RECT	199.487 47.621 199.519 47.685 ;
			RECT	199.655 47.621 199.687 47.685 ;
			RECT	199.823 47.621 199.855 47.685 ;
			RECT	199.991 47.621 200.023 47.685 ;
			RECT	200.362 47.621 200.394 47.685 ;
			RECT	200.9 47.621 200.932 47.685 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 48.003 201.665 48.123 ;
			LAYER	J3 ;
			RECT	1.661 48.031 1.693 48.095 ;
			RECT	2.323 48.031 2.387 48.095 ;
			RECT	3.451 48.031 3.483 48.095 ;
			RECT	4.179 48.047 4.211 48.079 ;
			RECT	4.568 48.047 4.632 48.079 ;
			RECT	4.805 48.031 4.837 48.095 ;
			RECT	4.96 48.031 4.992 48.095 ;
			RECT	5.252 48.031 5.284 48.095 ;
			RECT	5.808 48.047 5.84 48.079 ;
			RECT	6.179 48.031 6.211 48.095 ;
			RECT	6.347 48.031 6.379 48.095 ;
			RECT	6.515 48.031 6.547 48.095 ;
			RECT	6.683 48.031 6.715 48.095 ;
			RECT	6.851 48.031 6.883 48.095 ;
			RECT	7.019 48.031 7.051 48.095 ;
			RECT	7.187 48.031 7.219 48.095 ;
			RECT	7.355 48.031 7.387 48.095 ;
			RECT	7.523 48.031 7.555 48.095 ;
			RECT	7.691 48.031 7.723 48.095 ;
			RECT	7.859 48.031 7.891 48.095 ;
			RECT	8.027 48.031 8.059 48.095 ;
			RECT	8.195 48.031 8.227 48.095 ;
			RECT	8.363 48.031 8.395 48.095 ;
			RECT	8.531 48.031 8.563 48.095 ;
			RECT	8.699 48.031 8.731 48.095 ;
			RECT	8.867 48.031 8.899 48.095 ;
			RECT	9.035 48.031 9.067 48.095 ;
			RECT	9.203 48.031 9.235 48.095 ;
			RECT	9.371 48.031 9.403 48.095 ;
			RECT	9.539 48.031 9.571 48.095 ;
			RECT	9.707 48.031 9.739 48.095 ;
			RECT	9.875 48.031 9.907 48.095 ;
			RECT	10.043 48.031 10.075 48.095 ;
			RECT	10.211 48.031 10.243 48.095 ;
			RECT	10.379 48.031 10.411 48.095 ;
			RECT	10.547 48.031 10.579 48.095 ;
			RECT	10.715 48.031 10.747 48.095 ;
			RECT	10.883 48.031 10.915 48.095 ;
			RECT	11.051 48.031 11.083 48.095 ;
			RECT	11.219 48.031 11.251 48.095 ;
			RECT	11.387 48.031 11.419 48.095 ;
			RECT	11.555 48.031 11.587 48.095 ;
			RECT	11.723 48.031 11.755 48.095 ;
			RECT	11.891 48.031 11.923 48.095 ;
			RECT	12.059 48.031 12.091 48.095 ;
			RECT	12.227 48.031 12.259 48.095 ;
			RECT	12.395 48.031 12.427 48.095 ;
			RECT	12.563 48.031 12.595 48.095 ;
			RECT	12.731 48.031 12.763 48.095 ;
			RECT	12.899 48.031 12.931 48.095 ;
			RECT	13.067 48.031 13.099 48.095 ;
			RECT	13.235 48.031 13.267 48.095 ;
			RECT	13.403 48.031 13.435 48.095 ;
			RECT	13.571 48.031 13.603 48.095 ;
			RECT	13.739 48.031 13.771 48.095 ;
			RECT	13.907 48.031 13.939 48.095 ;
			RECT	14.075 48.031 14.107 48.095 ;
			RECT	14.243 48.031 14.275 48.095 ;
			RECT	14.411 48.031 14.443 48.095 ;
			RECT	14.579 48.031 14.611 48.095 ;
			RECT	14.747 48.031 14.779 48.095 ;
			RECT	14.915 48.031 14.947 48.095 ;
			RECT	15.083 48.031 15.115 48.095 ;
			RECT	15.251 48.031 15.283 48.095 ;
			RECT	15.419 48.031 15.451 48.095 ;
			RECT	15.587 48.031 15.619 48.095 ;
			RECT	15.755 48.031 15.787 48.095 ;
			RECT	15.923 48.031 15.955 48.095 ;
			RECT	16.091 48.031 16.123 48.095 ;
			RECT	16.259 48.031 16.291 48.095 ;
			RECT	16.427 48.031 16.459 48.095 ;
			RECT	16.595 48.031 16.627 48.095 ;
			RECT	16.763 48.031 16.795 48.095 ;
			RECT	16.931 48.031 16.963 48.095 ;
			RECT	17.099 48.031 17.131 48.095 ;
			RECT	17.267 48.031 17.299 48.095 ;
			RECT	17.435 48.031 17.467 48.095 ;
			RECT	17.603 48.031 17.635 48.095 ;
			RECT	17.771 48.031 17.803 48.095 ;
			RECT	17.939 48.031 17.971 48.095 ;
			RECT	18.107 48.031 18.139 48.095 ;
			RECT	18.275 48.031 18.307 48.095 ;
			RECT	18.443 48.031 18.475 48.095 ;
			RECT	18.611 48.031 18.643 48.095 ;
			RECT	18.779 48.031 18.811 48.095 ;
			RECT	18.947 48.031 18.979 48.095 ;
			RECT	19.115 48.031 19.147 48.095 ;
			RECT	19.283 48.031 19.315 48.095 ;
			RECT	19.451 48.031 19.483 48.095 ;
			RECT	19.619 48.031 19.651 48.095 ;
			RECT	19.787 48.031 19.819 48.095 ;
			RECT	19.955 48.031 19.987 48.095 ;
			RECT	20.123 48.031 20.155 48.095 ;
			RECT	20.291 48.031 20.323 48.095 ;
			RECT	20.459 48.031 20.491 48.095 ;
			RECT	20.627 48.031 20.659 48.095 ;
			RECT	20.795 48.031 20.827 48.095 ;
			RECT	20.963 48.031 20.995 48.095 ;
			RECT	21.131 48.031 21.163 48.095 ;
			RECT	21.299 48.031 21.331 48.095 ;
			RECT	21.467 48.031 21.499 48.095 ;
			RECT	21.635 48.031 21.667 48.095 ;
			RECT	21.803 48.031 21.835 48.095 ;
			RECT	21.971 48.031 22.003 48.095 ;
			RECT	22.139 48.031 22.171 48.095 ;
			RECT	22.307 48.031 22.339 48.095 ;
			RECT	22.475 48.031 22.507 48.095 ;
			RECT	22.643 48.031 22.675 48.095 ;
			RECT	22.811 48.031 22.843 48.095 ;
			RECT	22.979 48.031 23.011 48.095 ;
			RECT	23.147 48.031 23.179 48.095 ;
			RECT	23.315 48.031 23.347 48.095 ;
			RECT	23.483 48.031 23.515 48.095 ;
			RECT	23.651 48.031 23.683 48.095 ;
			RECT	23.819 48.031 23.851 48.095 ;
			RECT	23.987 48.031 24.019 48.095 ;
			RECT	24.155 48.031 24.187 48.095 ;
			RECT	24.323 48.031 24.355 48.095 ;
			RECT	24.491 48.031 24.523 48.095 ;
			RECT	24.659 48.031 24.691 48.095 ;
			RECT	24.827 48.031 24.859 48.095 ;
			RECT	24.995 48.031 25.027 48.095 ;
			RECT	25.163 48.031 25.195 48.095 ;
			RECT	25.331 48.031 25.363 48.095 ;
			RECT	25.499 48.031 25.531 48.095 ;
			RECT	25.667 48.031 25.699 48.095 ;
			RECT	25.835 48.031 25.867 48.095 ;
			RECT	26.003 48.031 26.035 48.095 ;
			RECT	26.171 48.031 26.203 48.095 ;
			RECT	26.339 48.031 26.371 48.095 ;
			RECT	26.507 48.031 26.539 48.095 ;
			RECT	26.675 48.031 26.707 48.095 ;
			RECT	26.843 48.031 26.875 48.095 ;
			RECT	27.011 48.031 27.043 48.095 ;
			RECT	27.179 48.031 27.211 48.095 ;
			RECT	27.347 48.031 27.379 48.095 ;
			RECT	27.515 48.031 27.547 48.095 ;
			RECT	27.683 48.031 27.715 48.095 ;
			RECT	27.851 48.031 27.883 48.095 ;
			RECT	28.019 48.031 28.051 48.095 ;
			RECT	28.187 48.031 28.219 48.095 ;
			RECT	28.355 48.031 28.387 48.095 ;
			RECT	28.523 48.031 28.555 48.095 ;
			RECT	28.691 48.031 28.723 48.095 ;
			RECT	28.859 48.031 28.891 48.095 ;
			RECT	29.027 48.031 29.059 48.095 ;
			RECT	29.195 48.031 29.227 48.095 ;
			RECT	29.363 48.031 29.395 48.095 ;
			RECT	29.531 48.031 29.563 48.095 ;
			RECT	29.699 48.031 29.731 48.095 ;
			RECT	29.867 48.031 29.899 48.095 ;
			RECT	30.035 48.031 30.067 48.095 ;
			RECT	30.203 48.031 30.235 48.095 ;
			RECT	30.371 48.031 30.403 48.095 ;
			RECT	30.539 48.031 30.571 48.095 ;
			RECT	30.707 48.031 30.739 48.095 ;
			RECT	30.875 48.031 30.907 48.095 ;
			RECT	31.043 48.031 31.075 48.095 ;
			RECT	31.211 48.031 31.243 48.095 ;
			RECT	31.379 48.031 31.411 48.095 ;
			RECT	31.547 48.031 31.579 48.095 ;
			RECT	31.715 48.031 31.747 48.095 ;
			RECT	31.883 48.031 31.915 48.095 ;
			RECT	32.051 48.031 32.083 48.095 ;
			RECT	32.219 48.031 32.251 48.095 ;
			RECT	32.387 48.031 32.419 48.095 ;
			RECT	32.555 48.031 32.587 48.095 ;
			RECT	32.723 48.031 32.755 48.095 ;
			RECT	32.891 48.031 32.923 48.095 ;
			RECT	33.059 48.031 33.091 48.095 ;
			RECT	33.227 48.031 33.259 48.095 ;
			RECT	33.395 48.031 33.427 48.095 ;
			RECT	33.563 48.031 33.595 48.095 ;
			RECT	33.731 48.031 33.763 48.095 ;
			RECT	33.899 48.031 33.931 48.095 ;
			RECT	34.067 48.031 34.099 48.095 ;
			RECT	34.235 48.031 34.267 48.095 ;
			RECT	34.403 48.031 34.435 48.095 ;
			RECT	34.571 48.031 34.603 48.095 ;
			RECT	34.739 48.031 34.771 48.095 ;
			RECT	34.907 48.031 34.939 48.095 ;
			RECT	35.075 48.031 35.107 48.095 ;
			RECT	35.243 48.031 35.275 48.095 ;
			RECT	35.411 48.031 35.443 48.095 ;
			RECT	35.579 48.031 35.611 48.095 ;
			RECT	35.747 48.031 35.779 48.095 ;
			RECT	35.915 48.031 35.947 48.095 ;
			RECT	36.083 48.031 36.115 48.095 ;
			RECT	36.251 48.031 36.283 48.095 ;
			RECT	36.419 48.031 36.451 48.095 ;
			RECT	36.587 48.031 36.619 48.095 ;
			RECT	36.755 48.031 36.787 48.095 ;
			RECT	36.923 48.031 36.955 48.095 ;
			RECT	37.091 48.031 37.123 48.095 ;
			RECT	37.259 48.031 37.291 48.095 ;
			RECT	37.427 48.031 37.459 48.095 ;
			RECT	37.595 48.031 37.627 48.095 ;
			RECT	37.763 48.031 37.795 48.095 ;
			RECT	37.931 48.031 37.963 48.095 ;
			RECT	38.099 48.031 38.131 48.095 ;
			RECT	38.267 48.031 38.299 48.095 ;
			RECT	38.435 48.031 38.467 48.095 ;
			RECT	38.603 48.031 38.635 48.095 ;
			RECT	38.771 48.031 38.803 48.095 ;
			RECT	38.939 48.031 38.971 48.095 ;
			RECT	39.107 48.031 39.139 48.095 ;
			RECT	39.275 48.031 39.307 48.095 ;
			RECT	39.443 48.031 39.475 48.095 ;
			RECT	39.611 48.031 39.643 48.095 ;
			RECT	39.779 48.031 39.811 48.095 ;
			RECT	39.947 48.031 39.979 48.095 ;
			RECT	40.115 48.031 40.147 48.095 ;
			RECT	40.283 48.031 40.315 48.095 ;
			RECT	40.451 48.031 40.483 48.095 ;
			RECT	40.619 48.031 40.651 48.095 ;
			RECT	40.787 48.031 40.819 48.095 ;
			RECT	40.955 48.031 40.987 48.095 ;
			RECT	41.123 48.031 41.155 48.095 ;
			RECT	41.291 48.031 41.323 48.095 ;
			RECT	41.459 48.031 41.491 48.095 ;
			RECT	41.627 48.031 41.659 48.095 ;
			RECT	41.795 48.031 41.827 48.095 ;
			RECT	41.963 48.031 41.995 48.095 ;
			RECT	42.131 48.031 42.163 48.095 ;
			RECT	42.299 48.031 42.331 48.095 ;
			RECT	42.467 48.031 42.499 48.095 ;
			RECT	42.635 48.031 42.667 48.095 ;
			RECT	42.803 48.031 42.835 48.095 ;
			RECT	42.971 48.031 43.003 48.095 ;
			RECT	43.139 48.031 43.171 48.095 ;
			RECT	43.307 48.031 43.339 48.095 ;
			RECT	43.475 48.031 43.507 48.095 ;
			RECT	43.643 48.031 43.675 48.095 ;
			RECT	43.811 48.031 43.843 48.095 ;
			RECT	43.979 48.031 44.011 48.095 ;
			RECT	44.147 48.031 44.179 48.095 ;
			RECT	44.315 48.031 44.347 48.095 ;
			RECT	44.483 48.031 44.515 48.095 ;
			RECT	44.651 48.031 44.683 48.095 ;
			RECT	44.819 48.031 44.851 48.095 ;
			RECT	44.987 48.031 45.019 48.095 ;
			RECT	45.155 48.031 45.187 48.095 ;
			RECT	45.323 48.031 45.355 48.095 ;
			RECT	45.491 48.031 45.523 48.095 ;
			RECT	45.659 48.031 45.691 48.095 ;
			RECT	45.827 48.031 45.859 48.095 ;
			RECT	45.995 48.031 46.027 48.095 ;
			RECT	46.163 48.031 46.195 48.095 ;
			RECT	46.331 48.031 46.363 48.095 ;
			RECT	46.499 48.031 46.531 48.095 ;
			RECT	46.667 48.031 46.699 48.095 ;
			RECT	46.835 48.031 46.867 48.095 ;
			RECT	47.003 48.031 47.035 48.095 ;
			RECT	47.171 48.031 47.203 48.095 ;
			RECT	47.339 48.031 47.371 48.095 ;
			RECT	47.507 48.031 47.539 48.095 ;
			RECT	47.675 48.031 47.707 48.095 ;
			RECT	47.843 48.031 47.875 48.095 ;
			RECT	48.011 48.031 48.043 48.095 ;
			RECT	48.179 48.031 48.211 48.095 ;
			RECT	48.347 48.031 48.379 48.095 ;
			RECT	48.515 48.031 48.547 48.095 ;
			RECT	48.683 48.031 48.715 48.095 ;
			RECT	48.851 48.031 48.883 48.095 ;
			RECT	49.019 48.031 49.051 48.095 ;
			RECT	49.187 48.031 49.219 48.095 ;
			RECT	49.557 48.047 49.589 48.079 ;
			RECT	51.92 48.031 51.952 48.095 ;
			RECT	52.96 48.031 53.024 48.095 ;
			RECT	53.91 48.031 53.942 48.095 ;
			RECT	54.251 48.031 54.283 48.095 ;
			RECT	54.812 48.031 54.844 48.095 ;
			RECT	55.562 48.031 55.626 48.095 ;
			RECT	55.842 48.031 55.874 48.095 ;
			RECT	55.969 48.031 56.033 48.095 ;
			RECT	57.372 48.031 57.404 48.095 ;
			RECT	58.615 48.047 58.647 48.079 ;
			RECT	58.985 48.031 59.017 48.095 ;
			RECT	59.153 48.031 59.185 48.095 ;
			RECT	59.321 48.031 59.353 48.095 ;
			RECT	59.489 48.031 59.521 48.095 ;
			RECT	59.657 48.031 59.689 48.095 ;
			RECT	59.825 48.031 59.857 48.095 ;
			RECT	59.993 48.031 60.025 48.095 ;
			RECT	60.161 48.031 60.193 48.095 ;
			RECT	60.329 48.031 60.361 48.095 ;
			RECT	60.497 48.031 60.529 48.095 ;
			RECT	60.665 48.031 60.697 48.095 ;
			RECT	60.833 48.031 60.865 48.095 ;
			RECT	61.001 48.031 61.033 48.095 ;
			RECT	61.169 48.031 61.201 48.095 ;
			RECT	61.337 48.031 61.369 48.095 ;
			RECT	61.505 48.031 61.537 48.095 ;
			RECT	61.673 48.031 61.705 48.095 ;
			RECT	61.841 48.031 61.873 48.095 ;
			RECT	62.009 48.031 62.041 48.095 ;
			RECT	62.177 48.031 62.209 48.095 ;
			RECT	62.345 48.031 62.377 48.095 ;
			RECT	62.513 48.031 62.545 48.095 ;
			RECT	62.681 48.031 62.713 48.095 ;
			RECT	62.849 48.031 62.881 48.095 ;
			RECT	63.017 48.031 63.049 48.095 ;
			RECT	63.185 48.031 63.217 48.095 ;
			RECT	63.353 48.031 63.385 48.095 ;
			RECT	63.521 48.031 63.553 48.095 ;
			RECT	63.689 48.031 63.721 48.095 ;
			RECT	63.857 48.031 63.889 48.095 ;
			RECT	64.025 48.031 64.057 48.095 ;
			RECT	64.193 48.031 64.225 48.095 ;
			RECT	64.361 48.031 64.393 48.095 ;
			RECT	64.529 48.031 64.561 48.095 ;
			RECT	64.697 48.031 64.729 48.095 ;
			RECT	64.865 48.031 64.897 48.095 ;
			RECT	65.033 48.031 65.065 48.095 ;
			RECT	65.201 48.031 65.233 48.095 ;
			RECT	65.369 48.031 65.401 48.095 ;
			RECT	65.537 48.031 65.569 48.095 ;
			RECT	65.705 48.031 65.737 48.095 ;
			RECT	65.873 48.031 65.905 48.095 ;
			RECT	66.041 48.031 66.073 48.095 ;
			RECT	66.209 48.031 66.241 48.095 ;
			RECT	66.377 48.031 66.409 48.095 ;
			RECT	66.545 48.031 66.577 48.095 ;
			RECT	66.713 48.031 66.745 48.095 ;
			RECT	66.881 48.031 66.913 48.095 ;
			RECT	67.049 48.031 67.081 48.095 ;
			RECT	67.217 48.031 67.249 48.095 ;
			RECT	67.385 48.031 67.417 48.095 ;
			RECT	67.553 48.031 67.585 48.095 ;
			RECT	67.721 48.031 67.753 48.095 ;
			RECT	67.889 48.031 67.921 48.095 ;
			RECT	68.057 48.031 68.089 48.095 ;
			RECT	68.225 48.031 68.257 48.095 ;
			RECT	68.393 48.031 68.425 48.095 ;
			RECT	68.561 48.031 68.593 48.095 ;
			RECT	68.729 48.031 68.761 48.095 ;
			RECT	68.897 48.031 68.929 48.095 ;
			RECT	69.065 48.031 69.097 48.095 ;
			RECT	69.233 48.031 69.265 48.095 ;
			RECT	69.401 48.031 69.433 48.095 ;
			RECT	69.569 48.031 69.601 48.095 ;
			RECT	69.737 48.031 69.769 48.095 ;
			RECT	69.905 48.031 69.937 48.095 ;
			RECT	70.073 48.031 70.105 48.095 ;
			RECT	70.241 48.031 70.273 48.095 ;
			RECT	70.409 48.031 70.441 48.095 ;
			RECT	70.577 48.031 70.609 48.095 ;
			RECT	70.745 48.031 70.777 48.095 ;
			RECT	70.913 48.031 70.945 48.095 ;
			RECT	71.081 48.031 71.113 48.095 ;
			RECT	71.249 48.031 71.281 48.095 ;
			RECT	71.417 48.031 71.449 48.095 ;
			RECT	71.585 48.031 71.617 48.095 ;
			RECT	71.753 48.031 71.785 48.095 ;
			RECT	71.921 48.031 71.953 48.095 ;
			RECT	72.089 48.031 72.121 48.095 ;
			RECT	72.257 48.031 72.289 48.095 ;
			RECT	72.425 48.031 72.457 48.095 ;
			RECT	72.593 48.031 72.625 48.095 ;
			RECT	72.761 48.031 72.793 48.095 ;
			RECT	72.929 48.031 72.961 48.095 ;
			RECT	73.097 48.031 73.129 48.095 ;
			RECT	73.265 48.031 73.297 48.095 ;
			RECT	73.433 48.031 73.465 48.095 ;
			RECT	73.601 48.031 73.633 48.095 ;
			RECT	73.769 48.031 73.801 48.095 ;
			RECT	73.937 48.031 73.969 48.095 ;
			RECT	74.105 48.031 74.137 48.095 ;
			RECT	74.273 48.031 74.305 48.095 ;
			RECT	74.441 48.031 74.473 48.095 ;
			RECT	74.609 48.031 74.641 48.095 ;
			RECT	74.777 48.031 74.809 48.095 ;
			RECT	74.945 48.031 74.977 48.095 ;
			RECT	75.113 48.031 75.145 48.095 ;
			RECT	75.281 48.031 75.313 48.095 ;
			RECT	75.449 48.031 75.481 48.095 ;
			RECT	75.617 48.031 75.649 48.095 ;
			RECT	75.785 48.031 75.817 48.095 ;
			RECT	75.953 48.031 75.985 48.095 ;
			RECT	76.121 48.031 76.153 48.095 ;
			RECT	76.289 48.031 76.321 48.095 ;
			RECT	76.457 48.031 76.489 48.095 ;
			RECT	76.625 48.031 76.657 48.095 ;
			RECT	76.793 48.031 76.825 48.095 ;
			RECT	76.961 48.031 76.993 48.095 ;
			RECT	77.129 48.031 77.161 48.095 ;
			RECT	77.297 48.031 77.329 48.095 ;
			RECT	77.465 48.031 77.497 48.095 ;
			RECT	77.633 48.031 77.665 48.095 ;
			RECT	77.801 48.031 77.833 48.095 ;
			RECT	77.969 48.031 78.001 48.095 ;
			RECT	78.137 48.031 78.169 48.095 ;
			RECT	78.305 48.031 78.337 48.095 ;
			RECT	78.473 48.031 78.505 48.095 ;
			RECT	78.641 48.031 78.673 48.095 ;
			RECT	78.809 48.031 78.841 48.095 ;
			RECT	78.977 48.031 79.009 48.095 ;
			RECT	79.145 48.031 79.177 48.095 ;
			RECT	79.313 48.031 79.345 48.095 ;
			RECT	79.481 48.031 79.513 48.095 ;
			RECT	79.649 48.031 79.681 48.095 ;
			RECT	79.817 48.031 79.849 48.095 ;
			RECT	79.985 48.031 80.017 48.095 ;
			RECT	80.153 48.031 80.185 48.095 ;
			RECT	80.321 48.031 80.353 48.095 ;
			RECT	80.489 48.031 80.521 48.095 ;
			RECT	80.657 48.031 80.689 48.095 ;
			RECT	80.825 48.031 80.857 48.095 ;
			RECT	80.993 48.031 81.025 48.095 ;
			RECT	81.161 48.031 81.193 48.095 ;
			RECT	81.329 48.031 81.361 48.095 ;
			RECT	81.497 48.031 81.529 48.095 ;
			RECT	81.665 48.031 81.697 48.095 ;
			RECT	81.833 48.031 81.865 48.095 ;
			RECT	82.001 48.031 82.033 48.095 ;
			RECT	82.169 48.031 82.201 48.095 ;
			RECT	82.337 48.031 82.369 48.095 ;
			RECT	82.505 48.031 82.537 48.095 ;
			RECT	82.673 48.031 82.705 48.095 ;
			RECT	82.841 48.031 82.873 48.095 ;
			RECT	83.009 48.031 83.041 48.095 ;
			RECT	83.177 48.031 83.209 48.095 ;
			RECT	83.345 48.031 83.377 48.095 ;
			RECT	83.513 48.031 83.545 48.095 ;
			RECT	83.681 48.031 83.713 48.095 ;
			RECT	83.849 48.031 83.881 48.095 ;
			RECT	84.017 48.031 84.049 48.095 ;
			RECT	84.185 48.031 84.217 48.095 ;
			RECT	84.353 48.031 84.385 48.095 ;
			RECT	84.521 48.031 84.553 48.095 ;
			RECT	84.689 48.031 84.721 48.095 ;
			RECT	84.857 48.031 84.889 48.095 ;
			RECT	85.025 48.031 85.057 48.095 ;
			RECT	85.193 48.031 85.225 48.095 ;
			RECT	85.361 48.031 85.393 48.095 ;
			RECT	85.529 48.031 85.561 48.095 ;
			RECT	85.697 48.031 85.729 48.095 ;
			RECT	85.865 48.031 85.897 48.095 ;
			RECT	86.033 48.031 86.065 48.095 ;
			RECT	86.201 48.031 86.233 48.095 ;
			RECT	86.369 48.031 86.401 48.095 ;
			RECT	86.537 48.031 86.569 48.095 ;
			RECT	86.705 48.031 86.737 48.095 ;
			RECT	86.873 48.031 86.905 48.095 ;
			RECT	87.041 48.031 87.073 48.095 ;
			RECT	87.209 48.031 87.241 48.095 ;
			RECT	87.377 48.031 87.409 48.095 ;
			RECT	87.545 48.031 87.577 48.095 ;
			RECT	87.713 48.031 87.745 48.095 ;
			RECT	87.881 48.031 87.913 48.095 ;
			RECT	88.049 48.031 88.081 48.095 ;
			RECT	88.217 48.031 88.249 48.095 ;
			RECT	88.385 48.031 88.417 48.095 ;
			RECT	88.553 48.031 88.585 48.095 ;
			RECT	88.721 48.031 88.753 48.095 ;
			RECT	88.889 48.031 88.921 48.095 ;
			RECT	89.057 48.031 89.089 48.095 ;
			RECT	89.225 48.031 89.257 48.095 ;
			RECT	89.393 48.031 89.425 48.095 ;
			RECT	89.561 48.031 89.593 48.095 ;
			RECT	89.729 48.031 89.761 48.095 ;
			RECT	89.897 48.031 89.929 48.095 ;
			RECT	90.065 48.031 90.097 48.095 ;
			RECT	90.233 48.031 90.265 48.095 ;
			RECT	90.401 48.031 90.433 48.095 ;
			RECT	90.569 48.031 90.601 48.095 ;
			RECT	90.737 48.031 90.769 48.095 ;
			RECT	90.905 48.031 90.937 48.095 ;
			RECT	91.073 48.031 91.105 48.095 ;
			RECT	91.241 48.031 91.273 48.095 ;
			RECT	91.409 48.031 91.441 48.095 ;
			RECT	91.577 48.031 91.609 48.095 ;
			RECT	91.745 48.031 91.777 48.095 ;
			RECT	91.913 48.031 91.945 48.095 ;
			RECT	92.081 48.031 92.113 48.095 ;
			RECT	92.249 48.031 92.281 48.095 ;
			RECT	92.417 48.031 92.449 48.095 ;
			RECT	92.585 48.031 92.617 48.095 ;
			RECT	92.753 48.031 92.785 48.095 ;
			RECT	92.921 48.031 92.953 48.095 ;
			RECT	93.089 48.031 93.121 48.095 ;
			RECT	93.257 48.031 93.289 48.095 ;
			RECT	93.425 48.031 93.457 48.095 ;
			RECT	93.593 48.031 93.625 48.095 ;
			RECT	93.761 48.031 93.793 48.095 ;
			RECT	93.929 48.031 93.961 48.095 ;
			RECT	94.097 48.031 94.129 48.095 ;
			RECT	94.265 48.031 94.297 48.095 ;
			RECT	94.433 48.031 94.465 48.095 ;
			RECT	94.601 48.031 94.633 48.095 ;
			RECT	94.769 48.031 94.801 48.095 ;
			RECT	94.937 48.031 94.969 48.095 ;
			RECT	95.105 48.031 95.137 48.095 ;
			RECT	95.273 48.031 95.305 48.095 ;
			RECT	95.441 48.031 95.473 48.095 ;
			RECT	95.609 48.031 95.641 48.095 ;
			RECT	95.777 48.031 95.809 48.095 ;
			RECT	95.945 48.031 95.977 48.095 ;
			RECT	96.113 48.031 96.145 48.095 ;
			RECT	96.281 48.031 96.313 48.095 ;
			RECT	96.449 48.031 96.481 48.095 ;
			RECT	96.617 48.031 96.649 48.095 ;
			RECT	96.785 48.031 96.817 48.095 ;
			RECT	96.953 48.031 96.985 48.095 ;
			RECT	97.121 48.031 97.153 48.095 ;
			RECT	97.289 48.031 97.321 48.095 ;
			RECT	97.457 48.031 97.489 48.095 ;
			RECT	97.625 48.031 97.657 48.095 ;
			RECT	97.793 48.031 97.825 48.095 ;
			RECT	97.961 48.031 97.993 48.095 ;
			RECT	98.129 48.031 98.161 48.095 ;
			RECT	98.297 48.031 98.329 48.095 ;
			RECT	98.465 48.031 98.497 48.095 ;
			RECT	98.633 48.031 98.665 48.095 ;
			RECT	98.801 48.031 98.833 48.095 ;
			RECT	98.969 48.031 99.001 48.095 ;
			RECT	99.137 48.031 99.169 48.095 ;
			RECT	99.305 48.031 99.337 48.095 ;
			RECT	99.473 48.031 99.505 48.095 ;
			RECT	99.641 48.031 99.673 48.095 ;
			RECT	99.809 48.031 99.841 48.095 ;
			RECT	99.977 48.031 100.009 48.095 ;
			RECT	100.145 48.031 100.177 48.095 ;
			RECT	100.313 48.031 100.345 48.095 ;
			RECT	100.481 48.031 100.513 48.095 ;
			RECT	100.649 48.031 100.681 48.095 ;
			RECT	100.817 48.031 100.849 48.095 ;
			RECT	100.985 48.031 101.017 48.095 ;
			RECT	101.153 48.031 101.185 48.095 ;
			RECT	101.321 48.031 101.353 48.095 ;
			RECT	101.489 48.031 101.521 48.095 ;
			RECT	101.657 48.031 101.689 48.095 ;
			RECT	101.825 48.031 101.857 48.095 ;
			RECT	101.993 48.031 102.025 48.095 ;
			RECT	102.364 48.047 102.396 48.079 ;
			RECT	103.806 48.047 103.838 48.079 ;
			RECT	104.177 48.031 104.209 48.095 ;
			RECT	104.345 48.031 104.377 48.095 ;
			RECT	104.513 48.031 104.545 48.095 ;
			RECT	104.681 48.031 104.713 48.095 ;
			RECT	104.849 48.031 104.881 48.095 ;
			RECT	105.017 48.031 105.049 48.095 ;
			RECT	105.185 48.031 105.217 48.095 ;
			RECT	105.353 48.031 105.385 48.095 ;
			RECT	105.521 48.031 105.553 48.095 ;
			RECT	105.689 48.031 105.721 48.095 ;
			RECT	105.857 48.031 105.889 48.095 ;
			RECT	106.025 48.031 106.057 48.095 ;
			RECT	106.193 48.031 106.225 48.095 ;
			RECT	106.361 48.031 106.393 48.095 ;
			RECT	106.529 48.031 106.561 48.095 ;
			RECT	106.697 48.031 106.729 48.095 ;
			RECT	106.865 48.031 106.897 48.095 ;
			RECT	107.033 48.031 107.065 48.095 ;
			RECT	107.201 48.031 107.233 48.095 ;
			RECT	107.369 48.031 107.401 48.095 ;
			RECT	107.537 48.031 107.569 48.095 ;
			RECT	107.705 48.031 107.737 48.095 ;
			RECT	107.873 48.031 107.905 48.095 ;
			RECT	108.041 48.031 108.073 48.095 ;
			RECT	108.209 48.031 108.241 48.095 ;
			RECT	108.377 48.031 108.409 48.095 ;
			RECT	108.545 48.031 108.577 48.095 ;
			RECT	108.713 48.031 108.745 48.095 ;
			RECT	108.881 48.031 108.913 48.095 ;
			RECT	109.049 48.031 109.081 48.095 ;
			RECT	109.217 48.031 109.249 48.095 ;
			RECT	109.385 48.031 109.417 48.095 ;
			RECT	109.553 48.031 109.585 48.095 ;
			RECT	109.721 48.031 109.753 48.095 ;
			RECT	109.889 48.031 109.921 48.095 ;
			RECT	110.057 48.031 110.089 48.095 ;
			RECT	110.225 48.031 110.257 48.095 ;
			RECT	110.393 48.031 110.425 48.095 ;
			RECT	110.561 48.031 110.593 48.095 ;
			RECT	110.729 48.031 110.761 48.095 ;
			RECT	110.897 48.031 110.929 48.095 ;
			RECT	111.065 48.031 111.097 48.095 ;
			RECT	111.233 48.031 111.265 48.095 ;
			RECT	111.401 48.031 111.433 48.095 ;
			RECT	111.569 48.031 111.601 48.095 ;
			RECT	111.737 48.031 111.769 48.095 ;
			RECT	111.905 48.031 111.937 48.095 ;
			RECT	112.073 48.031 112.105 48.095 ;
			RECT	112.241 48.031 112.273 48.095 ;
			RECT	112.409 48.031 112.441 48.095 ;
			RECT	112.577 48.031 112.609 48.095 ;
			RECT	112.745 48.031 112.777 48.095 ;
			RECT	112.913 48.031 112.945 48.095 ;
			RECT	113.081 48.031 113.113 48.095 ;
			RECT	113.249 48.031 113.281 48.095 ;
			RECT	113.417 48.031 113.449 48.095 ;
			RECT	113.585 48.031 113.617 48.095 ;
			RECT	113.753 48.031 113.785 48.095 ;
			RECT	113.921 48.031 113.953 48.095 ;
			RECT	114.089 48.031 114.121 48.095 ;
			RECT	114.257 48.031 114.289 48.095 ;
			RECT	114.425 48.031 114.457 48.095 ;
			RECT	114.593 48.031 114.625 48.095 ;
			RECT	114.761 48.031 114.793 48.095 ;
			RECT	114.929 48.031 114.961 48.095 ;
			RECT	115.097 48.031 115.129 48.095 ;
			RECT	115.265 48.031 115.297 48.095 ;
			RECT	115.433 48.031 115.465 48.095 ;
			RECT	115.601 48.031 115.633 48.095 ;
			RECT	115.769 48.031 115.801 48.095 ;
			RECT	115.937 48.031 115.969 48.095 ;
			RECT	116.105 48.031 116.137 48.095 ;
			RECT	116.273 48.031 116.305 48.095 ;
			RECT	116.441 48.031 116.473 48.095 ;
			RECT	116.609 48.031 116.641 48.095 ;
			RECT	116.777 48.031 116.809 48.095 ;
			RECT	116.945 48.031 116.977 48.095 ;
			RECT	117.113 48.031 117.145 48.095 ;
			RECT	117.281 48.031 117.313 48.095 ;
			RECT	117.449 48.031 117.481 48.095 ;
			RECT	117.617 48.031 117.649 48.095 ;
			RECT	117.785 48.031 117.817 48.095 ;
			RECT	117.953 48.031 117.985 48.095 ;
			RECT	118.121 48.031 118.153 48.095 ;
			RECT	118.289 48.031 118.321 48.095 ;
			RECT	118.457 48.031 118.489 48.095 ;
			RECT	118.625 48.031 118.657 48.095 ;
			RECT	118.793 48.031 118.825 48.095 ;
			RECT	118.961 48.031 118.993 48.095 ;
			RECT	119.129 48.031 119.161 48.095 ;
			RECT	119.297 48.031 119.329 48.095 ;
			RECT	119.465 48.031 119.497 48.095 ;
			RECT	119.633 48.031 119.665 48.095 ;
			RECT	119.801 48.031 119.833 48.095 ;
			RECT	119.969 48.031 120.001 48.095 ;
			RECT	120.137 48.031 120.169 48.095 ;
			RECT	120.305 48.031 120.337 48.095 ;
			RECT	120.473 48.031 120.505 48.095 ;
			RECT	120.641 48.031 120.673 48.095 ;
			RECT	120.809 48.031 120.841 48.095 ;
			RECT	120.977 48.031 121.009 48.095 ;
			RECT	121.145 48.031 121.177 48.095 ;
			RECT	121.313 48.031 121.345 48.095 ;
			RECT	121.481 48.031 121.513 48.095 ;
			RECT	121.649 48.031 121.681 48.095 ;
			RECT	121.817 48.031 121.849 48.095 ;
			RECT	121.985 48.031 122.017 48.095 ;
			RECT	122.153 48.031 122.185 48.095 ;
			RECT	122.321 48.031 122.353 48.095 ;
			RECT	122.489 48.031 122.521 48.095 ;
			RECT	122.657 48.031 122.689 48.095 ;
			RECT	122.825 48.031 122.857 48.095 ;
			RECT	122.993 48.031 123.025 48.095 ;
			RECT	123.161 48.031 123.193 48.095 ;
			RECT	123.329 48.031 123.361 48.095 ;
			RECT	123.497 48.031 123.529 48.095 ;
			RECT	123.665 48.031 123.697 48.095 ;
			RECT	123.833 48.031 123.865 48.095 ;
			RECT	124.001 48.031 124.033 48.095 ;
			RECT	124.169 48.031 124.201 48.095 ;
			RECT	124.337 48.031 124.369 48.095 ;
			RECT	124.505 48.031 124.537 48.095 ;
			RECT	124.673 48.031 124.705 48.095 ;
			RECT	124.841 48.031 124.873 48.095 ;
			RECT	125.009 48.031 125.041 48.095 ;
			RECT	125.177 48.031 125.209 48.095 ;
			RECT	125.345 48.031 125.377 48.095 ;
			RECT	125.513 48.031 125.545 48.095 ;
			RECT	125.681 48.031 125.713 48.095 ;
			RECT	125.849 48.031 125.881 48.095 ;
			RECT	126.017 48.031 126.049 48.095 ;
			RECT	126.185 48.031 126.217 48.095 ;
			RECT	126.353 48.031 126.385 48.095 ;
			RECT	126.521 48.031 126.553 48.095 ;
			RECT	126.689 48.031 126.721 48.095 ;
			RECT	126.857 48.031 126.889 48.095 ;
			RECT	127.025 48.031 127.057 48.095 ;
			RECT	127.193 48.031 127.225 48.095 ;
			RECT	127.361 48.031 127.393 48.095 ;
			RECT	127.529 48.031 127.561 48.095 ;
			RECT	127.697 48.031 127.729 48.095 ;
			RECT	127.865 48.031 127.897 48.095 ;
			RECT	128.033 48.031 128.065 48.095 ;
			RECT	128.201 48.031 128.233 48.095 ;
			RECT	128.369 48.031 128.401 48.095 ;
			RECT	128.537 48.031 128.569 48.095 ;
			RECT	128.705 48.031 128.737 48.095 ;
			RECT	128.873 48.031 128.905 48.095 ;
			RECT	129.041 48.031 129.073 48.095 ;
			RECT	129.209 48.031 129.241 48.095 ;
			RECT	129.377 48.031 129.409 48.095 ;
			RECT	129.545 48.031 129.577 48.095 ;
			RECT	129.713 48.031 129.745 48.095 ;
			RECT	129.881 48.031 129.913 48.095 ;
			RECT	130.049 48.031 130.081 48.095 ;
			RECT	130.217 48.031 130.249 48.095 ;
			RECT	130.385 48.031 130.417 48.095 ;
			RECT	130.553 48.031 130.585 48.095 ;
			RECT	130.721 48.031 130.753 48.095 ;
			RECT	130.889 48.031 130.921 48.095 ;
			RECT	131.057 48.031 131.089 48.095 ;
			RECT	131.225 48.031 131.257 48.095 ;
			RECT	131.393 48.031 131.425 48.095 ;
			RECT	131.561 48.031 131.593 48.095 ;
			RECT	131.729 48.031 131.761 48.095 ;
			RECT	131.897 48.031 131.929 48.095 ;
			RECT	132.065 48.031 132.097 48.095 ;
			RECT	132.233 48.031 132.265 48.095 ;
			RECT	132.401 48.031 132.433 48.095 ;
			RECT	132.569 48.031 132.601 48.095 ;
			RECT	132.737 48.031 132.769 48.095 ;
			RECT	132.905 48.031 132.937 48.095 ;
			RECT	133.073 48.031 133.105 48.095 ;
			RECT	133.241 48.031 133.273 48.095 ;
			RECT	133.409 48.031 133.441 48.095 ;
			RECT	133.577 48.031 133.609 48.095 ;
			RECT	133.745 48.031 133.777 48.095 ;
			RECT	133.913 48.031 133.945 48.095 ;
			RECT	134.081 48.031 134.113 48.095 ;
			RECT	134.249 48.031 134.281 48.095 ;
			RECT	134.417 48.031 134.449 48.095 ;
			RECT	134.585 48.031 134.617 48.095 ;
			RECT	134.753 48.031 134.785 48.095 ;
			RECT	134.921 48.031 134.953 48.095 ;
			RECT	135.089 48.031 135.121 48.095 ;
			RECT	135.257 48.031 135.289 48.095 ;
			RECT	135.425 48.031 135.457 48.095 ;
			RECT	135.593 48.031 135.625 48.095 ;
			RECT	135.761 48.031 135.793 48.095 ;
			RECT	135.929 48.031 135.961 48.095 ;
			RECT	136.097 48.031 136.129 48.095 ;
			RECT	136.265 48.031 136.297 48.095 ;
			RECT	136.433 48.031 136.465 48.095 ;
			RECT	136.601 48.031 136.633 48.095 ;
			RECT	136.769 48.031 136.801 48.095 ;
			RECT	136.937 48.031 136.969 48.095 ;
			RECT	137.105 48.031 137.137 48.095 ;
			RECT	137.273 48.031 137.305 48.095 ;
			RECT	137.441 48.031 137.473 48.095 ;
			RECT	137.609 48.031 137.641 48.095 ;
			RECT	137.777 48.031 137.809 48.095 ;
			RECT	137.945 48.031 137.977 48.095 ;
			RECT	138.113 48.031 138.145 48.095 ;
			RECT	138.281 48.031 138.313 48.095 ;
			RECT	138.449 48.031 138.481 48.095 ;
			RECT	138.617 48.031 138.649 48.095 ;
			RECT	138.785 48.031 138.817 48.095 ;
			RECT	138.953 48.031 138.985 48.095 ;
			RECT	139.121 48.031 139.153 48.095 ;
			RECT	139.289 48.031 139.321 48.095 ;
			RECT	139.457 48.031 139.489 48.095 ;
			RECT	139.625 48.031 139.657 48.095 ;
			RECT	139.793 48.031 139.825 48.095 ;
			RECT	139.961 48.031 139.993 48.095 ;
			RECT	140.129 48.031 140.161 48.095 ;
			RECT	140.297 48.031 140.329 48.095 ;
			RECT	140.465 48.031 140.497 48.095 ;
			RECT	140.633 48.031 140.665 48.095 ;
			RECT	140.801 48.031 140.833 48.095 ;
			RECT	140.969 48.031 141.001 48.095 ;
			RECT	141.137 48.031 141.169 48.095 ;
			RECT	141.305 48.031 141.337 48.095 ;
			RECT	141.473 48.031 141.505 48.095 ;
			RECT	141.641 48.031 141.673 48.095 ;
			RECT	141.809 48.031 141.841 48.095 ;
			RECT	141.977 48.031 142.009 48.095 ;
			RECT	142.145 48.031 142.177 48.095 ;
			RECT	142.313 48.031 142.345 48.095 ;
			RECT	142.481 48.031 142.513 48.095 ;
			RECT	142.649 48.031 142.681 48.095 ;
			RECT	142.817 48.031 142.849 48.095 ;
			RECT	142.985 48.031 143.017 48.095 ;
			RECT	143.153 48.031 143.185 48.095 ;
			RECT	143.321 48.031 143.353 48.095 ;
			RECT	143.489 48.031 143.521 48.095 ;
			RECT	143.657 48.031 143.689 48.095 ;
			RECT	143.825 48.031 143.857 48.095 ;
			RECT	143.993 48.031 144.025 48.095 ;
			RECT	144.161 48.031 144.193 48.095 ;
			RECT	144.329 48.031 144.361 48.095 ;
			RECT	144.497 48.031 144.529 48.095 ;
			RECT	144.665 48.031 144.697 48.095 ;
			RECT	144.833 48.031 144.865 48.095 ;
			RECT	145.001 48.031 145.033 48.095 ;
			RECT	145.169 48.031 145.201 48.095 ;
			RECT	145.337 48.031 145.369 48.095 ;
			RECT	145.505 48.031 145.537 48.095 ;
			RECT	145.673 48.031 145.705 48.095 ;
			RECT	145.841 48.031 145.873 48.095 ;
			RECT	146.009 48.031 146.041 48.095 ;
			RECT	146.177 48.031 146.209 48.095 ;
			RECT	146.345 48.031 146.377 48.095 ;
			RECT	146.513 48.031 146.545 48.095 ;
			RECT	146.681 48.031 146.713 48.095 ;
			RECT	146.849 48.031 146.881 48.095 ;
			RECT	147.017 48.031 147.049 48.095 ;
			RECT	147.185 48.031 147.217 48.095 ;
			RECT	147.555 48.047 147.587 48.079 ;
			RECT	149.918 48.031 149.95 48.095 ;
			RECT	150.958 48.031 151.022 48.095 ;
			RECT	151.908 48.031 151.94 48.095 ;
			RECT	152.249 48.031 152.281 48.095 ;
			RECT	152.81 48.031 152.842 48.095 ;
			RECT	153.56 48.031 153.624 48.095 ;
			RECT	153.84 48.031 153.872 48.095 ;
			RECT	153.967 48.031 154.031 48.095 ;
			RECT	155.37 48.031 155.402 48.095 ;
			RECT	156.613 48.047 156.645 48.079 ;
			RECT	156.983 48.031 157.015 48.095 ;
			RECT	157.151 48.031 157.183 48.095 ;
			RECT	157.319 48.031 157.351 48.095 ;
			RECT	157.487 48.031 157.519 48.095 ;
			RECT	157.655 48.031 157.687 48.095 ;
			RECT	157.823 48.031 157.855 48.095 ;
			RECT	157.991 48.031 158.023 48.095 ;
			RECT	158.159 48.031 158.191 48.095 ;
			RECT	158.327 48.031 158.359 48.095 ;
			RECT	158.495 48.031 158.527 48.095 ;
			RECT	158.663 48.031 158.695 48.095 ;
			RECT	158.831 48.031 158.863 48.095 ;
			RECT	158.999 48.031 159.031 48.095 ;
			RECT	159.167 48.031 159.199 48.095 ;
			RECT	159.335 48.031 159.367 48.095 ;
			RECT	159.503 48.031 159.535 48.095 ;
			RECT	159.671 48.031 159.703 48.095 ;
			RECT	159.839 48.031 159.871 48.095 ;
			RECT	160.007 48.031 160.039 48.095 ;
			RECT	160.175 48.031 160.207 48.095 ;
			RECT	160.343 48.031 160.375 48.095 ;
			RECT	160.511 48.031 160.543 48.095 ;
			RECT	160.679 48.031 160.711 48.095 ;
			RECT	160.847 48.031 160.879 48.095 ;
			RECT	161.015 48.031 161.047 48.095 ;
			RECT	161.183 48.031 161.215 48.095 ;
			RECT	161.351 48.031 161.383 48.095 ;
			RECT	161.519 48.031 161.551 48.095 ;
			RECT	161.687 48.031 161.719 48.095 ;
			RECT	161.855 48.031 161.887 48.095 ;
			RECT	162.023 48.031 162.055 48.095 ;
			RECT	162.191 48.031 162.223 48.095 ;
			RECT	162.359 48.031 162.391 48.095 ;
			RECT	162.527 48.031 162.559 48.095 ;
			RECT	162.695 48.031 162.727 48.095 ;
			RECT	162.863 48.031 162.895 48.095 ;
			RECT	163.031 48.031 163.063 48.095 ;
			RECT	163.199 48.031 163.231 48.095 ;
			RECT	163.367 48.031 163.399 48.095 ;
			RECT	163.535 48.031 163.567 48.095 ;
			RECT	163.703 48.031 163.735 48.095 ;
			RECT	163.871 48.031 163.903 48.095 ;
			RECT	164.039 48.031 164.071 48.095 ;
			RECT	164.207 48.031 164.239 48.095 ;
			RECT	164.375 48.031 164.407 48.095 ;
			RECT	164.543 48.031 164.575 48.095 ;
			RECT	164.711 48.031 164.743 48.095 ;
			RECT	164.879 48.031 164.911 48.095 ;
			RECT	165.047 48.031 165.079 48.095 ;
			RECT	165.215 48.031 165.247 48.095 ;
			RECT	165.383 48.031 165.415 48.095 ;
			RECT	165.551 48.031 165.583 48.095 ;
			RECT	165.719 48.031 165.751 48.095 ;
			RECT	165.887 48.031 165.919 48.095 ;
			RECT	166.055 48.031 166.087 48.095 ;
			RECT	166.223 48.031 166.255 48.095 ;
			RECT	166.391 48.031 166.423 48.095 ;
			RECT	166.559 48.031 166.591 48.095 ;
			RECT	166.727 48.031 166.759 48.095 ;
			RECT	166.895 48.031 166.927 48.095 ;
			RECT	167.063 48.031 167.095 48.095 ;
			RECT	167.231 48.031 167.263 48.095 ;
			RECT	167.399 48.031 167.431 48.095 ;
			RECT	167.567 48.031 167.599 48.095 ;
			RECT	167.735 48.031 167.767 48.095 ;
			RECT	167.903 48.031 167.935 48.095 ;
			RECT	168.071 48.031 168.103 48.095 ;
			RECT	168.239 48.031 168.271 48.095 ;
			RECT	168.407 48.031 168.439 48.095 ;
			RECT	168.575 48.031 168.607 48.095 ;
			RECT	168.743 48.031 168.775 48.095 ;
			RECT	168.911 48.031 168.943 48.095 ;
			RECT	169.079 48.031 169.111 48.095 ;
			RECT	169.247 48.031 169.279 48.095 ;
			RECT	169.415 48.031 169.447 48.095 ;
			RECT	169.583 48.031 169.615 48.095 ;
			RECT	169.751 48.031 169.783 48.095 ;
			RECT	169.919 48.031 169.951 48.095 ;
			RECT	170.087 48.031 170.119 48.095 ;
			RECT	170.255 48.031 170.287 48.095 ;
			RECT	170.423 48.031 170.455 48.095 ;
			RECT	170.591 48.031 170.623 48.095 ;
			RECT	170.759 48.031 170.791 48.095 ;
			RECT	170.927 48.031 170.959 48.095 ;
			RECT	171.095 48.031 171.127 48.095 ;
			RECT	171.263 48.031 171.295 48.095 ;
			RECT	171.431 48.031 171.463 48.095 ;
			RECT	171.599 48.031 171.631 48.095 ;
			RECT	171.767 48.031 171.799 48.095 ;
			RECT	171.935 48.031 171.967 48.095 ;
			RECT	172.103 48.031 172.135 48.095 ;
			RECT	172.271 48.031 172.303 48.095 ;
			RECT	172.439 48.031 172.471 48.095 ;
			RECT	172.607 48.031 172.639 48.095 ;
			RECT	172.775 48.031 172.807 48.095 ;
			RECT	172.943 48.031 172.975 48.095 ;
			RECT	173.111 48.031 173.143 48.095 ;
			RECT	173.279 48.031 173.311 48.095 ;
			RECT	173.447 48.031 173.479 48.095 ;
			RECT	173.615 48.031 173.647 48.095 ;
			RECT	173.783 48.031 173.815 48.095 ;
			RECT	173.951 48.031 173.983 48.095 ;
			RECT	174.119 48.031 174.151 48.095 ;
			RECT	174.287 48.031 174.319 48.095 ;
			RECT	174.455 48.031 174.487 48.095 ;
			RECT	174.623 48.031 174.655 48.095 ;
			RECT	174.791 48.031 174.823 48.095 ;
			RECT	174.959 48.031 174.991 48.095 ;
			RECT	175.127 48.031 175.159 48.095 ;
			RECT	175.295 48.031 175.327 48.095 ;
			RECT	175.463 48.031 175.495 48.095 ;
			RECT	175.631 48.031 175.663 48.095 ;
			RECT	175.799 48.031 175.831 48.095 ;
			RECT	175.967 48.031 175.999 48.095 ;
			RECT	176.135 48.031 176.167 48.095 ;
			RECT	176.303 48.031 176.335 48.095 ;
			RECT	176.471 48.031 176.503 48.095 ;
			RECT	176.639 48.031 176.671 48.095 ;
			RECT	176.807 48.031 176.839 48.095 ;
			RECT	176.975 48.031 177.007 48.095 ;
			RECT	177.143 48.031 177.175 48.095 ;
			RECT	177.311 48.031 177.343 48.095 ;
			RECT	177.479 48.031 177.511 48.095 ;
			RECT	177.647 48.031 177.679 48.095 ;
			RECT	177.815 48.031 177.847 48.095 ;
			RECT	177.983 48.031 178.015 48.095 ;
			RECT	178.151 48.031 178.183 48.095 ;
			RECT	178.319 48.031 178.351 48.095 ;
			RECT	178.487 48.031 178.519 48.095 ;
			RECT	178.655 48.031 178.687 48.095 ;
			RECT	178.823 48.031 178.855 48.095 ;
			RECT	178.991 48.031 179.023 48.095 ;
			RECT	179.159 48.031 179.191 48.095 ;
			RECT	179.327 48.031 179.359 48.095 ;
			RECT	179.495 48.031 179.527 48.095 ;
			RECT	179.663 48.031 179.695 48.095 ;
			RECT	179.831 48.031 179.863 48.095 ;
			RECT	179.999 48.031 180.031 48.095 ;
			RECT	180.167 48.031 180.199 48.095 ;
			RECT	180.335 48.031 180.367 48.095 ;
			RECT	180.503 48.031 180.535 48.095 ;
			RECT	180.671 48.031 180.703 48.095 ;
			RECT	180.839 48.031 180.871 48.095 ;
			RECT	181.007 48.031 181.039 48.095 ;
			RECT	181.175 48.031 181.207 48.095 ;
			RECT	181.343 48.031 181.375 48.095 ;
			RECT	181.511 48.031 181.543 48.095 ;
			RECT	181.679 48.031 181.711 48.095 ;
			RECT	181.847 48.031 181.879 48.095 ;
			RECT	182.015 48.031 182.047 48.095 ;
			RECT	182.183 48.031 182.215 48.095 ;
			RECT	182.351 48.031 182.383 48.095 ;
			RECT	182.519 48.031 182.551 48.095 ;
			RECT	182.687 48.031 182.719 48.095 ;
			RECT	182.855 48.031 182.887 48.095 ;
			RECT	183.023 48.031 183.055 48.095 ;
			RECT	183.191 48.031 183.223 48.095 ;
			RECT	183.359 48.031 183.391 48.095 ;
			RECT	183.527 48.031 183.559 48.095 ;
			RECT	183.695 48.031 183.727 48.095 ;
			RECT	183.863 48.031 183.895 48.095 ;
			RECT	184.031 48.031 184.063 48.095 ;
			RECT	184.199 48.031 184.231 48.095 ;
			RECT	184.367 48.031 184.399 48.095 ;
			RECT	184.535 48.031 184.567 48.095 ;
			RECT	184.703 48.031 184.735 48.095 ;
			RECT	184.871 48.031 184.903 48.095 ;
			RECT	185.039 48.031 185.071 48.095 ;
			RECT	185.207 48.031 185.239 48.095 ;
			RECT	185.375 48.031 185.407 48.095 ;
			RECT	185.543 48.031 185.575 48.095 ;
			RECT	185.711 48.031 185.743 48.095 ;
			RECT	185.879 48.031 185.911 48.095 ;
			RECT	186.047 48.031 186.079 48.095 ;
			RECT	186.215 48.031 186.247 48.095 ;
			RECT	186.383 48.031 186.415 48.095 ;
			RECT	186.551 48.031 186.583 48.095 ;
			RECT	186.719 48.031 186.751 48.095 ;
			RECT	186.887 48.031 186.919 48.095 ;
			RECT	187.055 48.031 187.087 48.095 ;
			RECT	187.223 48.031 187.255 48.095 ;
			RECT	187.391 48.031 187.423 48.095 ;
			RECT	187.559 48.031 187.591 48.095 ;
			RECT	187.727 48.031 187.759 48.095 ;
			RECT	187.895 48.031 187.927 48.095 ;
			RECT	188.063 48.031 188.095 48.095 ;
			RECT	188.231 48.031 188.263 48.095 ;
			RECT	188.399 48.031 188.431 48.095 ;
			RECT	188.567 48.031 188.599 48.095 ;
			RECT	188.735 48.031 188.767 48.095 ;
			RECT	188.903 48.031 188.935 48.095 ;
			RECT	189.071 48.031 189.103 48.095 ;
			RECT	189.239 48.031 189.271 48.095 ;
			RECT	189.407 48.031 189.439 48.095 ;
			RECT	189.575 48.031 189.607 48.095 ;
			RECT	189.743 48.031 189.775 48.095 ;
			RECT	189.911 48.031 189.943 48.095 ;
			RECT	190.079 48.031 190.111 48.095 ;
			RECT	190.247 48.031 190.279 48.095 ;
			RECT	190.415 48.031 190.447 48.095 ;
			RECT	190.583 48.031 190.615 48.095 ;
			RECT	190.751 48.031 190.783 48.095 ;
			RECT	190.919 48.031 190.951 48.095 ;
			RECT	191.087 48.031 191.119 48.095 ;
			RECT	191.255 48.031 191.287 48.095 ;
			RECT	191.423 48.031 191.455 48.095 ;
			RECT	191.591 48.031 191.623 48.095 ;
			RECT	191.759 48.031 191.791 48.095 ;
			RECT	191.927 48.031 191.959 48.095 ;
			RECT	192.095 48.031 192.127 48.095 ;
			RECT	192.263 48.031 192.295 48.095 ;
			RECT	192.431 48.031 192.463 48.095 ;
			RECT	192.599 48.031 192.631 48.095 ;
			RECT	192.767 48.031 192.799 48.095 ;
			RECT	192.935 48.031 192.967 48.095 ;
			RECT	193.103 48.031 193.135 48.095 ;
			RECT	193.271 48.031 193.303 48.095 ;
			RECT	193.439 48.031 193.471 48.095 ;
			RECT	193.607 48.031 193.639 48.095 ;
			RECT	193.775 48.031 193.807 48.095 ;
			RECT	193.943 48.031 193.975 48.095 ;
			RECT	194.111 48.031 194.143 48.095 ;
			RECT	194.279 48.031 194.311 48.095 ;
			RECT	194.447 48.031 194.479 48.095 ;
			RECT	194.615 48.031 194.647 48.095 ;
			RECT	194.783 48.031 194.815 48.095 ;
			RECT	194.951 48.031 194.983 48.095 ;
			RECT	195.119 48.031 195.151 48.095 ;
			RECT	195.287 48.031 195.319 48.095 ;
			RECT	195.455 48.031 195.487 48.095 ;
			RECT	195.623 48.031 195.655 48.095 ;
			RECT	195.791 48.031 195.823 48.095 ;
			RECT	195.959 48.031 195.991 48.095 ;
			RECT	196.127 48.031 196.159 48.095 ;
			RECT	196.295 48.031 196.327 48.095 ;
			RECT	196.463 48.031 196.495 48.095 ;
			RECT	196.631 48.031 196.663 48.095 ;
			RECT	196.799 48.031 196.831 48.095 ;
			RECT	196.967 48.031 196.999 48.095 ;
			RECT	197.135 48.031 197.167 48.095 ;
			RECT	197.303 48.031 197.335 48.095 ;
			RECT	197.471 48.031 197.503 48.095 ;
			RECT	197.639 48.031 197.671 48.095 ;
			RECT	197.807 48.031 197.839 48.095 ;
			RECT	197.975 48.031 198.007 48.095 ;
			RECT	198.143 48.031 198.175 48.095 ;
			RECT	198.311 48.031 198.343 48.095 ;
			RECT	198.479 48.031 198.511 48.095 ;
			RECT	198.647 48.031 198.679 48.095 ;
			RECT	198.815 48.031 198.847 48.095 ;
			RECT	198.983 48.031 199.015 48.095 ;
			RECT	199.151 48.031 199.183 48.095 ;
			RECT	199.319 48.031 199.351 48.095 ;
			RECT	199.487 48.031 199.519 48.095 ;
			RECT	199.655 48.031 199.687 48.095 ;
			RECT	199.823 48.031 199.855 48.095 ;
			RECT	199.991 48.031 200.023 48.095 ;
			RECT	200.362 48.047 200.394 48.079 ;
			RECT	200.9 48.031 200.932 48.095 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 50.158 201.665 50.268 ;
			LAYER	J3 ;
			RECT	1.645 50.181 1.709 50.245 ;
			RECT	2.323 50.181 2.387 50.245 ;
			RECT	3.438 50.199 3.47 50.263 ;
			RECT	4.195 50.181 4.227 50.245 ;
			RECT	4.96 50.181 4.992 50.245 ;
			RECT	5.252 50.181 5.284 50.245 ;
			RECT	5.927 50.181 5.959 50.245 ;
			RECT	6.179 50.181 6.211 50.245 ;
			RECT	6.347 50.181 6.379 50.245 ;
			RECT	6.515 50.181 6.547 50.245 ;
			RECT	6.683 50.181 6.715 50.245 ;
			RECT	6.851 50.181 6.883 50.245 ;
			RECT	7.019 50.181 7.051 50.245 ;
			RECT	7.187 50.181 7.219 50.245 ;
			RECT	7.355 50.181 7.387 50.245 ;
			RECT	7.523 50.181 7.555 50.245 ;
			RECT	7.691 50.181 7.723 50.245 ;
			RECT	7.859 50.181 7.891 50.245 ;
			RECT	8.027 50.181 8.059 50.245 ;
			RECT	8.195 50.181 8.227 50.245 ;
			RECT	8.363 50.181 8.395 50.245 ;
			RECT	8.531 50.181 8.563 50.245 ;
			RECT	8.699 50.181 8.731 50.245 ;
			RECT	8.867 50.181 8.899 50.245 ;
			RECT	9.035 50.181 9.067 50.245 ;
			RECT	9.203 50.181 9.235 50.245 ;
			RECT	9.371 50.181 9.403 50.245 ;
			RECT	9.539 50.181 9.571 50.245 ;
			RECT	9.707 50.181 9.739 50.245 ;
			RECT	9.875 50.181 9.907 50.245 ;
			RECT	10.043 50.181 10.075 50.245 ;
			RECT	10.211 50.181 10.243 50.245 ;
			RECT	10.379 50.181 10.411 50.245 ;
			RECT	10.547 50.181 10.579 50.245 ;
			RECT	10.715 50.181 10.747 50.245 ;
			RECT	10.883 50.181 10.915 50.245 ;
			RECT	11.051 50.181 11.083 50.245 ;
			RECT	11.219 50.181 11.251 50.245 ;
			RECT	11.387 50.181 11.419 50.245 ;
			RECT	11.555 50.181 11.587 50.245 ;
			RECT	11.723 50.181 11.755 50.245 ;
			RECT	11.891 50.181 11.923 50.245 ;
			RECT	12.059 50.181 12.091 50.245 ;
			RECT	12.227 50.181 12.259 50.245 ;
			RECT	12.395 50.181 12.427 50.245 ;
			RECT	12.563 50.181 12.595 50.245 ;
			RECT	12.731 50.181 12.763 50.245 ;
			RECT	12.899 50.181 12.931 50.245 ;
			RECT	13.067 50.181 13.099 50.245 ;
			RECT	13.235 50.181 13.267 50.245 ;
			RECT	13.403 50.181 13.435 50.245 ;
			RECT	13.571 50.181 13.603 50.245 ;
			RECT	13.739 50.181 13.771 50.245 ;
			RECT	13.907 50.181 13.939 50.245 ;
			RECT	14.075 50.181 14.107 50.245 ;
			RECT	14.243 50.181 14.275 50.245 ;
			RECT	14.411 50.181 14.443 50.245 ;
			RECT	14.579 50.181 14.611 50.245 ;
			RECT	14.747 50.181 14.779 50.245 ;
			RECT	14.915 50.181 14.947 50.245 ;
			RECT	15.083 50.181 15.115 50.245 ;
			RECT	15.251 50.181 15.283 50.245 ;
			RECT	15.419 50.181 15.451 50.245 ;
			RECT	15.587 50.181 15.619 50.245 ;
			RECT	15.755 50.181 15.787 50.245 ;
			RECT	15.923 50.181 15.955 50.245 ;
			RECT	16.091 50.181 16.123 50.245 ;
			RECT	16.259 50.181 16.291 50.245 ;
			RECT	16.427 50.181 16.459 50.245 ;
			RECT	16.595 50.181 16.627 50.245 ;
			RECT	16.763 50.181 16.795 50.245 ;
			RECT	16.931 50.181 16.963 50.245 ;
			RECT	17.099 50.181 17.131 50.245 ;
			RECT	17.267 50.181 17.299 50.245 ;
			RECT	17.435 50.181 17.467 50.245 ;
			RECT	17.603 50.181 17.635 50.245 ;
			RECT	17.771 50.181 17.803 50.245 ;
			RECT	17.939 50.181 17.971 50.245 ;
			RECT	18.107 50.181 18.139 50.245 ;
			RECT	18.275 50.181 18.307 50.245 ;
			RECT	18.443 50.181 18.475 50.245 ;
			RECT	18.611 50.181 18.643 50.245 ;
			RECT	18.779 50.181 18.811 50.245 ;
			RECT	18.947 50.181 18.979 50.245 ;
			RECT	19.115 50.181 19.147 50.245 ;
			RECT	19.283 50.181 19.315 50.245 ;
			RECT	19.451 50.181 19.483 50.245 ;
			RECT	19.619 50.181 19.651 50.245 ;
			RECT	19.787 50.181 19.819 50.245 ;
			RECT	19.955 50.181 19.987 50.245 ;
			RECT	20.123 50.181 20.155 50.245 ;
			RECT	20.291 50.181 20.323 50.245 ;
			RECT	20.459 50.181 20.491 50.245 ;
			RECT	20.627 50.181 20.659 50.245 ;
			RECT	20.795 50.181 20.827 50.245 ;
			RECT	20.963 50.181 20.995 50.245 ;
			RECT	21.131 50.181 21.163 50.245 ;
			RECT	21.299 50.181 21.331 50.245 ;
			RECT	21.467 50.181 21.499 50.245 ;
			RECT	21.635 50.181 21.667 50.245 ;
			RECT	21.803 50.181 21.835 50.245 ;
			RECT	21.971 50.181 22.003 50.245 ;
			RECT	22.139 50.181 22.171 50.245 ;
			RECT	22.307 50.181 22.339 50.245 ;
			RECT	22.475 50.181 22.507 50.245 ;
			RECT	22.643 50.181 22.675 50.245 ;
			RECT	22.811 50.181 22.843 50.245 ;
			RECT	22.979 50.181 23.011 50.245 ;
			RECT	23.147 50.181 23.179 50.245 ;
			RECT	23.315 50.181 23.347 50.245 ;
			RECT	23.483 50.181 23.515 50.245 ;
			RECT	23.651 50.181 23.683 50.245 ;
			RECT	23.819 50.181 23.851 50.245 ;
			RECT	23.987 50.181 24.019 50.245 ;
			RECT	24.155 50.181 24.187 50.245 ;
			RECT	24.323 50.181 24.355 50.245 ;
			RECT	24.491 50.181 24.523 50.245 ;
			RECT	24.659 50.181 24.691 50.245 ;
			RECT	24.827 50.181 24.859 50.245 ;
			RECT	24.995 50.181 25.027 50.245 ;
			RECT	25.163 50.181 25.195 50.245 ;
			RECT	25.331 50.181 25.363 50.245 ;
			RECT	25.499 50.181 25.531 50.245 ;
			RECT	25.667 50.181 25.699 50.245 ;
			RECT	25.835 50.181 25.867 50.245 ;
			RECT	26.003 50.181 26.035 50.245 ;
			RECT	26.171 50.181 26.203 50.245 ;
			RECT	26.339 50.181 26.371 50.245 ;
			RECT	26.507 50.181 26.539 50.245 ;
			RECT	26.675 50.181 26.707 50.245 ;
			RECT	26.843 50.181 26.875 50.245 ;
			RECT	27.011 50.181 27.043 50.245 ;
			RECT	27.179 50.181 27.211 50.245 ;
			RECT	27.347 50.181 27.379 50.245 ;
			RECT	27.515 50.181 27.547 50.245 ;
			RECT	27.683 50.181 27.715 50.245 ;
			RECT	27.851 50.181 27.883 50.245 ;
			RECT	28.019 50.181 28.051 50.245 ;
			RECT	28.187 50.181 28.219 50.245 ;
			RECT	28.355 50.181 28.387 50.245 ;
			RECT	28.523 50.181 28.555 50.245 ;
			RECT	28.691 50.181 28.723 50.245 ;
			RECT	28.859 50.181 28.891 50.245 ;
			RECT	29.027 50.181 29.059 50.245 ;
			RECT	29.195 50.181 29.227 50.245 ;
			RECT	29.363 50.181 29.395 50.245 ;
			RECT	29.531 50.181 29.563 50.245 ;
			RECT	29.699 50.181 29.731 50.245 ;
			RECT	29.867 50.181 29.899 50.245 ;
			RECT	30.035 50.181 30.067 50.245 ;
			RECT	30.203 50.181 30.235 50.245 ;
			RECT	30.371 50.181 30.403 50.245 ;
			RECT	30.539 50.181 30.571 50.245 ;
			RECT	30.707 50.181 30.739 50.245 ;
			RECT	30.875 50.181 30.907 50.245 ;
			RECT	31.043 50.181 31.075 50.245 ;
			RECT	31.211 50.181 31.243 50.245 ;
			RECT	31.379 50.181 31.411 50.245 ;
			RECT	31.547 50.181 31.579 50.245 ;
			RECT	31.715 50.181 31.747 50.245 ;
			RECT	31.883 50.181 31.915 50.245 ;
			RECT	32.051 50.181 32.083 50.245 ;
			RECT	32.219 50.181 32.251 50.245 ;
			RECT	32.387 50.181 32.419 50.245 ;
			RECT	32.555 50.181 32.587 50.245 ;
			RECT	32.723 50.181 32.755 50.245 ;
			RECT	32.891 50.181 32.923 50.245 ;
			RECT	33.059 50.181 33.091 50.245 ;
			RECT	33.227 50.181 33.259 50.245 ;
			RECT	33.395 50.181 33.427 50.245 ;
			RECT	33.563 50.181 33.595 50.245 ;
			RECT	33.731 50.181 33.763 50.245 ;
			RECT	33.899 50.181 33.931 50.245 ;
			RECT	34.067 50.181 34.099 50.245 ;
			RECT	34.235 50.181 34.267 50.245 ;
			RECT	34.403 50.181 34.435 50.245 ;
			RECT	34.571 50.181 34.603 50.245 ;
			RECT	34.739 50.181 34.771 50.245 ;
			RECT	34.907 50.181 34.939 50.245 ;
			RECT	35.075 50.181 35.107 50.245 ;
			RECT	35.243 50.181 35.275 50.245 ;
			RECT	35.411 50.181 35.443 50.245 ;
			RECT	35.579 50.181 35.611 50.245 ;
			RECT	35.747 50.181 35.779 50.245 ;
			RECT	35.915 50.181 35.947 50.245 ;
			RECT	36.083 50.181 36.115 50.245 ;
			RECT	36.251 50.181 36.283 50.245 ;
			RECT	36.419 50.181 36.451 50.245 ;
			RECT	36.587 50.181 36.619 50.245 ;
			RECT	36.755 50.181 36.787 50.245 ;
			RECT	36.923 50.181 36.955 50.245 ;
			RECT	37.091 50.181 37.123 50.245 ;
			RECT	37.259 50.181 37.291 50.245 ;
			RECT	37.427 50.181 37.459 50.245 ;
			RECT	37.595 50.181 37.627 50.245 ;
			RECT	37.763 50.181 37.795 50.245 ;
			RECT	37.931 50.181 37.963 50.245 ;
			RECT	38.099 50.181 38.131 50.245 ;
			RECT	38.267 50.181 38.299 50.245 ;
			RECT	38.435 50.181 38.467 50.245 ;
			RECT	38.603 50.181 38.635 50.245 ;
			RECT	38.771 50.181 38.803 50.245 ;
			RECT	38.939 50.181 38.971 50.245 ;
			RECT	39.107 50.181 39.139 50.245 ;
			RECT	39.275 50.181 39.307 50.245 ;
			RECT	39.443 50.181 39.475 50.245 ;
			RECT	39.611 50.181 39.643 50.245 ;
			RECT	39.779 50.181 39.811 50.245 ;
			RECT	39.947 50.181 39.979 50.245 ;
			RECT	40.115 50.181 40.147 50.245 ;
			RECT	40.283 50.181 40.315 50.245 ;
			RECT	40.451 50.181 40.483 50.245 ;
			RECT	40.619 50.181 40.651 50.245 ;
			RECT	40.787 50.181 40.819 50.245 ;
			RECT	40.955 50.181 40.987 50.245 ;
			RECT	41.123 50.181 41.155 50.245 ;
			RECT	41.291 50.181 41.323 50.245 ;
			RECT	41.459 50.181 41.491 50.245 ;
			RECT	41.627 50.181 41.659 50.245 ;
			RECT	41.795 50.181 41.827 50.245 ;
			RECT	41.963 50.181 41.995 50.245 ;
			RECT	42.131 50.181 42.163 50.245 ;
			RECT	42.299 50.181 42.331 50.245 ;
			RECT	42.467 50.181 42.499 50.245 ;
			RECT	42.635 50.181 42.667 50.245 ;
			RECT	42.803 50.181 42.835 50.245 ;
			RECT	42.971 50.181 43.003 50.245 ;
			RECT	43.139 50.181 43.171 50.245 ;
			RECT	43.307 50.181 43.339 50.245 ;
			RECT	43.475 50.181 43.507 50.245 ;
			RECT	43.643 50.181 43.675 50.245 ;
			RECT	43.811 50.181 43.843 50.245 ;
			RECT	43.979 50.181 44.011 50.245 ;
			RECT	44.147 50.181 44.179 50.245 ;
			RECT	44.315 50.181 44.347 50.245 ;
			RECT	44.483 50.181 44.515 50.245 ;
			RECT	44.651 50.181 44.683 50.245 ;
			RECT	44.819 50.181 44.851 50.245 ;
			RECT	44.987 50.181 45.019 50.245 ;
			RECT	45.155 50.181 45.187 50.245 ;
			RECT	45.323 50.181 45.355 50.245 ;
			RECT	45.491 50.181 45.523 50.245 ;
			RECT	45.659 50.181 45.691 50.245 ;
			RECT	45.827 50.181 45.859 50.245 ;
			RECT	45.995 50.181 46.027 50.245 ;
			RECT	46.163 50.181 46.195 50.245 ;
			RECT	46.331 50.181 46.363 50.245 ;
			RECT	46.499 50.181 46.531 50.245 ;
			RECT	46.667 50.181 46.699 50.245 ;
			RECT	46.835 50.181 46.867 50.245 ;
			RECT	47.003 50.181 47.035 50.245 ;
			RECT	47.171 50.181 47.203 50.245 ;
			RECT	47.339 50.181 47.371 50.245 ;
			RECT	47.507 50.181 47.539 50.245 ;
			RECT	47.675 50.181 47.707 50.245 ;
			RECT	47.843 50.181 47.875 50.245 ;
			RECT	48.011 50.181 48.043 50.245 ;
			RECT	48.179 50.181 48.211 50.245 ;
			RECT	48.347 50.181 48.379 50.245 ;
			RECT	48.515 50.181 48.547 50.245 ;
			RECT	48.683 50.181 48.715 50.245 ;
			RECT	48.851 50.181 48.883 50.245 ;
			RECT	49.019 50.181 49.051 50.245 ;
			RECT	49.187 50.181 49.219 50.245 ;
			RECT	49.439 50.181 49.471 50.245 ;
			RECT	52.944 50.181 52.976 50.245 ;
			RECT	53.91 50.181 53.942 50.245 ;
			RECT	54.812 50.181 54.844 50.245 ;
			RECT	55.969 50.181 56.033 50.245 ;
			RECT	58.733 50.181 58.765 50.245 ;
			RECT	58.985 50.181 59.017 50.245 ;
			RECT	59.153 50.181 59.185 50.245 ;
			RECT	59.321 50.181 59.353 50.245 ;
			RECT	59.489 50.181 59.521 50.245 ;
			RECT	59.657 50.181 59.689 50.245 ;
			RECT	59.825 50.181 59.857 50.245 ;
			RECT	59.993 50.181 60.025 50.245 ;
			RECT	60.161 50.181 60.193 50.245 ;
			RECT	60.329 50.181 60.361 50.245 ;
			RECT	60.497 50.181 60.529 50.245 ;
			RECT	60.665 50.181 60.697 50.245 ;
			RECT	60.833 50.181 60.865 50.245 ;
			RECT	61.001 50.181 61.033 50.245 ;
			RECT	61.169 50.181 61.201 50.245 ;
			RECT	61.337 50.181 61.369 50.245 ;
			RECT	61.505 50.181 61.537 50.245 ;
			RECT	61.673 50.181 61.705 50.245 ;
			RECT	61.841 50.181 61.873 50.245 ;
			RECT	62.009 50.181 62.041 50.245 ;
			RECT	62.177 50.181 62.209 50.245 ;
			RECT	62.345 50.181 62.377 50.245 ;
			RECT	62.513 50.181 62.545 50.245 ;
			RECT	62.681 50.181 62.713 50.245 ;
			RECT	62.849 50.181 62.881 50.245 ;
			RECT	63.017 50.181 63.049 50.245 ;
			RECT	63.185 50.181 63.217 50.245 ;
			RECT	63.353 50.181 63.385 50.245 ;
			RECT	63.521 50.181 63.553 50.245 ;
			RECT	63.689 50.181 63.721 50.245 ;
			RECT	63.857 50.181 63.889 50.245 ;
			RECT	64.025 50.181 64.057 50.245 ;
			RECT	64.193 50.181 64.225 50.245 ;
			RECT	64.361 50.181 64.393 50.245 ;
			RECT	64.529 50.181 64.561 50.245 ;
			RECT	64.697 50.181 64.729 50.245 ;
			RECT	64.865 50.181 64.897 50.245 ;
			RECT	65.033 50.181 65.065 50.245 ;
			RECT	65.201 50.181 65.233 50.245 ;
			RECT	65.369 50.181 65.401 50.245 ;
			RECT	65.537 50.181 65.569 50.245 ;
			RECT	65.705 50.181 65.737 50.245 ;
			RECT	65.873 50.181 65.905 50.245 ;
			RECT	66.041 50.181 66.073 50.245 ;
			RECT	66.209 50.181 66.241 50.245 ;
			RECT	66.377 50.181 66.409 50.245 ;
			RECT	66.545 50.181 66.577 50.245 ;
			RECT	66.713 50.181 66.745 50.245 ;
			RECT	66.881 50.181 66.913 50.245 ;
			RECT	67.049 50.181 67.081 50.245 ;
			RECT	67.217 50.181 67.249 50.245 ;
			RECT	67.385 50.181 67.417 50.245 ;
			RECT	67.553 50.181 67.585 50.245 ;
			RECT	67.721 50.181 67.753 50.245 ;
			RECT	67.889 50.181 67.921 50.245 ;
			RECT	68.057 50.181 68.089 50.245 ;
			RECT	68.225 50.181 68.257 50.245 ;
			RECT	68.393 50.181 68.425 50.245 ;
			RECT	68.561 50.181 68.593 50.245 ;
			RECT	68.729 50.181 68.761 50.245 ;
			RECT	68.897 50.181 68.929 50.245 ;
			RECT	69.065 50.181 69.097 50.245 ;
			RECT	69.233 50.181 69.265 50.245 ;
			RECT	69.401 50.181 69.433 50.245 ;
			RECT	69.569 50.181 69.601 50.245 ;
			RECT	69.737 50.181 69.769 50.245 ;
			RECT	69.905 50.181 69.937 50.245 ;
			RECT	70.073 50.181 70.105 50.245 ;
			RECT	70.241 50.181 70.273 50.245 ;
			RECT	70.409 50.181 70.441 50.245 ;
			RECT	70.577 50.181 70.609 50.245 ;
			RECT	70.745 50.181 70.777 50.245 ;
			RECT	70.913 50.181 70.945 50.245 ;
			RECT	71.081 50.181 71.113 50.245 ;
			RECT	71.249 50.181 71.281 50.245 ;
			RECT	71.417 50.181 71.449 50.245 ;
			RECT	71.585 50.181 71.617 50.245 ;
			RECT	71.753 50.181 71.785 50.245 ;
			RECT	71.921 50.181 71.953 50.245 ;
			RECT	72.089 50.181 72.121 50.245 ;
			RECT	72.257 50.181 72.289 50.245 ;
			RECT	72.425 50.181 72.457 50.245 ;
			RECT	72.593 50.181 72.625 50.245 ;
			RECT	72.761 50.181 72.793 50.245 ;
			RECT	72.929 50.181 72.961 50.245 ;
			RECT	73.097 50.181 73.129 50.245 ;
			RECT	73.265 50.181 73.297 50.245 ;
			RECT	73.433 50.181 73.465 50.245 ;
			RECT	73.601 50.181 73.633 50.245 ;
			RECT	73.769 50.181 73.801 50.245 ;
			RECT	73.937 50.181 73.969 50.245 ;
			RECT	74.105 50.181 74.137 50.245 ;
			RECT	74.273 50.181 74.305 50.245 ;
			RECT	74.441 50.181 74.473 50.245 ;
			RECT	74.609 50.181 74.641 50.245 ;
			RECT	74.777 50.181 74.809 50.245 ;
			RECT	74.945 50.181 74.977 50.245 ;
			RECT	75.113 50.181 75.145 50.245 ;
			RECT	75.281 50.181 75.313 50.245 ;
			RECT	75.449 50.181 75.481 50.245 ;
			RECT	75.617 50.181 75.649 50.245 ;
			RECT	75.785 50.181 75.817 50.245 ;
			RECT	75.953 50.181 75.985 50.245 ;
			RECT	76.121 50.181 76.153 50.245 ;
			RECT	76.289 50.181 76.321 50.245 ;
			RECT	76.457 50.181 76.489 50.245 ;
			RECT	76.625 50.181 76.657 50.245 ;
			RECT	76.793 50.181 76.825 50.245 ;
			RECT	76.961 50.181 76.993 50.245 ;
			RECT	77.129 50.181 77.161 50.245 ;
			RECT	77.297 50.181 77.329 50.245 ;
			RECT	77.465 50.181 77.497 50.245 ;
			RECT	77.633 50.181 77.665 50.245 ;
			RECT	77.801 50.181 77.833 50.245 ;
			RECT	77.969 50.181 78.001 50.245 ;
			RECT	78.137 50.181 78.169 50.245 ;
			RECT	78.305 50.181 78.337 50.245 ;
			RECT	78.473 50.181 78.505 50.245 ;
			RECT	78.641 50.181 78.673 50.245 ;
			RECT	78.809 50.181 78.841 50.245 ;
			RECT	78.977 50.181 79.009 50.245 ;
			RECT	79.145 50.181 79.177 50.245 ;
			RECT	79.313 50.181 79.345 50.245 ;
			RECT	79.481 50.181 79.513 50.245 ;
			RECT	79.649 50.181 79.681 50.245 ;
			RECT	79.817 50.181 79.849 50.245 ;
			RECT	79.985 50.181 80.017 50.245 ;
			RECT	80.153 50.181 80.185 50.245 ;
			RECT	80.321 50.181 80.353 50.245 ;
			RECT	80.489 50.181 80.521 50.245 ;
			RECT	80.657 50.181 80.689 50.245 ;
			RECT	80.825 50.181 80.857 50.245 ;
			RECT	80.993 50.181 81.025 50.245 ;
			RECT	81.161 50.181 81.193 50.245 ;
			RECT	81.329 50.181 81.361 50.245 ;
			RECT	81.497 50.181 81.529 50.245 ;
			RECT	81.665 50.181 81.697 50.245 ;
			RECT	81.833 50.181 81.865 50.245 ;
			RECT	82.001 50.181 82.033 50.245 ;
			RECT	82.169 50.181 82.201 50.245 ;
			RECT	82.337 50.181 82.369 50.245 ;
			RECT	82.505 50.181 82.537 50.245 ;
			RECT	82.673 50.181 82.705 50.245 ;
			RECT	82.841 50.181 82.873 50.245 ;
			RECT	83.009 50.181 83.041 50.245 ;
			RECT	83.177 50.181 83.209 50.245 ;
			RECT	83.345 50.181 83.377 50.245 ;
			RECT	83.513 50.181 83.545 50.245 ;
			RECT	83.681 50.181 83.713 50.245 ;
			RECT	83.849 50.181 83.881 50.245 ;
			RECT	84.017 50.181 84.049 50.245 ;
			RECT	84.185 50.181 84.217 50.245 ;
			RECT	84.353 50.181 84.385 50.245 ;
			RECT	84.521 50.181 84.553 50.245 ;
			RECT	84.689 50.181 84.721 50.245 ;
			RECT	84.857 50.181 84.889 50.245 ;
			RECT	85.025 50.181 85.057 50.245 ;
			RECT	85.193 50.181 85.225 50.245 ;
			RECT	85.361 50.181 85.393 50.245 ;
			RECT	85.529 50.181 85.561 50.245 ;
			RECT	85.697 50.181 85.729 50.245 ;
			RECT	85.865 50.181 85.897 50.245 ;
			RECT	86.033 50.181 86.065 50.245 ;
			RECT	86.201 50.181 86.233 50.245 ;
			RECT	86.369 50.181 86.401 50.245 ;
			RECT	86.537 50.181 86.569 50.245 ;
			RECT	86.705 50.181 86.737 50.245 ;
			RECT	86.873 50.181 86.905 50.245 ;
			RECT	87.041 50.181 87.073 50.245 ;
			RECT	87.209 50.181 87.241 50.245 ;
			RECT	87.377 50.181 87.409 50.245 ;
			RECT	87.545 50.181 87.577 50.245 ;
			RECT	87.713 50.181 87.745 50.245 ;
			RECT	87.881 50.181 87.913 50.245 ;
			RECT	88.049 50.181 88.081 50.245 ;
			RECT	88.217 50.181 88.249 50.245 ;
			RECT	88.385 50.181 88.417 50.245 ;
			RECT	88.553 50.181 88.585 50.245 ;
			RECT	88.721 50.181 88.753 50.245 ;
			RECT	88.889 50.181 88.921 50.245 ;
			RECT	89.057 50.181 89.089 50.245 ;
			RECT	89.225 50.181 89.257 50.245 ;
			RECT	89.393 50.181 89.425 50.245 ;
			RECT	89.561 50.181 89.593 50.245 ;
			RECT	89.729 50.181 89.761 50.245 ;
			RECT	89.897 50.181 89.929 50.245 ;
			RECT	90.065 50.181 90.097 50.245 ;
			RECT	90.233 50.181 90.265 50.245 ;
			RECT	90.401 50.181 90.433 50.245 ;
			RECT	90.569 50.181 90.601 50.245 ;
			RECT	90.737 50.181 90.769 50.245 ;
			RECT	90.905 50.181 90.937 50.245 ;
			RECT	91.073 50.181 91.105 50.245 ;
			RECT	91.241 50.181 91.273 50.245 ;
			RECT	91.409 50.181 91.441 50.245 ;
			RECT	91.577 50.181 91.609 50.245 ;
			RECT	91.745 50.181 91.777 50.245 ;
			RECT	91.913 50.181 91.945 50.245 ;
			RECT	92.081 50.181 92.113 50.245 ;
			RECT	92.249 50.181 92.281 50.245 ;
			RECT	92.417 50.181 92.449 50.245 ;
			RECT	92.585 50.181 92.617 50.245 ;
			RECT	92.753 50.181 92.785 50.245 ;
			RECT	92.921 50.181 92.953 50.245 ;
			RECT	93.089 50.181 93.121 50.245 ;
			RECT	93.257 50.181 93.289 50.245 ;
			RECT	93.425 50.181 93.457 50.245 ;
			RECT	93.593 50.181 93.625 50.245 ;
			RECT	93.761 50.181 93.793 50.245 ;
			RECT	93.929 50.181 93.961 50.245 ;
			RECT	94.097 50.181 94.129 50.245 ;
			RECT	94.265 50.181 94.297 50.245 ;
			RECT	94.433 50.181 94.465 50.245 ;
			RECT	94.601 50.181 94.633 50.245 ;
			RECT	94.769 50.181 94.801 50.245 ;
			RECT	94.937 50.181 94.969 50.245 ;
			RECT	95.105 50.181 95.137 50.245 ;
			RECT	95.273 50.181 95.305 50.245 ;
			RECT	95.441 50.181 95.473 50.245 ;
			RECT	95.609 50.181 95.641 50.245 ;
			RECT	95.777 50.181 95.809 50.245 ;
			RECT	95.945 50.181 95.977 50.245 ;
			RECT	96.113 50.181 96.145 50.245 ;
			RECT	96.281 50.181 96.313 50.245 ;
			RECT	96.449 50.181 96.481 50.245 ;
			RECT	96.617 50.181 96.649 50.245 ;
			RECT	96.785 50.181 96.817 50.245 ;
			RECT	96.953 50.181 96.985 50.245 ;
			RECT	97.121 50.181 97.153 50.245 ;
			RECT	97.289 50.181 97.321 50.245 ;
			RECT	97.457 50.181 97.489 50.245 ;
			RECT	97.625 50.181 97.657 50.245 ;
			RECT	97.793 50.181 97.825 50.245 ;
			RECT	97.961 50.181 97.993 50.245 ;
			RECT	98.129 50.181 98.161 50.245 ;
			RECT	98.297 50.181 98.329 50.245 ;
			RECT	98.465 50.181 98.497 50.245 ;
			RECT	98.633 50.181 98.665 50.245 ;
			RECT	98.801 50.181 98.833 50.245 ;
			RECT	98.969 50.181 99.001 50.245 ;
			RECT	99.137 50.181 99.169 50.245 ;
			RECT	99.305 50.181 99.337 50.245 ;
			RECT	99.473 50.181 99.505 50.245 ;
			RECT	99.641 50.181 99.673 50.245 ;
			RECT	99.809 50.181 99.841 50.245 ;
			RECT	99.977 50.181 100.009 50.245 ;
			RECT	100.145 50.181 100.177 50.245 ;
			RECT	100.313 50.181 100.345 50.245 ;
			RECT	100.481 50.181 100.513 50.245 ;
			RECT	100.649 50.181 100.681 50.245 ;
			RECT	100.817 50.181 100.849 50.245 ;
			RECT	100.985 50.181 101.017 50.245 ;
			RECT	101.153 50.181 101.185 50.245 ;
			RECT	101.321 50.181 101.353 50.245 ;
			RECT	101.489 50.181 101.521 50.245 ;
			RECT	101.657 50.181 101.689 50.245 ;
			RECT	101.825 50.181 101.857 50.245 ;
			RECT	101.993 50.181 102.025 50.245 ;
			RECT	102.245 50.181 102.277 50.245 ;
			RECT	103.085 50.181 103.117 50.245 ;
			RECT	103.925 50.181 103.957 50.245 ;
			RECT	104.177 50.181 104.209 50.245 ;
			RECT	104.345 50.181 104.377 50.245 ;
			RECT	104.513 50.181 104.545 50.245 ;
			RECT	104.681 50.181 104.713 50.245 ;
			RECT	104.849 50.181 104.881 50.245 ;
			RECT	105.017 50.181 105.049 50.245 ;
			RECT	105.185 50.181 105.217 50.245 ;
			RECT	105.353 50.181 105.385 50.245 ;
			RECT	105.521 50.181 105.553 50.245 ;
			RECT	105.689 50.181 105.721 50.245 ;
			RECT	105.857 50.181 105.889 50.245 ;
			RECT	106.025 50.181 106.057 50.245 ;
			RECT	106.193 50.181 106.225 50.245 ;
			RECT	106.361 50.181 106.393 50.245 ;
			RECT	106.529 50.181 106.561 50.245 ;
			RECT	106.697 50.181 106.729 50.245 ;
			RECT	106.865 50.181 106.897 50.245 ;
			RECT	107.033 50.181 107.065 50.245 ;
			RECT	107.201 50.181 107.233 50.245 ;
			RECT	107.369 50.181 107.401 50.245 ;
			RECT	107.537 50.181 107.569 50.245 ;
			RECT	107.705 50.181 107.737 50.245 ;
			RECT	107.873 50.181 107.905 50.245 ;
			RECT	108.041 50.181 108.073 50.245 ;
			RECT	108.209 50.181 108.241 50.245 ;
			RECT	108.377 50.181 108.409 50.245 ;
			RECT	108.545 50.181 108.577 50.245 ;
			RECT	108.713 50.181 108.745 50.245 ;
			RECT	108.881 50.181 108.913 50.245 ;
			RECT	109.049 50.181 109.081 50.245 ;
			RECT	109.217 50.181 109.249 50.245 ;
			RECT	109.385 50.181 109.417 50.245 ;
			RECT	109.553 50.181 109.585 50.245 ;
			RECT	109.721 50.181 109.753 50.245 ;
			RECT	109.889 50.181 109.921 50.245 ;
			RECT	110.057 50.181 110.089 50.245 ;
			RECT	110.225 50.181 110.257 50.245 ;
			RECT	110.393 50.181 110.425 50.245 ;
			RECT	110.561 50.181 110.593 50.245 ;
			RECT	110.729 50.181 110.761 50.245 ;
			RECT	110.897 50.181 110.929 50.245 ;
			RECT	111.065 50.181 111.097 50.245 ;
			RECT	111.233 50.181 111.265 50.245 ;
			RECT	111.401 50.181 111.433 50.245 ;
			RECT	111.569 50.181 111.601 50.245 ;
			RECT	111.737 50.181 111.769 50.245 ;
			RECT	111.905 50.181 111.937 50.245 ;
			RECT	112.073 50.181 112.105 50.245 ;
			RECT	112.241 50.181 112.273 50.245 ;
			RECT	112.409 50.181 112.441 50.245 ;
			RECT	112.577 50.181 112.609 50.245 ;
			RECT	112.745 50.181 112.777 50.245 ;
			RECT	112.913 50.181 112.945 50.245 ;
			RECT	113.081 50.181 113.113 50.245 ;
			RECT	113.249 50.181 113.281 50.245 ;
			RECT	113.417 50.181 113.449 50.245 ;
			RECT	113.585 50.181 113.617 50.245 ;
			RECT	113.753 50.181 113.785 50.245 ;
			RECT	113.921 50.181 113.953 50.245 ;
			RECT	114.089 50.181 114.121 50.245 ;
			RECT	114.257 50.181 114.289 50.245 ;
			RECT	114.425 50.181 114.457 50.245 ;
			RECT	114.593 50.181 114.625 50.245 ;
			RECT	114.761 50.181 114.793 50.245 ;
			RECT	114.929 50.181 114.961 50.245 ;
			RECT	115.097 50.181 115.129 50.245 ;
			RECT	115.265 50.181 115.297 50.245 ;
			RECT	115.433 50.181 115.465 50.245 ;
			RECT	115.601 50.181 115.633 50.245 ;
			RECT	115.769 50.181 115.801 50.245 ;
			RECT	115.937 50.181 115.969 50.245 ;
			RECT	116.105 50.181 116.137 50.245 ;
			RECT	116.273 50.181 116.305 50.245 ;
			RECT	116.441 50.181 116.473 50.245 ;
			RECT	116.609 50.181 116.641 50.245 ;
			RECT	116.777 50.181 116.809 50.245 ;
			RECT	116.945 50.181 116.977 50.245 ;
			RECT	117.113 50.181 117.145 50.245 ;
			RECT	117.281 50.181 117.313 50.245 ;
			RECT	117.449 50.181 117.481 50.245 ;
			RECT	117.617 50.181 117.649 50.245 ;
			RECT	117.785 50.181 117.817 50.245 ;
			RECT	117.953 50.181 117.985 50.245 ;
			RECT	118.121 50.181 118.153 50.245 ;
			RECT	118.289 50.181 118.321 50.245 ;
			RECT	118.457 50.181 118.489 50.245 ;
			RECT	118.625 50.181 118.657 50.245 ;
			RECT	118.793 50.181 118.825 50.245 ;
			RECT	118.961 50.181 118.993 50.245 ;
			RECT	119.129 50.181 119.161 50.245 ;
			RECT	119.297 50.181 119.329 50.245 ;
			RECT	119.465 50.181 119.497 50.245 ;
			RECT	119.633 50.181 119.665 50.245 ;
			RECT	119.801 50.181 119.833 50.245 ;
			RECT	119.969 50.181 120.001 50.245 ;
			RECT	120.137 50.181 120.169 50.245 ;
			RECT	120.305 50.181 120.337 50.245 ;
			RECT	120.473 50.181 120.505 50.245 ;
			RECT	120.641 50.181 120.673 50.245 ;
			RECT	120.809 50.181 120.841 50.245 ;
			RECT	120.977 50.181 121.009 50.245 ;
			RECT	121.145 50.181 121.177 50.245 ;
			RECT	121.313 50.181 121.345 50.245 ;
			RECT	121.481 50.181 121.513 50.245 ;
			RECT	121.649 50.181 121.681 50.245 ;
			RECT	121.817 50.181 121.849 50.245 ;
			RECT	121.985 50.181 122.017 50.245 ;
			RECT	122.153 50.181 122.185 50.245 ;
			RECT	122.321 50.181 122.353 50.245 ;
			RECT	122.489 50.181 122.521 50.245 ;
			RECT	122.657 50.181 122.689 50.245 ;
			RECT	122.825 50.181 122.857 50.245 ;
			RECT	122.993 50.181 123.025 50.245 ;
			RECT	123.161 50.181 123.193 50.245 ;
			RECT	123.329 50.181 123.361 50.245 ;
			RECT	123.497 50.181 123.529 50.245 ;
			RECT	123.665 50.181 123.697 50.245 ;
			RECT	123.833 50.181 123.865 50.245 ;
			RECT	124.001 50.181 124.033 50.245 ;
			RECT	124.169 50.181 124.201 50.245 ;
			RECT	124.337 50.181 124.369 50.245 ;
			RECT	124.505 50.181 124.537 50.245 ;
			RECT	124.673 50.181 124.705 50.245 ;
			RECT	124.841 50.181 124.873 50.245 ;
			RECT	125.009 50.181 125.041 50.245 ;
			RECT	125.177 50.181 125.209 50.245 ;
			RECT	125.345 50.181 125.377 50.245 ;
			RECT	125.513 50.181 125.545 50.245 ;
			RECT	125.681 50.181 125.713 50.245 ;
			RECT	125.849 50.181 125.881 50.245 ;
			RECT	126.017 50.181 126.049 50.245 ;
			RECT	126.185 50.181 126.217 50.245 ;
			RECT	126.353 50.181 126.385 50.245 ;
			RECT	126.521 50.181 126.553 50.245 ;
			RECT	126.689 50.181 126.721 50.245 ;
			RECT	126.857 50.181 126.889 50.245 ;
			RECT	127.025 50.181 127.057 50.245 ;
			RECT	127.193 50.181 127.225 50.245 ;
			RECT	127.361 50.181 127.393 50.245 ;
			RECT	127.529 50.181 127.561 50.245 ;
			RECT	127.697 50.181 127.729 50.245 ;
			RECT	127.865 50.181 127.897 50.245 ;
			RECT	128.033 50.181 128.065 50.245 ;
			RECT	128.201 50.181 128.233 50.245 ;
			RECT	128.369 50.181 128.401 50.245 ;
			RECT	128.537 50.181 128.569 50.245 ;
			RECT	128.705 50.181 128.737 50.245 ;
			RECT	128.873 50.181 128.905 50.245 ;
			RECT	129.041 50.181 129.073 50.245 ;
			RECT	129.209 50.181 129.241 50.245 ;
			RECT	129.377 50.181 129.409 50.245 ;
			RECT	129.545 50.181 129.577 50.245 ;
			RECT	129.713 50.181 129.745 50.245 ;
			RECT	129.881 50.181 129.913 50.245 ;
			RECT	130.049 50.181 130.081 50.245 ;
			RECT	130.217 50.181 130.249 50.245 ;
			RECT	130.385 50.181 130.417 50.245 ;
			RECT	130.553 50.181 130.585 50.245 ;
			RECT	130.721 50.181 130.753 50.245 ;
			RECT	130.889 50.181 130.921 50.245 ;
			RECT	131.057 50.181 131.089 50.245 ;
			RECT	131.225 50.181 131.257 50.245 ;
			RECT	131.393 50.181 131.425 50.245 ;
			RECT	131.561 50.181 131.593 50.245 ;
			RECT	131.729 50.181 131.761 50.245 ;
			RECT	131.897 50.181 131.929 50.245 ;
			RECT	132.065 50.181 132.097 50.245 ;
			RECT	132.233 50.181 132.265 50.245 ;
			RECT	132.401 50.181 132.433 50.245 ;
			RECT	132.569 50.181 132.601 50.245 ;
			RECT	132.737 50.181 132.769 50.245 ;
			RECT	132.905 50.181 132.937 50.245 ;
			RECT	133.073 50.181 133.105 50.245 ;
			RECT	133.241 50.181 133.273 50.245 ;
			RECT	133.409 50.181 133.441 50.245 ;
			RECT	133.577 50.181 133.609 50.245 ;
			RECT	133.745 50.181 133.777 50.245 ;
			RECT	133.913 50.181 133.945 50.245 ;
			RECT	134.081 50.181 134.113 50.245 ;
			RECT	134.249 50.181 134.281 50.245 ;
			RECT	134.417 50.181 134.449 50.245 ;
			RECT	134.585 50.181 134.617 50.245 ;
			RECT	134.753 50.181 134.785 50.245 ;
			RECT	134.921 50.181 134.953 50.245 ;
			RECT	135.089 50.181 135.121 50.245 ;
			RECT	135.257 50.181 135.289 50.245 ;
			RECT	135.425 50.181 135.457 50.245 ;
			RECT	135.593 50.181 135.625 50.245 ;
			RECT	135.761 50.181 135.793 50.245 ;
			RECT	135.929 50.181 135.961 50.245 ;
			RECT	136.097 50.181 136.129 50.245 ;
			RECT	136.265 50.181 136.297 50.245 ;
			RECT	136.433 50.181 136.465 50.245 ;
			RECT	136.601 50.181 136.633 50.245 ;
			RECT	136.769 50.181 136.801 50.245 ;
			RECT	136.937 50.181 136.969 50.245 ;
			RECT	137.105 50.181 137.137 50.245 ;
			RECT	137.273 50.181 137.305 50.245 ;
			RECT	137.441 50.181 137.473 50.245 ;
			RECT	137.609 50.181 137.641 50.245 ;
			RECT	137.777 50.181 137.809 50.245 ;
			RECT	137.945 50.181 137.977 50.245 ;
			RECT	138.113 50.181 138.145 50.245 ;
			RECT	138.281 50.181 138.313 50.245 ;
			RECT	138.449 50.181 138.481 50.245 ;
			RECT	138.617 50.181 138.649 50.245 ;
			RECT	138.785 50.181 138.817 50.245 ;
			RECT	138.953 50.181 138.985 50.245 ;
			RECT	139.121 50.181 139.153 50.245 ;
			RECT	139.289 50.181 139.321 50.245 ;
			RECT	139.457 50.181 139.489 50.245 ;
			RECT	139.625 50.181 139.657 50.245 ;
			RECT	139.793 50.181 139.825 50.245 ;
			RECT	139.961 50.181 139.993 50.245 ;
			RECT	140.129 50.181 140.161 50.245 ;
			RECT	140.297 50.181 140.329 50.245 ;
			RECT	140.465 50.181 140.497 50.245 ;
			RECT	140.633 50.181 140.665 50.245 ;
			RECT	140.801 50.181 140.833 50.245 ;
			RECT	140.969 50.181 141.001 50.245 ;
			RECT	141.137 50.181 141.169 50.245 ;
			RECT	141.305 50.181 141.337 50.245 ;
			RECT	141.473 50.181 141.505 50.245 ;
			RECT	141.641 50.181 141.673 50.245 ;
			RECT	141.809 50.181 141.841 50.245 ;
			RECT	141.977 50.181 142.009 50.245 ;
			RECT	142.145 50.181 142.177 50.245 ;
			RECT	142.313 50.181 142.345 50.245 ;
			RECT	142.481 50.181 142.513 50.245 ;
			RECT	142.649 50.181 142.681 50.245 ;
			RECT	142.817 50.181 142.849 50.245 ;
			RECT	142.985 50.181 143.017 50.245 ;
			RECT	143.153 50.181 143.185 50.245 ;
			RECT	143.321 50.181 143.353 50.245 ;
			RECT	143.489 50.181 143.521 50.245 ;
			RECT	143.657 50.181 143.689 50.245 ;
			RECT	143.825 50.181 143.857 50.245 ;
			RECT	143.993 50.181 144.025 50.245 ;
			RECT	144.161 50.181 144.193 50.245 ;
			RECT	144.329 50.181 144.361 50.245 ;
			RECT	144.497 50.181 144.529 50.245 ;
			RECT	144.665 50.181 144.697 50.245 ;
			RECT	144.833 50.181 144.865 50.245 ;
			RECT	145.001 50.181 145.033 50.245 ;
			RECT	145.169 50.181 145.201 50.245 ;
			RECT	145.337 50.181 145.369 50.245 ;
			RECT	145.505 50.181 145.537 50.245 ;
			RECT	145.673 50.181 145.705 50.245 ;
			RECT	145.841 50.181 145.873 50.245 ;
			RECT	146.009 50.181 146.041 50.245 ;
			RECT	146.177 50.181 146.209 50.245 ;
			RECT	146.345 50.181 146.377 50.245 ;
			RECT	146.513 50.181 146.545 50.245 ;
			RECT	146.681 50.181 146.713 50.245 ;
			RECT	146.849 50.181 146.881 50.245 ;
			RECT	147.017 50.181 147.049 50.245 ;
			RECT	147.185 50.181 147.217 50.245 ;
			RECT	147.437 50.181 147.469 50.245 ;
			RECT	150.942 50.181 150.974 50.245 ;
			RECT	151.908 50.181 151.94 50.245 ;
			RECT	152.81 50.181 152.842 50.245 ;
			RECT	153.967 50.181 154.031 50.245 ;
			RECT	156.731 50.181 156.763 50.245 ;
			RECT	156.983 50.181 157.015 50.245 ;
			RECT	157.151 50.181 157.183 50.245 ;
			RECT	157.319 50.181 157.351 50.245 ;
			RECT	157.487 50.181 157.519 50.245 ;
			RECT	157.655 50.181 157.687 50.245 ;
			RECT	157.823 50.181 157.855 50.245 ;
			RECT	157.991 50.181 158.023 50.245 ;
			RECT	158.159 50.181 158.191 50.245 ;
			RECT	158.327 50.181 158.359 50.245 ;
			RECT	158.495 50.181 158.527 50.245 ;
			RECT	158.663 50.181 158.695 50.245 ;
			RECT	158.831 50.181 158.863 50.245 ;
			RECT	158.999 50.181 159.031 50.245 ;
			RECT	159.167 50.181 159.199 50.245 ;
			RECT	159.335 50.181 159.367 50.245 ;
			RECT	159.503 50.181 159.535 50.245 ;
			RECT	159.671 50.181 159.703 50.245 ;
			RECT	159.839 50.181 159.871 50.245 ;
			RECT	160.007 50.181 160.039 50.245 ;
			RECT	160.175 50.181 160.207 50.245 ;
			RECT	160.343 50.181 160.375 50.245 ;
			RECT	160.511 50.181 160.543 50.245 ;
			RECT	160.679 50.181 160.711 50.245 ;
			RECT	160.847 50.181 160.879 50.245 ;
			RECT	161.015 50.181 161.047 50.245 ;
			RECT	161.183 50.181 161.215 50.245 ;
			RECT	161.351 50.181 161.383 50.245 ;
			RECT	161.519 50.181 161.551 50.245 ;
			RECT	161.687 50.181 161.719 50.245 ;
			RECT	161.855 50.181 161.887 50.245 ;
			RECT	162.023 50.181 162.055 50.245 ;
			RECT	162.191 50.181 162.223 50.245 ;
			RECT	162.359 50.181 162.391 50.245 ;
			RECT	162.527 50.181 162.559 50.245 ;
			RECT	162.695 50.181 162.727 50.245 ;
			RECT	162.863 50.181 162.895 50.245 ;
			RECT	163.031 50.181 163.063 50.245 ;
			RECT	163.199 50.181 163.231 50.245 ;
			RECT	163.367 50.181 163.399 50.245 ;
			RECT	163.535 50.181 163.567 50.245 ;
			RECT	163.703 50.181 163.735 50.245 ;
			RECT	163.871 50.181 163.903 50.245 ;
			RECT	164.039 50.181 164.071 50.245 ;
			RECT	164.207 50.181 164.239 50.245 ;
			RECT	164.375 50.181 164.407 50.245 ;
			RECT	164.543 50.181 164.575 50.245 ;
			RECT	164.711 50.181 164.743 50.245 ;
			RECT	164.879 50.181 164.911 50.245 ;
			RECT	165.047 50.181 165.079 50.245 ;
			RECT	165.215 50.181 165.247 50.245 ;
			RECT	165.383 50.181 165.415 50.245 ;
			RECT	165.551 50.181 165.583 50.245 ;
			RECT	165.719 50.181 165.751 50.245 ;
			RECT	165.887 50.181 165.919 50.245 ;
			RECT	166.055 50.181 166.087 50.245 ;
			RECT	166.223 50.181 166.255 50.245 ;
			RECT	166.391 50.181 166.423 50.245 ;
			RECT	166.559 50.181 166.591 50.245 ;
			RECT	166.727 50.181 166.759 50.245 ;
			RECT	166.895 50.181 166.927 50.245 ;
			RECT	167.063 50.181 167.095 50.245 ;
			RECT	167.231 50.181 167.263 50.245 ;
			RECT	167.399 50.181 167.431 50.245 ;
			RECT	167.567 50.181 167.599 50.245 ;
			RECT	167.735 50.181 167.767 50.245 ;
			RECT	167.903 50.181 167.935 50.245 ;
			RECT	168.071 50.181 168.103 50.245 ;
			RECT	168.239 50.181 168.271 50.245 ;
			RECT	168.407 50.181 168.439 50.245 ;
			RECT	168.575 50.181 168.607 50.245 ;
			RECT	168.743 50.181 168.775 50.245 ;
			RECT	168.911 50.181 168.943 50.245 ;
			RECT	169.079 50.181 169.111 50.245 ;
			RECT	169.247 50.181 169.279 50.245 ;
			RECT	169.415 50.181 169.447 50.245 ;
			RECT	169.583 50.181 169.615 50.245 ;
			RECT	169.751 50.181 169.783 50.245 ;
			RECT	169.919 50.181 169.951 50.245 ;
			RECT	170.087 50.181 170.119 50.245 ;
			RECT	170.255 50.181 170.287 50.245 ;
			RECT	170.423 50.181 170.455 50.245 ;
			RECT	170.591 50.181 170.623 50.245 ;
			RECT	170.759 50.181 170.791 50.245 ;
			RECT	170.927 50.181 170.959 50.245 ;
			RECT	171.095 50.181 171.127 50.245 ;
			RECT	171.263 50.181 171.295 50.245 ;
			RECT	171.431 50.181 171.463 50.245 ;
			RECT	171.599 50.181 171.631 50.245 ;
			RECT	171.767 50.181 171.799 50.245 ;
			RECT	171.935 50.181 171.967 50.245 ;
			RECT	172.103 50.181 172.135 50.245 ;
			RECT	172.271 50.181 172.303 50.245 ;
			RECT	172.439 50.181 172.471 50.245 ;
			RECT	172.607 50.181 172.639 50.245 ;
			RECT	172.775 50.181 172.807 50.245 ;
			RECT	172.943 50.181 172.975 50.245 ;
			RECT	173.111 50.181 173.143 50.245 ;
			RECT	173.279 50.181 173.311 50.245 ;
			RECT	173.447 50.181 173.479 50.245 ;
			RECT	173.615 50.181 173.647 50.245 ;
			RECT	173.783 50.181 173.815 50.245 ;
			RECT	173.951 50.181 173.983 50.245 ;
			RECT	174.119 50.181 174.151 50.245 ;
			RECT	174.287 50.181 174.319 50.245 ;
			RECT	174.455 50.181 174.487 50.245 ;
			RECT	174.623 50.181 174.655 50.245 ;
			RECT	174.791 50.181 174.823 50.245 ;
			RECT	174.959 50.181 174.991 50.245 ;
			RECT	175.127 50.181 175.159 50.245 ;
			RECT	175.295 50.181 175.327 50.245 ;
			RECT	175.463 50.181 175.495 50.245 ;
			RECT	175.631 50.181 175.663 50.245 ;
			RECT	175.799 50.181 175.831 50.245 ;
			RECT	175.967 50.181 175.999 50.245 ;
			RECT	176.135 50.181 176.167 50.245 ;
			RECT	176.303 50.181 176.335 50.245 ;
			RECT	176.471 50.181 176.503 50.245 ;
			RECT	176.639 50.181 176.671 50.245 ;
			RECT	176.807 50.181 176.839 50.245 ;
			RECT	176.975 50.181 177.007 50.245 ;
			RECT	177.143 50.181 177.175 50.245 ;
			RECT	177.311 50.181 177.343 50.245 ;
			RECT	177.479 50.181 177.511 50.245 ;
			RECT	177.647 50.181 177.679 50.245 ;
			RECT	177.815 50.181 177.847 50.245 ;
			RECT	177.983 50.181 178.015 50.245 ;
			RECT	178.151 50.181 178.183 50.245 ;
			RECT	178.319 50.181 178.351 50.245 ;
			RECT	178.487 50.181 178.519 50.245 ;
			RECT	178.655 50.181 178.687 50.245 ;
			RECT	178.823 50.181 178.855 50.245 ;
			RECT	178.991 50.181 179.023 50.245 ;
			RECT	179.159 50.181 179.191 50.245 ;
			RECT	179.327 50.181 179.359 50.245 ;
			RECT	179.495 50.181 179.527 50.245 ;
			RECT	179.663 50.181 179.695 50.245 ;
			RECT	179.831 50.181 179.863 50.245 ;
			RECT	179.999 50.181 180.031 50.245 ;
			RECT	180.167 50.181 180.199 50.245 ;
			RECT	180.335 50.181 180.367 50.245 ;
			RECT	180.503 50.181 180.535 50.245 ;
			RECT	180.671 50.181 180.703 50.245 ;
			RECT	180.839 50.181 180.871 50.245 ;
			RECT	181.007 50.181 181.039 50.245 ;
			RECT	181.175 50.181 181.207 50.245 ;
			RECT	181.343 50.181 181.375 50.245 ;
			RECT	181.511 50.181 181.543 50.245 ;
			RECT	181.679 50.181 181.711 50.245 ;
			RECT	181.847 50.181 181.879 50.245 ;
			RECT	182.015 50.181 182.047 50.245 ;
			RECT	182.183 50.181 182.215 50.245 ;
			RECT	182.351 50.181 182.383 50.245 ;
			RECT	182.519 50.181 182.551 50.245 ;
			RECT	182.687 50.181 182.719 50.245 ;
			RECT	182.855 50.181 182.887 50.245 ;
			RECT	183.023 50.181 183.055 50.245 ;
			RECT	183.191 50.181 183.223 50.245 ;
			RECT	183.359 50.181 183.391 50.245 ;
			RECT	183.527 50.181 183.559 50.245 ;
			RECT	183.695 50.181 183.727 50.245 ;
			RECT	183.863 50.181 183.895 50.245 ;
			RECT	184.031 50.181 184.063 50.245 ;
			RECT	184.199 50.181 184.231 50.245 ;
			RECT	184.367 50.181 184.399 50.245 ;
			RECT	184.535 50.181 184.567 50.245 ;
			RECT	184.703 50.181 184.735 50.245 ;
			RECT	184.871 50.181 184.903 50.245 ;
			RECT	185.039 50.181 185.071 50.245 ;
			RECT	185.207 50.181 185.239 50.245 ;
			RECT	185.375 50.181 185.407 50.245 ;
			RECT	185.543 50.181 185.575 50.245 ;
			RECT	185.711 50.181 185.743 50.245 ;
			RECT	185.879 50.181 185.911 50.245 ;
			RECT	186.047 50.181 186.079 50.245 ;
			RECT	186.215 50.181 186.247 50.245 ;
			RECT	186.383 50.181 186.415 50.245 ;
			RECT	186.551 50.181 186.583 50.245 ;
			RECT	186.719 50.181 186.751 50.245 ;
			RECT	186.887 50.181 186.919 50.245 ;
			RECT	187.055 50.181 187.087 50.245 ;
			RECT	187.223 50.181 187.255 50.245 ;
			RECT	187.391 50.181 187.423 50.245 ;
			RECT	187.559 50.181 187.591 50.245 ;
			RECT	187.727 50.181 187.759 50.245 ;
			RECT	187.895 50.181 187.927 50.245 ;
			RECT	188.063 50.181 188.095 50.245 ;
			RECT	188.231 50.181 188.263 50.245 ;
			RECT	188.399 50.181 188.431 50.245 ;
			RECT	188.567 50.181 188.599 50.245 ;
			RECT	188.735 50.181 188.767 50.245 ;
			RECT	188.903 50.181 188.935 50.245 ;
			RECT	189.071 50.181 189.103 50.245 ;
			RECT	189.239 50.181 189.271 50.245 ;
			RECT	189.407 50.181 189.439 50.245 ;
			RECT	189.575 50.181 189.607 50.245 ;
			RECT	189.743 50.181 189.775 50.245 ;
			RECT	189.911 50.181 189.943 50.245 ;
			RECT	190.079 50.181 190.111 50.245 ;
			RECT	190.247 50.181 190.279 50.245 ;
			RECT	190.415 50.181 190.447 50.245 ;
			RECT	190.583 50.181 190.615 50.245 ;
			RECT	190.751 50.181 190.783 50.245 ;
			RECT	190.919 50.181 190.951 50.245 ;
			RECT	191.087 50.181 191.119 50.245 ;
			RECT	191.255 50.181 191.287 50.245 ;
			RECT	191.423 50.181 191.455 50.245 ;
			RECT	191.591 50.181 191.623 50.245 ;
			RECT	191.759 50.181 191.791 50.245 ;
			RECT	191.927 50.181 191.959 50.245 ;
			RECT	192.095 50.181 192.127 50.245 ;
			RECT	192.263 50.181 192.295 50.245 ;
			RECT	192.431 50.181 192.463 50.245 ;
			RECT	192.599 50.181 192.631 50.245 ;
			RECT	192.767 50.181 192.799 50.245 ;
			RECT	192.935 50.181 192.967 50.245 ;
			RECT	193.103 50.181 193.135 50.245 ;
			RECT	193.271 50.181 193.303 50.245 ;
			RECT	193.439 50.181 193.471 50.245 ;
			RECT	193.607 50.181 193.639 50.245 ;
			RECT	193.775 50.181 193.807 50.245 ;
			RECT	193.943 50.181 193.975 50.245 ;
			RECT	194.111 50.181 194.143 50.245 ;
			RECT	194.279 50.181 194.311 50.245 ;
			RECT	194.447 50.181 194.479 50.245 ;
			RECT	194.615 50.181 194.647 50.245 ;
			RECT	194.783 50.181 194.815 50.245 ;
			RECT	194.951 50.181 194.983 50.245 ;
			RECT	195.119 50.181 195.151 50.245 ;
			RECT	195.287 50.181 195.319 50.245 ;
			RECT	195.455 50.181 195.487 50.245 ;
			RECT	195.623 50.181 195.655 50.245 ;
			RECT	195.791 50.181 195.823 50.245 ;
			RECT	195.959 50.181 195.991 50.245 ;
			RECT	196.127 50.181 196.159 50.245 ;
			RECT	196.295 50.181 196.327 50.245 ;
			RECT	196.463 50.181 196.495 50.245 ;
			RECT	196.631 50.181 196.663 50.245 ;
			RECT	196.799 50.181 196.831 50.245 ;
			RECT	196.967 50.181 196.999 50.245 ;
			RECT	197.135 50.181 197.167 50.245 ;
			RECT	197.303 50.181 197.335 50.245 ;
			RECT	197.471 50.181 197.503 50.245 ;
			RECT	197.639 50.181 197.671 50.245 ;
			RECT	197.807 50.181 197.839 50.245 ;
			RECT	197.975 50.181 198.007 50.245 ;
			RECT	198.143 50.181 198.175 50.245 ;
			RECT	198.311 50.181 198.343 50.245 ;
			RECT	198.479 50.181 198.511 50.245 ;
			RECT	198.647 50.181 198.679 50.245 ;
			RECT	198.815 50.181 198.847 50.245 ;
			RECT	198.983 50.181 199.015 50.245 ;
			RECT	199.151 50.181 199.183 50.245 ;
			RECT	199.319 50.181 199.351 50.245 ;
			RECT	199.487 50.181 199.519 50.245 ;
			RECT	199.655 50.181 199.687 50.245 ;
			RECT	199.823 50.181 199.855 50.245 ;
			RECT	199.991 50.181 200.023 50.245 ;
			RECT	200.243 50.181 200.275 50.245 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 79.736 201.665 79.856 ;
			LAYER	J3 ;
			RECT	0.755 79.764 0.787 79.828 ;
			RECT	1.645 79.764 1.709 79.828 ;
			RECT	2.323 79.764 2.387 79.828 ;
			RECT	3.438 79.764 3.47 79.828 ;
			RECT	3.585 79.764 3.617 79.828 ;
			RECT	4.195 79.764 4.227 79.828 ;
			RECT	4.72 79.764 4.752 79.828 ;
			RECT	4.944 79.764 5.008 79.828 ;
			RECT	5.267 79.764 5.299 79.828 ;
			RECT	5.797 79.764 5.829 79.828 ;
			RECT	5.927 79.775 5.959 79.807 ;
			RECT	6.049 79.78 6.081 79.812 ;
			RECT	6.179 79.764 6.211 79.828 ;
			RECT	6.347 79.764 6.379 79.828 ;
			RECT	6.515 79.764 6.547 79.828 ;
			RECT	6.683 79.764 6.715 79.828 ;
			RECT	6.851 79.764 6.883 79.828 ;
			RECT	7.019 79.764 7.051 79.828 ;
			RECT	7.187 79.764 7.219 79.828 ;
			RECT	7.355 79.764 7.387 79.828 ;
			RECT	7.523 79.764 7.555 79.828 ;
			RECT	7.691 79.764 7.723 79.828 ;
			RECT	7.859 79.764 7.891 79.828 ;
			RECT	8.027 79.764 8.059 79.828 ;
			RECT	8.195 79.764 8.227 79.828 ;
			RECT	8.363 79.764 8.395 79.828 ;
			RECT	8.531 79.764 8.563 79.828 ;
			RECT	8.699 79.764 8.731 79.828 ;
			RECT	8.867 79.764 8.899 79.828 ;
			RECT	9.035 79.764 9.067 79.828 ;
			RECT	9.203 79.764 9.235 79.828 ;
			RECT	9.371 79.764 9.403 79.828 ;
			RECT	9.539 79.764 9.571 79.828 ;
			RECT	9.707 79.764 9.739 79.828 ;
			RECT	9.875 79.764 9.907 79.828 ;
			RECT	10.043 79.764 10.075 79.828 ;
			RECT	10.211 79.764 10.243 79.828 ;
			RECT	10.379 79.764 10.411 79.828 ;
			RECT	10.547 79.764 10.579 79.828 ;
			RECT	10.715 79.764 10.747 79.828 ;
			RECT	10.883 79.764 10.915 79.828 ;
			RECT	11.051 79.764 11.083 79.828 ;
			RECT	11.219 79.764 11.251 79.828 ;
			RECT	11.387 79.764 11.419 79.828 ;
			RECT	11.555 79.764 11.587 79.828 ;
			RECT	11.723 79.764 11.755 79.828 ;
			RECT	11.891 79.764 11.923 79.828 ;
			RECT	12.059 79.764 12.091 79.828 ;
			RECT	12.227 79.764 12.259 79.828 ;
			RECT	12.395 79.764 12.427 79.828 ;
			RECT	12.563 79.764 12.595 79.828 ;
			RECT	12.731 79.764 12.763 79.828 ;
			RECT	12.899 79.764 12.931 79.828 ;
			RECT	13.067 79.764 13.099 79.828 ;
			RECT	13.235 79.764 13.267 79.828 ;
			RECT	13.403 79.764 13.435 79.828 ;
			RECT	13.571 79.764 13.603 79.828 ;
			RECT	13.739 79.764 13.771 79.828 ;
			RECT	13.907 79.764 13.939 79.828 ;
			RECT	14.075 79.764 14.107 79.828 ;
			RECT	14.243 79.764 14.275 79.828 ;
			RECT	14.411 79.764 14.443 79.828 ;
			RECT	14.579 79.764 14.611 79.828 ;
			RECT	14.747 79.764 14.779 79.828 ;
			RECT	14.915 79.764 14.947 79.828 ;
			RECT	15.083 79.764 15.115 79.828 ;
			RECT	15.251 79.764 15.283 79.828 ;
			RECT	15.419 79.764 15.451 79.828 ;
			RECT	15.587 79.764 15.619 79.828 ;
			RECT	15.755 79.764 15.787 79.828 ;
			RECT	15.923 79.764 15.955 79.828 ;
			RECT	16.091 79.764 16.123 79.828 ;
			RECT	16.259 79.764 16.291 79.828 ;
			RECT	16.427 79.764 16.459 79.828 ;
			RECT	16.595 79.764 16.627 79.828 ;
			RECT	16.763 79.764 16.795 79.828 ;
			RECT	16.931 79.764 16.963 79.828 ;
			RECT	17.099 79.764 17.131 79.828 ;
			RECT	17.267 79.764 17.299 79.828 ;
			RECT	17.435 79.764 17.467 79.828 ;
			RECT	17.603 79.764 17.635 79.828 ;
			RECT	17.771 79.764 17.803 79.828 ;
			RECT	17.939 79.764 17.971 79.828 ;
			RECT	18.107 79.764 18.139 79.828 ;
			RECT	18.275 79.764 18.307 79.828 ;
			RECT	18.443 79.764 18.475 79.828 ;
			RECT	18.611 79.764 18.643 79.828 ;
			RECT	18.779 79.764 18.811 79.828 ;
			RECT	18.947 79.764 18.979 79.828 ;
			RECT	19.115 79.764 19.147 79.828 ;
			RECT	19.283 79.764 19.315 79.828 ;
			RECT	19.451 79.764 19.483 79.828 ;
			RECT	19.619 79.764 19.651 79.828 ;
			RECT	19.787 79.764 19.819 79.828 ;
			RECT	19.955 79.764 19.987 79.828 ;
			RECT	20.123 79.764 20.155 79.828 ;
			RECT	20.291 79.764 20.323 79.828 ;
			RECT	20.459 79.764 20.491 79.828 ;
			RECT	20.627 79.764 20.659 79.828 ;
			RECT	20.795 79.764 20.827 79.828 ;
			RECT	20.963 79.764 20.995 79.828 ;
			RECT	21.131 79.764 21.163 79.828 ;
			RECT	21.299 79.764 21.331 79.828 ;
			RECT	21.467 79.764 21.499 79.828 ;
			RECT	21.635 79.764 21.667 79.828 ;
			RECT	21.803 79.764 21.835 79.828 ;
			RECT	21.971 79.764 22.003 79.828 ;
			RECT	22.139 79.764 22.171 79.828 ;
			RECT	22.307 79.764 22.339 79.828 ;
			RECT	22.475 79.764 22.507 79.828 ;
			RECT	22.643 79.764 22.675 79.828 ;
			RECT	22.811 79.764 22.843 79.828 ;
			RECT	22.979 79.764 23.011 79.828 ;
			RECT	23.147 79.764 23.179 79.828 ;
			RECT	23.315 79.764 23.347 79.828 ;
			RECT	23.483 79.764 23.515 79.828 ;
			RECT	23.651 79.764 23.683 79.828 ;
			RECT	23.819 79.764 23.851 79.828 ;
			RECT	23.987 79.764 24.019 79.828 ;
			RECT	24.155 79.764 24.187 79.828 ;
			RECT	24.323 79.764 24.355 79.828 ;
			RECT	24.491 79.764 24.523 79.828 ;
			RECT	24.659 79.764 24.691 79.828 ;
			RECT	24.827 79.764 24.859 79.828 ;
			RECT	24.995 79.764 25.027 79.828 ;
			RECT	25.163 79.764 25.195 79.828 ;
			RECT	25.331 79.764 25.363 79.828 ;
			RECT	25.499 79.764 25.531 79.828 ;
			RECT	25.667 79.764 25.699 79.828 ;
			RECT	25.835 79.764 25.867 79.828 ;
			RECT	26.003 79.764 26.035 79.828 ;
			RECT	26.171 79.764 26.203 79.828 ;
			RECT	26.339 79.764 26.371 79.828 ;
			RECT	26.507 79.764 26.539 79.828 ;
			RECT	26.675 79.764 26.707 79.828 ;
			RECT	26.843 79.764 26.875 79.828 ;
			RECT	27.011 79.764 27.043 79.828 ;
			RECT	27.179 79.764 27.211 79.828 ;
			RECT	27.347 79.764 27.379 79.828 ;
			RECT	27.515 79.764 27.547 79.828 ;
			RECT	27.683 79.764 27.715 79.828 ;
			RECT	27.851 79.764 27.883 79.828 ;
			RECT	28.019 79.764 28.051 79.828 ;
			RECT	28.187 79.764 28.219 79.828 ;
			RECT	28.355 79.764 28.387 79.828 ;
			RECT	28.523 79.764 28.555 79.828 ;
			RECT	28.691 79.764 28.723 79.828 ;
			RECT	28.859 79.764 28.891 79.828 ;
			RECT	29.027 79.764 29.059 79.828 ;
			RECT	29.195 79.764 29.227 79.828 ;
			RECT	29.363 79.764 29.395 79.828 ;
			RECT	29.531 79.764 29.563 79.828 ;
			RECT	29.699 79.764 29.731 79.828 ;
			RECT	29.867 79.764 29.899 79.828 ;
			RECT	30.035 79.764 30.067 79.828 ;
			RECT	30.203 79.764 30.235 79.828 ;
			RECT	30.371 79.764 30.403 79.828 ;
			RECT	30.539 79.764 30.571 79.828 ;
			RECT	30.707 79.764 30.739 79.828 ;
			RECT	30.875 79.764 30.907 79.828 ;
			RECT	31.043 79.764 31.075 79.828 ;
			RECT	31.211 79.764 31.243 79.828 ;
			RECT	31.379 79.764 31.411 79.828 ;
			RECT	31.547 79.764 31.579 79.828 ;
			RECT	31.715 79.764 31.747 79.828 ;
			RECT	31.883 79.764 31.915 79.828 ;
			RECT	32.051 79.764 32.083 79.828 ;
			RECT	32.219 79.764 32.251 79.828 ;
			RECT	32.387 79.764 32.419 79.828 ;
			RECT	32.555 79.764 32.587 79.828 ;
			RECT	32.723 79.764 32.755 79.828 ;
			RECT	32.891 79.764 32.923 79.828 ;
			RECT	33.059 79.764 33.091 79.828 ;
			RECT	33.227 79.764 33.259 79.828 ;
			RECT	33.395 79.764 33.427 79.828 ;
			RECT	33.563 79.764 33.595 79.828 ;
			RECT	33.731 79.764 33.763 79.828 ;
			RECT	33.899 79.764 33.931 79.828 ;
			RECT	34.067 79.764 34.099 79.828 ;
			RECT	34.235 79.764 34.267 79.828 ;
			RECT	34.403 79.764 34.435 79.828 ;
			RECT	34.571 79.764 34.603 79.828 ;
			RECT	34.739 79.764 34.771 79.828 ;
			RECT	34.907 79.764 34.939 79.828 ;
			RECT	35.075 79.764 35.107 79.828 ;
			RECT	35.243 79.764 35.275 79.828 ;
			RECT	35.411 79.764 35.443 79.828 ;
			RECT	35.579 79.764 35.611 79.828 ;
			RECT	35.747 79.764 35.779 79.828 ;
			RECT	35.915 79.764 35.947 79.828 ;
			RECT	36.083 79.764 36.115 79.828 ;
			RECT	36.251 79.764 36.283 79.828 ;
			RECT	36.419 79.764 36.451 79.828 ;
			RECT	36.587 79.764 36.619 79.828 ;
			RECT	36.755 79.764 36.787 79.828 ;
			RECT	36.923 79.764 36.955 79.828 ;
			RECT	37.091 79.764 37.123 79.828 ;
			RECT	37.259 79.764 37.291 79.828 ;
			RECT	37.427 79.764 37.459 79.828 ;
			RECT	37.595 79.764 37.627 79.828 ;
			RECT	37.763 79.764 37.795 79.828 ;
			RECT	37.931 79.764 37.963 79.828 ;
			RECT	38.099 79.764 38.131 79.828 ;
			RECT	38.267 79.764 38.299 79.828 ;
			RECT	38.435 79.764 38.467 79.828 ;
			RECT	38.603 79.764 38.635 79.828 ;
			RECT	38.771 79.764 38.803 79.828 ;
			RECT	38.939 79.764 38.971 79.828 ;
			RECT	39.107 79.764 39.139 79.828 ;
			RECT	39.275 79.764 39.307 79.828 ;
			RECT	39.443 79.764 39.475 79.828 ;
			RECT	39.611 79.764 39.643 79.828 ;
			RECT	39.779 79.764 39.811 79.828 ;
			RECT	39.947 79.764 39.979 79.828 ;
			RECT	40.115 79.764 40.147 79.828 ;
			RECT	40.283 79.764 40.315 79.828 ;
			RECT	40.451 79.764 40.483 79.828 ;
			RECT	40.619 79.764 40.651 79.828 ;
			RECT	40.787 79.764 40.819 79.828 ;
			RECT	40.955 79.764 40.987 79.828 ;
			RECT	41.123 79.764 41.155 79.828 ;
			RECT	41.291 79.764 41.323 79.828 ;
			RECT	41.459 79.764 41.491 79.828 ;
			RECT	41.627 79.764 41.659 79.828 ;
			RECT	41.795 79.764 41.827 79.828 ;
			RECT	41.963 79.764 41.995 79.828 ;
			RECT	42.131 79.764 42.163 79.828 ;
			RECT	42.299 79.764 42.331 79.828 ;
			RECT	42.467 79.764 42.499 79.828 ;
			RECT	42.635 79.764 42.667 79.828 ;
			RECT	42.803 79.764 42.835 79.828 ;
			RECT	42.971 79.764 43.003 79.828 ;
			RECT	43.139 79.764 43.171 79.828 ;
			RECT	43.307 79.764 43.339 79.828 ;
			RECT	43.475 79.764 43.507 79.828 ;
			RECT	43.643 79.764 43.675 79.828 ;
			RECT	43.811 79.764 43.843 79.828 ;
			RECT	43.979 79.764 44.011 79.828 ;
			RECT	44.147 79.764 44.179 79.828 ;
			RECT	44.315 79.764 44.347 79.828 ;
			RECT	44.483 79.764 44.515 79.828 ;
			RECT	44.651 79.764 44.683 79.828 ;
			RECT	44.819 79.764 44.851 79.828 ;
			RECT	44.987 79.764 45.019 79.828 ;
			RECT	45.155 79.764 45.187 79.828 ;
			RECT	45.323 79.764 45.355 79.828 ;
			RECT	45.491 79.764 45.523 79.828 ;
			RECT	45.659 79.764 45.691 79.828 ;
			RECT	45.827 79.764 45.859 79.828 ;
			RECT	45.995 79.764 46.027 79.828 ;
			RECT	46.163 79.764 46.195 79.828 ;
			RECT	46.331 79.764 46.363 79.828 ;
			RECT	46.499 79.764 46.531 79.828 ;
			RECT	46.667 79.764 46.699 79.828 ;
			RECT	46.835 79.764 46.867 79.828 ;
			RECT	47.003 79.764 47.035 79.828 ;
			RECT	47.171 79.764 47.203 79.828 ;
			RECT	47.339 79.764 47.371 79.828 ;
			RECT	47.507 79.764 47.539 79.828 ;
			RECT	47.675 79.764 47.707 79.828 ;
			RECT	47.843 79.764 47.875 79.828 ;
			RECT	48.011 79.764 48.043 79.828 ;
			RECT	48.179 79.764 48.211 79.828 ;
			RECT	48.347 79.764 48.379 79.828 ;
			RECT	48.515 79.764 48.547 79.828 ;
			RECT	48.683 79.764 48.715 79.828 ;
			RECT	48.851 79.764 48.883 79.828 ;
			RECT	49.019 79.764 49.051 79.828 ;
			RECT	49.187 79.764 49.219 79.828 ;
			RECT	49.318 79.78 49.35 79.812 ;
			RECT	49.439 79.78 49.471 79.812 ;
			RECT	49.569 79.764 49.601 79.828 ;
			RECT	51.881 79.764 51.913 79.828 ;
			RECT	53.132 79.764 53.196 79.828 ;
			RECT	53.812 79.764 53.844 79.828 ;
			RECT	54.251 79.764 54.283 79.828 ;
			RECT	55.562 79.764 55.626 79.828 ;
			RECT	58.603 79.764 58.635 79.828 ;
			RECT	58.733 79.78 58.765 79.812 ;
			RECT	58.854 79.78 58.886 79.812 ;
			RECT	58.985 79.764 59.017 79.828 ;
			RECT	59.153 79.764 59.185 79.828 ;
			RECT	59.321 79.764 59.353 79.828 ;
			RECT	59.489 79.764 59.521 79.828 ;
			RECT	59.657 79.764 59.689 79.828 ;
			RECT	59.825 79.764 59.857 79.828 ;
			RECT	59.993 79.764 60.025 79.828 ;
			RECT	60.161 79.764 60.193 79.828 ;
			RECT	60.329 79.764 60.361 79.828 ;
			RECT	60.497 79.764 60.529 79.828 ;
			RECT	60.665 79.764 60.697 79.828 ;
			RECT	60.833 79.764 60.865 79.828 ;
			RECT	61.001 79.764 61.033 79.828 ;
			RECT	61.169 79.764 61.201 79.828 ;
			RECT	61.337 79.764 61.369 79.828 ;
			RECT	61.505 79.764 61.537 79.828 ;
			RECT	61.673 79.764 61.705 79.828 ;
			RECT	61.841 79.764 61.873 79.828 ;
			RECT	62.009 79.764 62.041 79.828 ;
			RECT	62.177 79.764 62.209 79.828 ;
			RECT	62.345 79.764 62.377 79.828 ;
			RECT	62.513 79.764 62.545 79.828 ;
			RECT	62.681 79.764 62.713 79.828 ;
			RECT	62.849 79.764 62.881 79.828 ;
			RECT	63.017 79.764 63.049 79.828 ;
			RECT	63.185 79.764 63.217 79.828 ;
			RECT	63.353 79.764 63.385 79.828 ;
			RECT	63.521 79.764 63.553 79.828 ;
			RECT	63.689 79.764 63.721 79.828 ;
			RECT	63.857 79.764 63.889 79.828 ;
			RECT	64.025 79.764 64.057 79.828 ;
			RECT	64.193 79.764 64.225 79.828 ;
			RECT	64.361 79.764 64.393 79.828 ;
			RECT	64.529 79.764 64.561 79.828 ;
			RECT	64.697 79.764 64.729 79.828 ;
			RECT	64.865 79.764 64.897 79.828 ;
			RECT	65.033 79.764 65.065 79.828 ;
			RECT	65.201 79.764 65.233 79.828 ;
			RECT	65.369 79.764 65.401 79.828 ;
			RECT	65.537 79.764 65.569 79.828 ;
			RECT	65.705 79.764 65.737 79.828 ;
			RECT	65.873 79.764 65.905 79.828 ;
			RECT	66.041 79.764 66.073 79.828 ;
			RECT	66.209 79.764 66.241 79.828 ;
			RECT	66.377 79.764 66.409 79.828 ;
			RECT	66.545 79.764 66.577 79.828 ;
			RECT	66.713 79.764 66.745 79.828 ;
			RECT	66.881 79.764 66.913 79.828 ;
			RECT	67.049 79.764 67.081 79.828 ;
			RECT	67.217 79.764 67.249 79.828 ;
			RECT	67.385 79.764 67.417 79.828 ;
			RECT	67.553 79.764 67.585 79.828 ;
			RECT	67.721 79.764 67.753 79.828 ;
			RECT	67.889 79.764 67.921 79.828 ;
			RECT	68.057 79.764 68.089 79.828 ;
			RECT	68.225 79.764 68.257 79.828 ;
			RECT	68.393 79.764 68.425 79.828 ;
			RECT	68.561 79.764 68.593 79.828 ;
			RECT	68.729 79.764 68.761 79.828 ;
			RECT	68.897 79.764 68.929 79.828 ;
			RECT	69.065 79.764 69.097 79.828 ;
			RECT	69.233 79.764 69.265 79.828 ;
			RECT	69.401 79.764 69.433 79.828 ;
			RECT	69.569 79.764 69.601 79.828 ;
			RECT	69.737 79.764 69.769 79.828 ;
			RECT	69.905 79.764 69.937 79.828 ;
			RECT	70.073 79.764 70.105 79.828 ;
			RECT	70.241 79.764 70.273 79.828 ;
			RECT	70.409 79.764 70.441 79.828 ;
			RECT	70.577 79.764 70.609 79.828 ;
			RECT	70.745 79.764 70.777 79.828 ;
			RECT	70.913 79.764 70.945 79.828 ;
			RECT	71.081 79.764 71.113 79.828 ;
			RECT	71.249 79.764 71.281 79.828 ;
			RECT	71.417 79.764 71.449 79.828 ;
			RECT	71.585 79.764 71.617 79.828 ;
			RECT	71.753 79.764 71.785 79.828 ;
			RECT	71.921 79.764 71.953 79.828 ;
			RECT	72.089 79.764 72.121 79.828 ;
			RECT	72.257 79.764 72.289 79.828 ;
			RECT	72.425 79.764 72.457 79.828 ;
			RECT	72.593 79.764 72.625 79.828 ;
			RECT	72.761 79.764 72.793 79.828 ;
			RECT	72.929 79.764 72.961 79.828 ;
			RECT	73.097 79.764 73.129 79.828 ;
			RECT	73.265 79.764 73.297 79.828 ;
			RECT	73.433 79.764 73.465 79.828 ;
			RECT	73.601 79.764 73.633 79.828 ;
			RECT	73.769 79.764 73.801 79.828 ;
			RECT	73.937 79.764 73.969 79.828 ;
			RECT	74.105 79.764 74.137 79.828 ;
			RECT	74.273 79.764 74.305 79.828 ;
			RECT	74.441 79.764 74.473 79.828 ;
			RECT	74.609 79.764 74.641 79.828 ;
			RECT	74.777 79.764 74.809 79.828 ;
			RECT	74.945 79.764 74.977 79.828 ;
			RECT	75.113 79.764 75.145 79.828 ;
			RECT	75.281 79.764 75.313 79.828 ;
			RECT	75.449 79.764 75.481 79.828 ;
			RECT	75.617 79.764 75.649 79.828 ;
			RECT	75.785 79.764 75.817 79.828 ;
			RECT	75.953 79.764 75.985 79.828 ;
			RECT	76.121 79.764 76.153 79.828 ;
			RECT	76.289 79.764 76.321 79.828 ;
			RECT	76.457 79.764 76.489 79.828 ;
			RECT	76.625 79.764 76.657 79.828 ;
			RECT	76.793 79.764 76.825 79.828 ;
			RECT	76.961 79.764 76.993 79.828 ;
			RECT	77.129 79.764 77.161 79.828 ;
			RECT	77.297 79.764 77.329 79.828 ;
			RECT	77.465 79.764 77.497 79.828 ;
			RECT	77.633 79.764 77.665 79.828 ;
			RECT	77.801 79.764 77.833 79.828 ;
			RECT	77.969 79.764 78.001 79.828 ;
			RECT	78.137 79.764 78.169 79.828 ;
			RECT	78.305 79.764 78.337 79.828 ;
			RECT	78.473 79.764 78.505 79.828 ;
			RECT	78.641 79.764 78.673 79.828 ;
			RECT	78.809 79.764 78.841 79.828 ;
			RECT	78.977 79.764 79.009 79.828 ;
			RECT	79.145 79.764 79.177 79.828 ;
			RECT	79.313 79.764 79.345 79.828 ;
			RECT	79.481 79.764 79.513 79.828 ;
			RECT	79.649 79.764 79.681 79.828 ;
			RECT	79.817 79.764 79.849 79.828 ;
			RECT	79.985 79.764 80.017 79.828 ;
			RECT	80.153 79.764 80.185 79.828 ;
			RECT	80.321 79.764 80.353 79.828 ;
			RECT	80.489 79.764 80.521 79.828 ;
			RECT	80.657 79.764 80.689 79.828 ;
			RECT	80.825 79.764 80.857 79.828 ;
			RECT	80.993 79.764 81.025 79.828 ;
			RECT	81.161 79.764 81.193 79.828 ;
			RECT	81.329 79.764 81.361 79.828 ;
			RECT	81.497 79.764 81.529 79.828 ;
			RECT	81.665 79.764 81.697 79.828 ;
			RECT	81.833 79.764 81.865 79.828 ;
			RECT	82.001 79.764 82.033 79.828 ;
			RECT	82.169 79.764 82.201 79.828 ;
			RECT	82.337 79.764 82.369 79.828 ;
			RECT	82.505 79.764 82.537 79.828 ;
			RECT	82.673 79.764 82.705 79.828 ;
			RECT	82.841 79.764 82.873 79.828 ;
			RECT	83.009 79.764 83.041 79.828 ;
			RECT	83.177 79.764 83.209 79.828 ;
			RECT	83.345 79.764 83.377 79.828 ;
			RECT	83.513 79.764 83.545 79.828 ;
			RECT	83.681 79.764 83.713 79.828 ;
			RECT	83.849 79.764 83.881 79.828 ;
			RECT	84.017 79.764 84.049 79.828 ;
			RECT	84.185 79.764 84.217 79.828 ;
			RECT	84.353 79.764 84.385 79.828 ;
			RECT	84.521 79.764 84.553 79.828 ;
			RECT	84.689 79.764 84.721 79.828 ;
			RECT	84.857 79.764 84.889 79.828 ;
			RECT	85.025 79.764 85.057 79.828 ;
			RECT	85.193 79.764 85.225 79.828 ;
			RECT	85.361 79.764 85.393 79.828 ;
			RECT	85.529 79.764 85.561 79.828 ;
			RECT	85.697 79.764 85.729 79.828 ;
			RECT	85.865 79.764 85.897 79.828 ;
			RECT	86.033 79.764 86.065 79.828 ;
			RECT	86.201 79.764 86.233 79.828 ;
			RECT	86.369 79.764 86.401 79.828 ;
			RECT	86.537 79.764 86.569 79.828 ;
			RECT	86.705 79.764 86.737 79.828 ;
			RECT	86.873 79.764 86.905 79.828 ;
			RECT	87.041 79.764 87.073 79.828 ;
			RECT	87.209 79.764 87.241 79.828 ;
			RECT	87.377 79.764 87.409 79.828 ;
			RECT	87.545 79.764 87.577 79.828 ;
			RECT	87.713 79.764 87.745 79.828 ;
			RECT	87.881 79.764 87.913 79.828 ;
			RECT	88.049 79.764 88.081 79.828 ;
			RECT	88.217 79.764 88.249 79.828 ;
			RECT	88.385 79.764 88.417 79.828 ;
			RECT	88.553 79.764 88.585 79.828 ;
			RECT	88.721 79.764 88.753 79.828 ;
			RECT	88.889 79.764 88.921 79.828 ;
			RECT	89.057 79.764 89.089 79.828 ;
			RECT	89.225 79.764 89.257 79.828 ;
			RECT	89.393 79.764 89.425 79.828 ;
			RECT	89.561 79.764 89.593 79.828 ;
			RECT	89.729 79.764 89.761 79.828 ;
			RECT	89.897 79.764 89.929 79.828 ;
			RECT	90.065 79.764 90.097 79.828 ;
			RECT	90.233 79.764 90.265 79.828 ;
			RECT	90.401 79.764 90.433 79.828 ;
			RECT	90.569 79.764 90.601 79.828 ;
			RECT	90.737 79.764 90.769 79.828 ;
			RECT	90.905 79.764 90.937 79.828 ;
			RECT	91.073 79.764 91.105 79.828 ;
			RECT	91.241 79.764 91.273 79.828 ;
			RECT	91.409 79.764 91.441 79.828 ;
			RECT	91.577 79.764 91.609 79.828 ;
			RECT	91.745 79.764 91.777 79.828 ;
			RECT	91.913 79.764 91.945 79.828 ;
			RECT	92.081 79.764 92.113 79.828 ;
			RECT	92.249 79.764 92.281 79.828 ;
			RECT	92.417 79.764 92.449 79.828 ;
			RECT	92.585 79.764 92.617 79.828 ;
			RECT	92.753 79.764 92.785 79.828 ;
			RECT	92.921 79.764 92.953 79.828 ;
			RECT	93.089 79.764 93.121 79.828 ;
			RECT	93.257 79.764 93.289 79.828 ;
			RECT	93.425 79.764 93.457 79.828 ;
			RECT	93.593 79.764 93.625 79.828 ;
			RECT	93.761 79.764 93.793 79.828 ;
			RECT	93.929 79.764 93.961 79.828 ;
			RECT	94.097 79.764 94.129 79.828 ;
			RECT	94.265 79.764 94.297 79.828 ;
			RECT	94.433 79.764 94.465 79.828 ;
			RECT	94.601 79.764 94.633 79.828 ;
			RECT	94.769 79.764 94.801 79.828 ;
			RECT	94.937 79.764 94.969 79.828 ;
			RECT	95.105 79.764 95.137 79.828 ;
			RECT	95.273 79.764 95.305 79.828 ;
			RECT	95.441 79.764 95.473 79.828 ;
			RECT	95.609 79.764 95.641 79.828 ;
			RECT	95.777 79.764 95.809 79.828 ;
			RECT	95.945 79.764 95.977 79.828 ;
			RECT	96.113 79.764 96.145 79.828 ;
			RECT	96.281 79.764 96.313 79.828 ;
			RECT	96.449 79.764 96.481 79.828 ;
			RECT	96.617 79.764 96.649 79.828 ;
			RECT	96.785 79.764 96.817 79.828 ;
			RECT	96.953 79.764 96.985 79.828 ;
			RECT	97.121 79.764 97.153 79.828 ;
			RECT	97.289 79.764 97.321 79.828 ;
			RECT	97.457 79.764 97.489 79.828 ;
			RECT	97.625 79.764 97.657 79.828 ;
			RECT	97.793 79.764 97.825 79.828 ;
			RECT	97.961 79.764 97.993 79.828 ;
			RECT	98.129 79.764 98.161 79.828 ;
			RECT	98.297 79.764 98.329 79.828 ;
			RECT	98.465 79.764 98.497 79.828 ;
			RECT	98.633 79.764 98.665 79.828 ;
			RECT	98.801 79.764 98.833 79.828 ;
			RECT	98.969 79.764 99.001 79.828 ;
			RECT	99.137 79.764 99.169 79.828 ;
			RECT	99.305 79.764 99.337 79.828 ;
			RECT	99.473 79.764 99.505 79.828 ;
			RECT	99.641 79.764 99.673 79.828 ;
			RECT	99.809 79.764 99.841 79.828 ;
			RECT	99.977 79.764 100.009 79.828 ;
			RECT	100.145 79.764 100.177 79.828 ;
			RECT	100.313 79.764 100.345 79.828 ;
			RECT	100.481 79.764 100.513 79.828 ;
			RECT	100.649 79.764 100.681 79.828 ;
			RECT	100.817 79.764 100.849 79.828 ;
			RECT	100.985 79.764 101.017 79.828 ;
			RECT	101.153 79.764 101.185 79.828 ;
			RECT	101.321 79.764 101.353 79.828 ;
			RECT	101.489 79.764 101.521 79.828 ;
			RECT	101.657 79.764 101.689 79.828 ;
			RECT	101.825 79.764 101.857 79.828 ;
			RECT	101.993 79.764 102.025 79.828 ;
			RECT	102.123 79.78 102.155 79.812 ;
			RECT	102.245 79.775 102.277 79.807 ;
			RECT	102.375 79.764 102.407 79.828 ;
			RECT	103.795 79.764 103.827 79.828 ;
			RECT	103.925 79.775 103.957 79.807 ;
			RECT	104.047 79.78 104.079 79.812 ;
			RECT	104.177 79.764 104.209 79.828 ;
			RECT	104.345 79.764 104.377 79.828 ;
			RECT	104.513 79.764 104.545 79.828 ;
			RECT	104.681 79.764 104.713 79.828 ;
			RECT	104.849 79.764 104.881 79.828 ;
			RECT	105.017 79.764 105.049 79.828 ;
			RECT	105.185 79.764 105.217 79.828 ;
			RECT	105.353 79.764 105.385 79.828 ;
			RECT	105.521 79.764 105.553 79.828 ;
			RECT	105.689 79.764 105.721 79.828 ;
			RECT	105.857 79.764 105.889 79.828 ;
			RECT	106.025 79.764 106.057 79.828 ;
			RECT	106.193 79.764 106.225 79.828 ;
			RECT	106.361 79.764 106.393 79.828 ;
			RECT	106.529 79.764 106.561 79.828 ;
			RECT	106.697 79.764 106.729 79.828 ;
			RECT	106.865 79.764 106.897 79.828 ;
			RECT	107.033 79.764 107.065 79.828 ;
			RECT	107.201 79.764 107.233 79.828 ;
			RECT	107.369 79.764 107.401 79.828 ;
			RECT	107.537 79.764 107.569 79.828 ;
			RECT	107.705 79.764 107.737 79.828 ;
			RECT	107.873 79.764 107.905 79.828 ;
			RECT	108.041 79.764 108.073 79.828 ;
			RECT	108.209 79.764 108.241 79.828 ;
			RECT	108.377 79.764 108.409 79.828 ;
			RECT	108.545 79.764 108.577 79.828 ;
			RECT	108.713 79.764 108.745 79.828 ;
			RECT	108.881 79.764 108.913 79.828 ;
			RECT	109.049 79.764 109.081 79.828 ;
			RECT	109.217 79.764 109.249 79.828 ;
			RECT	109.385 79.764 109.417 79.828 ;
			RECT	109.553 79.764 109.585 79.828 ;
			RECT	109.721 79.764 109.753 79.828 ;
			RECT	109.889 79.764 109.921 79.828 ;
			RECT	110.057 79.764 110.089 79.828 ;
			RECT	110.225 79.764 110.257 79.828 ;
			RECT	110.393 79.764 110.425 79.828 ;
			RECT	110.561 79.764 110.593 79.828 ;
			RECT	110.729 79.764 110.761 79.828 ;
			RECT	110.897 79.764 110.929 79.828 ;
			RECT	111.065 79.764 111.097 79.828 ;
			RECT	111.233 79.764 111.265 79.828 ;
			RECT	111.401 79.764 111.433 79.828 ;
			RECT	111.569 79.764 111.601 79.828 ;
			RECT	111.737 79.764 111.769 79.828 ;
			RECT	111.905 79.764 111.937 79.828 ;
			RECT	112.073 79.764 112.105 79.828 ;
			RECT	112.241 79.764 112.273 79.828 ;
			RECT	112.409 79.764 112.441 79.828 ;
			RECT	112.577 79.764 112.609 79.828 ;
			RECT	112.745 79.764 112.777 79.828 ;
			RECT	112.913 79.764 112.945 79.828 ;
			RECT	113.081 79.764 113.113 79.828 ;
			RECT	113.249 79.764 113.281 79.828 ;
			RECT	113.417 79.764 113.449 79.828 ;
			RECT	113.585 79.764 113.617 79.828 ;
			RECT	113.753 79.764 113.785 79.828 ;
			RECT	113.921 79.764 113.953 79.828 ;
			RECT	114.089 79.764 114.121 79.828 ;
			RECT	114.257 79.764 114.289 79.828 ;
			RECT	114.425 79.764 114.457 79.828 ;
			RECT	114.593 79.764 114.625 79.828 ;
			RECT	114.761 79.764 114.793 79.828 ;
			RECT	114.929 79.764 114.961 79.828 ;
			RECT	115.097 79.764 115.129 79.828 ;
			RECT	115.265 79.764 115.297 79.828 ;
			RECT	115.433 79.764 115.465 79.828 ;
			RECT	115.601 79.764 115.633 79.828 ;
			RECT	115.769 79.764 115.801 79.828 ;
			RECT	115.937 79.764 115.969 79.828 ;
			RECT	116.105 79.764 116.137 79.828 ;
			RECT	116.273 79.764 116.305 79.828 ;
			RECT	116.441 79.764 116.473 79.828 ;
			RECT	116.609 79.764 116.641 79.828 ;
			RECT	116.777 79.764 116.809 79.828 ;
			RECT	116.945 79.764 116.977 79.828 ;
			RECT	117.113 79.764 117.145 79.828 ;
			RECT	117.281 79.764 117.313 79.828 ;
			RECT	117.449 79.764 117.481 79.828 ;
			RECT	117.617 79.764 117.649 79.828 ;
			RECT	117.785 79.764 117.817 79.828 ;
			RECT	117.953 79.764 117.985 79.828 ;
			RECT	118.121 79.764 118.153 79.828 ;
			RECT	118.289 79.764 118.321 79.828 ;
			RECT	118.457 79.764 118.489 79.828 ;
			RECT	118.625 79.764 118.657 79.828 ;
			RECT	118.793 79.764 118.825 79.828 ;
			RECT	118.961 79.764 118.993 79.828 ;
			RECT	119.129 79.764 119.161 79.828 ;
			RECT	119.297 79.764 119.329 79.828 ;
			RECT	119.465 79.764 119.497 79.828 ;
			RECT	119.633 79.764 119.665 79.828 ;
			RECT	119.801 79.764 119.833 79.828 ;
			RECT	119.969 79.764 120.001 79.828 ;
			RECT	120.137 79.764 120.169 79.828 ;
			RECT	120.305 79.764 120.337 79.828 ;
			RECT	120.473 79.764 120.505 79.828 ;
			RECT	120.641 79.764 120.673 79.828 ;
			RECT	120.809 79.764 120.841 79.828 ;
			RECT	120.977 79.764 121.009 79.828 ;
			RECT	121.145 79.764 121.177 79.828 ;
			RECT	121.313 79.764 121.345 79.828 ;
			RECT	121.481 79.764 121.513 79.828 ;
			RECT	121.649 79.764 121.681 79.828 ;
			RECT	121.817 79.764 121.849 79.828 ;
			RECT	121.985 79.764 122.017 79.828 ;
			RECT	122.153 79.764 122.185 79.828 ;
			RECT	122.321 79.764 122.353 79.828 ;
			RECT	122.489 79.764 122.521 79.828 ;
			RECT	122.657 79.764 122.689 79.828 ;
			RECT	122.825 79.764 122.857 79.828 ;
			RECT	122.993 79.764 123.025 79.828 ;
			RECT	123.161 79.764 123.193 79.828 ;
			RECT	123.329 79.764 123.361 79.828 ;
			RECT	123.497 79.764 123.529 79.828 ;
			RECT	123.665 79.764 123.697 79.828 ;
			RECT	123.833 79.764 123.865 79.828 ;
			RECT	124.001 79.764 124.033 79.828 ;
			RECT	124.169 79.764 124.201 79.828 ;
			RECT	124.337 79.764 124.369 79.828 ;
			RECT	124.505 79.764 124.537 79.828 ;
			RECT	124.673 79.764 124.705 79.828 ;
			RECT	124.841 79.764 124.873 79.828 ;
			RECT	125.009 79.764 125.041 79.828 ;
			RECT	125.177 79.764 125.209 79.828 ;
			RECT	125.345 79.764 125.377 79.828 ;
			RECT	125.513 79.764 125.545 79.828 ;
			RECT	125.681 79.764 125.713 79.828 ;
			RECT	125.849 79.764 125.881 79.828 ;
			RECT	126.017 79.764 126.049 79.828 ;
			RECT	126.185 79.764 126.217 79.828 ;
			RECT	126.353 79.764 126.385 79.828 ;
			RECT	126.521 79.764 126.553 79.828 ;
			RECT	126.689 79.764 126.721 79.828 ;
			RECT	126.857 79.764 126.889 79.828 ;
			RECT	127.025 79.764 127.057 79.828 ;
			RECT	127.193 79.764 127.225 79.828 ;
			RECT	127.361 79.764 127.393 79.828 ;
			RECT	127.529 79.764 127.561 79.828 ;
			RECT	127.697 79.764 127.729 79.828 ;
			RECT	127.865 79.764 127.897 79.828 ;
			RECT	128.033 79.764 128.065 79.828 ;
			RECT	128.201 79.764 128.233 79.828 ;
			RECT	128.369 79.764 128.401 79.828 ;
			RECT	128.537 79.764 128.569 79.828 ;
			RECT	128.705 79.764 128.737 79.828 ;
			RECT	128.873 79.764 128.905 79.828 ;
			RECT	129.041 79.764 129.073 79.828 ;
			RECT	129.209 79.764 129.241 79.828 ;
			RECT	129.377 79.764 129.409 79.828 ;
			RECT	129.545 79.764 129.577 79.828 ;
			RECT	129.713 79.764 129.745 79.828 ;
			RECT	129.881 79.764 129.913 79.828 ;
			RECT	130.049 79.764 130.081 79.828 ;
			RECT	130.217 79.764 130.249 79.828 ;
			RECT	130.385 79.764 130.417 79.828 ;
			RECT	130.553 79.764 130.585 79.828 ;
			RECT	130.721 79.764 130.753 79.828 ;
			RECT	130.889 79.764 130.921 79.828 ;
			RECT	131.057 79.764 131.089 79.828 ;
			RECT	131.225 79.764 131.257 79.828 ;
			RECT	131.393 79.764 131.425 79.828 ;
			RECT	131.561 79.764 131.593 79.828 ;
			RECT	131.729 79.764 131.761 79.828 ;
			RECT	131.897 79.764 131.929 79.828 ;
			RECT	132.065 79.764 132.097 79.828 ;
			RECT	132.233 79.764 132.265 79.828 ;
			RECT	132.401 79.764 132.433 79.828 ;
			RECT	132.569 79.764 132.601 79.828 ;
			RECT	132.737 79.764 132.769 79.828 ;
			RECT	132.905 79.764 132.937 79.828 ;
			RECT	133.073 79.764 133.105 79.828 ;
			RECT	133.241 79.764 133.273 79.828 ;
			RECT	133.409 79.764 133.441 79.828 ;
			RECT	133.577 79.764 133.609 79.828 ;
			RECT	133.745 79.764 133.777 79.828 ;
			RECT	133.913 79.764 133.945 79.828 ;
			RECT	134.081 79.764 134.113 79.828 ;
			RECT	134.249 79.764 134.281 79.828 ;
			RECT	134.417 79.764 134.449 79.828 ;
			RECT	134.585 79.764 134.617 79.828 ;
			RECT	134.753 79.764 134.785 79.828 ;
			RECT	134.921 79.764 134.953 79.828 ;
			RECT	135.089 79.764 135.121 79.828 ;
			RECT	135.257 79.764 135.289 79.828 ;
			RECT	135.425 79.764 135.457 79.828 ;
			RECT	135.593 79.764 135.625 79.828 ;
			RECT	135.761 79.764 135.793 79.828 ;
			RECT	135.929 79.764 135.961 79.828 ;
			RECT	136.097 79.764 136.129 79.828 ;
			RECT	136.265 79.764 136.297 79.828 ;
			RECT	136.433 79.764 136.465 79.828 ;
			RECT	136.601 79.764 136.633 79.828 ;
			RECT	136.769 79.764 136.801 79.828 ;
			RECT	136.937 79.764 136.969 79.828 ;
			RECT	137.105 79.764 137.137 79.828 ;
			RECT	137.273 79.764 137.305 79.828 ;
			RECT	137.441 79.764 137.473 79.828 ;
			RECT	137.609 79.764 137.641 79.828 ;
			RECT	137.777 79.764 137.809 79.828 ;
			RECT	137.945 79.764 137.977 79.828 ;
			RECT	138.113 79.764 138.145 79.828 ;
			RECT	138.281 79.764 138.313 79.828 ;
			RECT	138.449 79.764 138.481 79.828 ;
			RECT	138.617 79.764 138.649 79.828 ;
			RECT	138.785 79.764 138.817 79.828 ;
			RECT	138.953 79.764 138.985 79.828 ;
			RECT	139.121 79.764 139.153 79.828 ;
			RECT	139.289 79.764 139.321 79.828 ;
			RECT	139.457 79.764 139.489 79.828 ;
			RECT	139.625 79.764 139.657 79.828 ;
			RECT	139.793 79.764 139.825 79.828 ;
			RECT	139.961 79.764 139.993 79.828 ;
			RECT	140.129 79.764 140.161 79.828 ;
			RECT	140.297 79.764 140.329 79.828 ;
			RECT	140.465 79.764 140.497 79.828 ;
			RECT	140.633 79.764 140.665 79.828 ;
			RECT	140.801 79.764 140.833 79.828 ;
			RECT	140.969 79.764 141.001 79.828 ;
			RECT	141.137 79.764 141.169 79.828 ;
			RECT	141.305 79.764 141.337 79.828 ;
			RECT	141.473 79.764 141.505 79.828 ;
			RECT	141.641 79.764 141.673 79.828 ;
			RECT	141.809 79.764 141.841 79.828 ;
			RECT	141.977 79.764 142.009 79.828 ;
			RECT	142.145 79.764 142.177 79.828 ;
			RECT	142.313 79.764 142.345 79.828 ;
			RECT	142.481 79.764 142.513 79.828 ;
			RECT	142.649 79.764 142.681 79.828 ;
			RECT	142.817 79.764 142.849 79.828 ;
			RECT	142.985 79.764 143.017 79.828 ;
			RECT	143.153 79.764 143.185 79.828 ;
			RECT	143.321 79.764 143.353 79.828 ;
			RECT	143.489 79.764 143.521 79.828 ;
			RECT	143.657 79.764 143.689 79.828 ;
			RECT	143.825 79.764 143.857 79.828 ;
			RECT	143.993 79.764 144.025 79.828 ;
			RECT	144.161 79.764 144.193 79.828 ;
			RECT	144.329 79.764 144.361 79.828 ;
			RECT	144.497 79.764 144.529 79.828 ;
			RECT	144.665 79.764 144.697 79.828 ;
			RECT	144.833 79.764 144.865 79.828 ;
			RECT	145.001 79.764 145.033 79.828 ;
			RECT	145.169 79.764 145.201 79.828 ;
			RECT	145.337 79.764 145.369 79.828 ;
			RECT	145.505 79.764 145.537 79.828 ;
			RECT	145.673 79.764 145.705 79.828 ;
			RECT	145.841 79.764 145.873 79.828 ;
			RECT	146.009 79.764 146.041 79.828 ;
			RECT	146.177 79.764 146.209 79.828 ;
			RECT	146.345 79.764 146.377 79.828 ;
			RECT	146.513 79.764 146.545 79.828 ;
			RECT	146.681 79.764 146.713 79.828 ;
			RECT	146.849 79.764 146.881 79.828 ;
			RECT	147.017 79.764 147.049 79.828 ;
			RECT	147.185 79.764 147.217 79.828 ;
			RECT	147.316 79.78 147.348 79.812 ;
			RECT	147.437 79.78 147.469 79.812 ;
			RECT	147.567 79.764 147.599 79.828 ;
			RECT	149.879 79.764 149.911 79.828 ;
			RECT	151.13 79.764 151.194 79.828 ;
			RECT	151.81 79.764 151.842 79.828 ;
			RECT	152.249 79.764 152.281 79.828 ;
			RECT	153.56 79.764 153.624 79.828 ;
			RECT	156.601 79.764 156.633 79.828 ;
			RECT	156.731 79.78 156.763 79.812 ;
			RECT	156.852 79.78 156.884 79.812 ;
			RECT	156.983 79.764 157.015 79.828 ;
			RECT	157.151 79.764 157.183 79.828 ;
			RECT	157.319 79.764 157.351 79.828 ;
			RECT	157.487 79.764 157.519 79.828 ;
			RECT	157.655 79.764 157.687 79.828 ;
			RECT	157.823 79.764 157.855 79.828 ;
			RECT	157.991 79.764 158.023 79.828 ;
			RECT	158.159 79.764 158.191 79.828 ;
			RECT	158.327 79.764 158.359 79.828 ;
			RECT	158.495 79.764 158.527 79.828 ;
			RECT	158.663 79.764 158.695 79.828 ;
			RECT	158.831 79.764 158.863 79.828 ;
			RECT	158.999 79.764 159.031 79.828 ;
			RECT	159.167 79.764 159.199 79.828 ;
			RECT	159.335 79.764 159.367 79.828 ;
			RECT	159.503 79.764 159.535 79.828 ;
			RECT	159.671 79.764 159.703 79.828 ;
			RECT	159.839 79.764 159.871 79.828 ;
			RECT	160.007 79.764 160.039 79.828 ;
			RECT	160.175 79.764 160.207 79.828 ;
			RECT	160.343 79.764 160.375 79.828 ;
			RECT	160.511 79.764 160.543 79.828 ;
			RECT	160.679 79.764 160.711 79.828 ;
			RECT	160.847 79.764 160.879 79.828 ;
			RECT	161.015 79.764 161.047 79.828 ;
			RECT	161.183 79.764 161.215 79.828 ;
			RECT	161.351 79.764 161.383 79.828 ;
			RECT	161.519 79.764 161.551 79.828 ;
			RECT	161.687 79.764 161.719 79.828 ;
			RECT	161.855 79.764 161.887 79.828 ;
			RECT	162.023 79.764 162.055 79.828 ;
			RECT	162.191 79.764 162.223 79.828 ;
			RECT	162.359 79.764 162.391 79.828 ;
			RECT	162.527 79.764 162.559 79.828 ;
			RECT	162.695 79.764 162.727 79.828 ;
			RECT	162.863 79.764 162.895 79.828 ;
			RECT	163.031 79.764 163.063 79.828 ;
			RECT	163.199 79.764 163.231 79.828 ;
			RECT	163.367 79.764 163.399 79.828 ;
			RECT	163.535 79.764 163.567 79.828 ;
			RECT	163.703 79.764 163.735 79.828 ;
			RECT	163.871 79.764 163.903 79.828 ;
			RECT	164.039 79.764 164.071 79.828 ;
			RECT	164.207 79.764 164.239 79.828 ;
			RECT	164.375 79.764 164.407 79.828 ;
			RECT	164.543 79.764 164.575 79.828 ;
			RECT	164.711 79.764 164.743 79.828 ;
			RECT	164.879 79.764 164.911 79.828 ;
			RECT	165.047 79.764 165.079 79.828 ;
			RECT	165.215 79.764 165.247 79.828 ;
			RECT	165.383 79.764 165.415 79.828 ;
			RECT	165.551 79.764 165.583 79.828 ;
			RECT	165.719 79.764 165.751 79.828 ;
			RECT	165.887 79.764 165.919 79.828 ;
			RECT	166.055 79.764 166.087 79.828 ;
			RECT	166.223 79.764 166.255 79.828 ;
			RECT	166.391 79.764 166.423 79.828 ;
			RECT	166.559 79.764 166.591 79.828 ;
			RECT	166.727 79.764 166.759 79.828 ;
			RECT	166.895 79.764 166.927 79.828 ;
			RECT	167.063 79.764 167.095 79.828 ;
			RECT	167.231 79.764 167.263 79.828 ;
			RECT	167.399 79.764 167.431 79.828 ;
			RECT	167.567 79.764 167.599 79.828 ;
			RECT	167.735 79.764 167.767 79.828 ;
			RECT	167.903 79.764 167.935 79.828 ;
			RECT	168.071 79.764 168.103 79.828 ;
			RECT	168.239 79.764 168.271 79.828 ;
			RECT	168.407 79.764 168.439 79.828 ;
			RECT	168.575 79.764 168.607 79.828 ;
			RECT	168.743 79.764 168.775 79.828 ;
			RECT	168.911 79.764 168.943 79.828 ;
			RECT	169.079 79.764 169.111 79.828 ;
			RECT	169.247 79.764 169.279 79.828 ;
			RECT	169.415 79.764 169.447 79.828 ;
			RECT	169.583 79.764 169.615 79.828 ;
			RECT	169.751 79.764 169.783 79.828 ;
			RECT	169.919 79.764 169.951 79.828 ;
			RECT	170.087 79.764 170.119 79.828 ;
			RECT	170.255 79.764 170.287 79.828 ;
			RECT	170.423 79.764 170.455 79.828 ;
			RECT	170.591 79.764 170.623 79.828 ;
			RECT	170.759 79.764 170.791 79.828 ;
			RECT	170.927 79.764 170.959 79.828 ;
			RECT	171.095 79.764 171.127 79.828 ;
			RECT	171.263 79.764 171.295 79.828 ;
			RECT	171.431 79.764 171.463 79.828 ;
			RECT	171.599 79.764 171.631 79.828 ;
			RECT	171.767 79.764 171.799 79.828 ;
			RECT	171.935 79.764 171.967 79.828 ;
			RECT	172.103 79.764 172.135 79.828 ;
			RECT	172.271 79.764 172.303 79.828 ;
			RECT	172.439 79.764 172.471 79.828 ;
			RECT	172.607 79.764 172.639 79.828 ;
			RECT	172.775 79.764 172.807 79.828 ;
			RECT	172.943 79.764 172.975 79.828 ;
			RECT	173.111 79.764 173.143 79.828 ;
			RECT	173.279 79.764 173.311 79.828 ;
			RECT	173.447 79.764 173.479 79.828 ;
			RECT	173.615 79.764 173.647 79.828 ;
			RECT	173.783 79.764 173.815 79.828 ;
			RECT	173.951 79.764 173.983 79.828 ;
			RECT	174.119 79.764 174.151 79.828 ;
			RECT	174.287 79.764 174.319 79.828 ;
			RECT	174.455 79.764 174.487 79.828 ;
			RECT	174.623 79.764 174.655 79.828 ;
			RECT	174.791 79.764 174.823 79.828 ;
			RECT	174.959 79.764 174.991 79.828 ;
			RECT	175.127 79.764 175.159 79.828 ;
			RECT	175.295 79.764 175.327 79.828 ;
			RECT	175.463 79.764 175.495 79.828 ;
			RECT	175.631 79.764 175.663 79.828 ;
			RECT	175.799 79.764 175.831 79.828 ;
			RECT	175.967 79.764 175.999 79.828 ;
			RECT	176.135 79.764 176.167 79.828 ;
			RECT	176.303 79.764 176.335 79.828 ;
			RECT	176.471 79.764 176.503 79.828 ;
			RECT	176.639 79.764 176.671 79.828 ;
			RECT	176.807 79.764 176.839 79.828 ;
			RECT	176.975 79.764 177.007 79.828 ;
			RECT	177.143 79.764 177.175 79.828 ;
			RECT	177.311 79.764 177.343 79.828 ;
			RECT	177.479 79.764 177.511 79.828 ;
			RECT	177.647 79.764 177.679 79.828 ;
			RECT	177.815 79.764 177.847 79.828 ;
			RECT	177.983 79.764 178.015 79.828 ;
			RECT	178.151 79.764 178.183 79.828 ;
			RECT	178.319 79.764 178.351 79.828 ;
			RECT	178.487 79.764 178.519 79.828 ;
			RECT	178.655 79.764 178.687 79.828 ;
			RECT	178.823 79.764 178.855 79.828 ;
			RECT	178.991 79.764 179.023 79.828 ;
			RECT	179.159 79.764 179.191 79.828 ;
			RECT	179.327 79.764 179.359 79.828 ;
			RECT	179.495 79.764 179.527 79.828 ;
			RECT	179.663 79.764 179.695 79.828 ;
			RECT	179.831 79.764 179.863 79.828 ;
			RECT	179.999 79.764 180.031 79.828 ;
			RECT	180.167 79.764 180.199 79.828 ;
			RECT	180.335 79.764 180.367 79.828 ;
			RECT	180.503 79.764 180.535 79.828 ;
			RECT	180.671 79.764 180.703 79.828 ;
			RECT	180.839 79.764 180.871 79.828 ;
			RECT	181.007 79.764 181.039 79.828 ;
			RECT	181.175 79.764 181.207 79.828 ;
			RECT	181.343 79.764 181.375 79.828 ;
			RECT	181.511 79.764 181.543 79.828 ;
			RECT	181.679 79.764 181.711 79.828 ;
			RECT	181.847 79.764 181.879 79.828 ;
			RECT	182.015 79.764 182.047 79.828 ;
			RECT	182.183 79.764 182.215 79.828 ;
			RECT	182.351 79.764 182.383 79.828 ;
			RECT	182.519 79.764 182.551 79.828 ;
			RECT	182.687 79.764 182.719 79.828 ;
			RECT	182.855 79.764 182.887 79.828 ;
			RECT	183.023 79.764 183.055 79.828 ;
			RECT	183.191 79.764 183.223 79.828 ;
			RECT	183.359 79.764 183.391 79.828 ;
			RECT	183.527 79.764 183.559 79.828 ;
			RECT	183.695 79.764 183.727 79.828 ;
			RECT	183.863 79.764 183.895 79.828 ;
			RECT	184.031 79.764 184.063 79.828 ;
			RECT	184.199 79.764 184.231 79.828 ;
			RECT	184.367 79.764 184.399 79.828 ;
			RECT	184.535 79.764 184.567 79.828 ;
			RECT	184.703 79.764 184.735 79.828 ;
			RECT	184.871 79.764 184.903 79.828 ;
			RECT	185.039 79.764 185.071 79.828 ;
			RECT	185.207 79.764 185.239 79.828 ;
			RECT	185.375 79.764 185.407 79.828 ;
			RECT	185.543 79.764 185.575 79.828 ;
			RECT	185.711 79.764 185.743 79.828 ;
			RECT	185.879 79.764 185.911 79.828 ;
			RECT	186.047 79.764 186.079 79.828 ;
			RECT	186.215 79.764 186.247 79.828 ;
			RECT	186.383 79.764 186.415 79.828 ;
			RECT	186.551 79.764 186.583 79.828 ;
			RECT	186.719 79.764 186.751 79.828 ;
			RECT	186.887 79.764 186.919 79.828 ;
			RECT	187.055 79.764 187.087 79.828 ;
			RECT	187.223 79.764 187.255 79.828 ;
			RECT	187.391 79.764 187.423 79.828 ;
			RECT	187.559 79.764 187.591 79.828 ;
			RECT	187.727 79.764 187.759 79.828 ;
			RECT	187.895 79.764 187.927 79.828 ;
			RECT	188.063 79.764 188.095 79.828 ;
			RECT	188.231 79.764 188.263 79.828 ;
			RECT	188.399 79.764 188.431 79.828 ;
			RECT	188.567 79.764 188.599 79.828 ;
			RECT	188.735 79.764 188.767 79.828 ;
			RECT	188.903 79.764 188.935 79.828 ;
			RECT	189.071 79.764 189.103 79.828 ;
			RECT	189.239 79.764 189.271 79.828 ;
			RECT	189.407 79.764 189.439 79.828 ;
			RECT	189.575 79.764 189.607 79.828 ;
			RECT	189.743 79.764 189.775 79.828 ;
			RECT	189.911 79.764 189.943 79.828 ;
			RECT	190.079 79.764 190.111 79.828 ;
			RECT	190.247 79.764 190.279 79.828 ;
			RECT	190.415 79.764 190.447 79.828 ;
			RECT	190.583 79.764 190.615 79.828 ;
			RECT	190.751 79.764 190.783 79.828 ;
			RECT	190.919 79.764 190.951 79.828 ;
			RECT	191.087 79.764 191.119 79.828 ;
			RECT	191.255 79.764 191.287 79.828 ;
			RECT	191.423 79.764 191.455 79.828 ;
			RECT	191.591 79.764 191.623 79.828 ;
			RECT	191.759 79.764 191.791 79.828 ;
			RECT	191.927 79.764 191.959 79.828 ;
			RECT	192.095 79.764 192.127 79.828 ;
			RECT	192.263 79.764 192.295 79.828 ;
			RECT	192.431 79.764 192.463 79.828 ;
			RECT	192.599 79.764 192.631 79.828 ;
			RECT	192.767 79.764 192.799 79.828 ;
			RECT	192.935 79.764 192.967 79.828 ;
			RECT	193.103 79.764 193.135 79.828 ;
			RECT	193.271 79.764 193.303 79.828 ;
			RECT	193.439 79.764 193.471 79.828 ;
			RECT	193.607 79.764 193.639 79.828 ;
			RECT	193.775 79.764 193.807 79.828 ;
			RECT	193.943 79.764 193.975 79.828 ;
			RECT	194.111 79.764 194.143 79.828 ;
			RECT	194.279 79.764 194.311 79.828 ;
			RECT	194.447 79.764 194.479 79.828 ;
			RECT	194.615 79.764 194.647 79.828 ;
			RECT	194.783 79.764 194.815 79.828 ;
			RECT	194.951 79.764 194.983 79.828 ;
			RECT	195.119 79.764 195.151 79.828 ;
			RECT	195.287 79.764 195.319 79.828 ;
			RECT	195.455 79.764 195.487 79.828 ;
			RECT	195.623 79.764 195.655 79.828 ;
			RECT	195.791 79.764 195.823 79.828 ;
			RECT	195.959 79.764 195.991 79.828 ;
			RECT	196.127 79.764 196.159 79.828 ;
			RECT	196.295 79.764 196.327 79.828 ;
			RECT	196.463 79.764 196.495 79.828 ;
			RECT	196.631 79.764 196.663 79.828 ;
			RECT	196.799 79.764 196.831 79.828 ;
			RECT	196.967 79.764 196.999 79.828 ;
			RECT	197.135 79.764 197.167 79.828 ;
			RECT	197.303 79.764 197.335 79.828 ;
			RECT	197.471 79.764 197.503 79.828 ;
			RECT	197.639 79.764 197.671 79.828 ;
			RECT	197.807 79.764 197.839 79.828 ;
			RECT	197.975 79.764 198.007 79.828 ;
			RECT	198.143 79.764 198.175 79.828 ;
			RECT	198.311 79.764 198.343 79.828 ;
			RECT	198.479 79.764 198.511 79.828 ;
			RECT	198.647 79.764 198.679 79.828 ;
			RECT	198.815 79.764 198.847 79.828 ;
			RECT	198.983 79.764 199.015 79.828 ;
			RECT	199.151 79.764 199.183 79.828 ;
			RECT	199.319 79.764 199.351 79.828 ;
			RECT	199.487 79.764 199.519 79.828 ;
			RECT	199.655 79.764 199.687 79.828 ;
			RECT	199.823 79.764 199.855 79.828 ;
			RECT	199.991 79.764 200.023 79.828 ;
			RECT	200.121 79.78 200.153 79.812 ;
			RECT	200.243 79.775 200.275 79.807 ;
			RECT	200.373 79.764 200.405 79.828 ;
			RECT	200.9 79.764 200.932 79.828 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 31.12 201.665 31.24 ;
			LAYER	J3 ;
			RECT	0.755 31.148 0.787 31.212 ;
			RECT	1.645 31.148 1.709 31.212 ;
			RECT	2.323 31.148 2.387 31.212 ;
			RECT	3.438 31.148 3.47 31.212 ;
			RECT	3.585 31.148 3.617 31.212 ;
			RECT	4.195 31.148 4.227 31.212 ;
			RECT	4.72 31.148 4.752 31.212 ;
			RECT	4.944 31.148 5.008 31.212 ;
			RECT	5.267 31.148 5.299 31.212 ;
			RECT	5.797 31.148 5.829 31.212 ;
			RECT	5.927 31.169 5.959 31.201 ;
			RECT	6.049 31.164 6.081 31.196 ;
			RECT	6.179 31.148 6.211 31.212 ;
			RECT	6.347 31.148 6.379 31.212 ;
			RECT	6.515 31.148 6.547 31.212 ;
			RECT	6.683 31.148 6.715 31.212 ;
			RECT	6.851 31.148 6.883 31.212 ;
			RECT	7.019 31.148 7.051 31.212 ;
			RECT	7.187 31.148 7.219 31.212 ;
			RECT	7.355 31.148 7.387 31.212 ;
			RECT	7.523 31.148 7.555 31.212 ;
			RECT	7.691 31.148 7.723 31.212 ;
			RECT	7.859 31.148 7.891 31.212 ;
			RECT	8.027 31.148 8.059 31.212 ;
			RECT	8.195 31.148 8.227 31.212 ;
			RECT	8.363 31.148 8.395 31.212 ;
			RECT	8.531 31.148 8.563 31.212 ;
			RECT	8.699 31.148 8.731 31.212 ;
			RECT	8.867 31.148 8.899 31.212 ;
			RECT	9.035 31.148 9.067 31.212 ;
			RECT	9.203 31.148 9.235 31.212 ;
			RECT	9.371 31.148 9.403 31.212 ;
			RECT	9.539 31.148 9.571 31.212 ;
			RECT	9.707 31.148 9.739 31.212 ;
			RECT	9.875 31.148 9.907 31.212 ;
			RECT	10.043 31.148 10.075 31.212 ;
			RECT	10.211 31.148 10.243 31.212 ;
			RECT	10.379 31.148 10.411 31.212 ;
			RECT	10.547 31.148 10.579 31.212 ;
			RECT	10.715 31.148 10.747 31.212 ;
			RECT	10.883 31.148 10.915 31.212 ;
			RECT	11.051 31.148 11.083 31.212 ;
			RECT	11.219 31.148 11.251 31.212 ;
			RECT	11.387 31.148 11.419 31.212 ;
			RECT	11.555 31.148 11.587 31.212 ;
			RECT	11.723 31.148 11.755 31.212 ;
			RECT	11.891 31.148 11.923 31.212 ;
			RECT	12.059 31.148 12.091 31.212 ;
			RECT	12.227 31.148 12.259 31.212 ;
			RECT	12.395 31.148 12.427 31.212 ;
			RECT	12.563 31.148 12.595 31.212 ;
			RECT	12.731 31.148 12.763 31.212 ;
			RECT	12.899 31.148 12.931 31.212 ;
			RECT	13.067 31.148 13.099 31.212 ;
			RECT	13.235 31.148 13.267 31.212 ;
			RECT	13.403 31.148 13.435 31.212 ;
			RECT	13.571 31.148 13.603 31.212 ;
			RECT	13.739 31.148 13.771 31.212 ;
			RECT	13.907 31.148 13.939 31.212 ;
			RECT	14.075 31.148 14.107 31.212 ;
			RECT	14.243 31.148 14.275 31.212 ;
			RECT	14.411 31.148 14.443 31.212 ;
			RECT	14.579 31.148 14.611 31.212 ;
			RECT	14.747 31.148 14.779 31.212 ;
			RECT	14.915 31.148 14.947 31.212 ;
			RECT	15.083 31.148 15.115 31.212 ;
			RECT	15.251 31.148 15.283 31.212 ;
			RECT	15.419 31.148 15.451 31.212 ;
			RECT	15.587 31.148 15.619 31.212 ;
			RECT	15.755 31.148 15.787 31.212 ;
			RECT	15.923 31.148 15.955 31.212 ;
			RECT	16.091 31.148 16.123 31.212 ;
			RECT	16.259 31.148 16.291 31.212 ;
			RECT	16.427 31.148 16.459 31.212 ;
			RECT	16.595 31.148 16.627 31.212 ;
			RECT	16.763 31.148 16.795 31.212 ;
			RECT	16.931 31.148 16.963 31.212 ;
			RECT	17.099 31.148 17.131 31.212 ;
			RECT	17.267 31.148 17.299 31.212 ;
			RECT	17.435 31.148 17.467 31.212 ;
			RECT	17.603 31.148 17.635 31.212 ;
			RECT	17.771 31.148 17.803 31.212 ;
			RECT	17.939 31.148 17.971 31.212 ;
			RECT	18.107 31.148 18.139 31.212 ;
			RECT	18.275 31.148 18.307 31.212 ;
			RECT	18.443 31.148 18.475 31.212 ;
			RECT	18.611 31.148 18.643 31.212 ;
			RECT	18.779 31.148 18.811 31.212 ;
			RECT	18.947 31.148 18.979 31.212 ;
			RECT	19.115 31.148 19.147 31.212 ;
			RECT	19.283 31.148 19.315 31.212 ;
			RECT	19.451 31.148 19.483 31.212 ;
			RECT	19.619 31.148 19.651 31.212 ;
			RECT	19.787 31.148 19.819 31.212 ;
			RECT	19.955 31.148 19.987 31.212 ;
			RECT	20.123 31.148 20.155 31.212 ;
			RECT	20.291 31.148 20.323 31.212 ;
			RECT	20.459 31.148 20.491 31.212 ;
			RECT	20.627 31.148 20.659 31.212 ;
			RECT	20.795 31.148 20.827 31.212 ;
			RECT	20.963 31.148 20.995 31.212 ;
			RECT	21.131 31.148 21.163 31.212 ;
			RECT	21.299 31.148 21.331 31.212 ;
			RECT	21.467 31.148 21.499 31.212 ;
			RECT	21.635 31.148 21.667 31.212 ;
			RECT	21.803 31.148 21.835 31.212 ;
			RECT	21.971 31.148 22.003 31.212 ;
			RECT	22.139 31.148 22.171 31.212 ;
			RECT	22.307 31.148 22.339 31.212 ;
			RECT	22.475 31.148 22.507 31.212 ;
			RECT	22.643 31.148 22.675 31.212 ;
			RECT	22.811 31.148 22.843 31.212 ;
			RECT	22.979 31.148 23.011 31.212 ;
			RECT	23.147 31.148 23.179 31.212 ;
			RECT	23.315 31.148 23.347 31.212 ;
			RECT	23.483 31.148 23.515 31.212 ;
			RECT	23.651 31.148 23.683 31.212 ;
			RECT	23.819 31.148 23.851 31.212 ;
			RECT	23.987 31.148 24.019 31.212 ;
			RECT	24.155 31.148 24.187 31.212 ;
			RECT	24.323 31.148 24.355 31.212 ;
			RECT	24.491 31.148 24.523 31.212 ;
			RECT	24.659 31.148 24.691 31.212 ;
			RECT	24.827 31.148 24.859 31.212 ;
			RECT	24.995 31.148 25.027 31.212 ;
			RECT	25.163 31.148 25.195 31.212 ;
			RECT	25.331 31.148 25.363 31.212 ;
			RECT	25.499 31.148 25.531 31.212 ;
			RECT	25.667 31.148 25.699 31.212 ;
			RECT	25.835 31.148 25.867 31.212 ;
			RECT	26.003 31.148 26.035 31.212 ;
			RECT	26.171 31.148 26.203 31.212 ;
			RECT	26.339 31.148 26.371 31.212 ;
			RECT	26.507 31.148 26.539 31.212 ;
			RECT	26.675 31.148 26.707 31.212 ;
			RECT	26.843 31.148 26.875 31.212 ;
			RECT	27.011 31.148 27.043 31.212 ;
			RECT	27.179 31.148 27.211 31.212 ;
			RECT	27.347 31.148 27.379 31.212 ;
			RECT	27.515 31.148 27.547 31.212 ;
			RECT	27.683 31.148 27.715 31.212 ;
			RECT	27.851 31.148 27.883 31.212 ;
			RECT	28.019 31.148 28.051 31.212 ;
			RECT	28.187 31.148 28.219 31.212 ;
			RECT	28.355 31.148 28.387 31.212 ;
			RECT	28.523 31.148 28.555 31.212 ;
			RECT	28.691 31.148 28.723 31.212 ;
			RECT	28.859 31.148 28.891 31.212 ;
			RECT	29.027 31.148 29.059 31.212 ;
			RECT	29.195 31.148 29.227 31.212 ;
			RECT	29.363 31.148 29.395 31.212 ;
			RECT	29.531 31.148 29.563 31.212 ;
			RECT	29.699 31.148 29.731 31.212 ;
			RECT	29.867 31.148 29.899 31.212 ;
			RECT	30.035 31.148 30.067 31.212 ;
			RECT	30.203 31.148 30.235 31.212 ;
			RECT	30.371 31.148 30.403 31.212 ;
			RECT	30.539 31.148 30.571 31.212 ;
			RECT	30.707 31.148 30.739 31.212 ;
			RECT	30.875 31.148 30.907 31.212 ;
			RECT	31.043 31.148 31.075 31.212 ;
			RECT	31.211 31.148 31.243 31.212 ;
			RECT	31.379 31.148 31.411 31.212 ;
			RECT	31.547 31.148 31.579 31.212 ;
			RECT	31.715 31.148 31.747 31.212 ;
			RECT	31.883 31.148 31.915 31.212 ;
			RECT	32.051 31.148 32.083 31.212 ;
			RECT	32.219 31.148 32.251 31.212 ;
			RECT	32.387 31.148 32.419 31.212 ;
			RECT	32.555 31.148 32.587 31.212 ;
			RECT	32.723 31.148 32.755 31.212 ;
			RECT	32.891 31.148 32.923 31.212 ;
			RECT	33.059 31.148 33.091 31.212 ;
			RECT	33.227 31.148 33.259 31.212 ;
			RECT	33.395 31.148 33.427 31.212 ;
			RECT	33.563 31.148 33.595 31.212 ;
			RECT	33.731 31.148 33.763 31.212 ;
			RECT	33.899 31.148 33.931 31.212 ;
			RECT	34.067 31.148 34.099 31.212 ;
			RECT	34.235 31.148 34.267 31.212 ;
			RECT	34.403 31.148 34.435 31.212 ;
			RECT	34.571 31.148 34.603 31.212 ;
			RECT	34.739 31.148 34.771 31.212 ;
			RECT	34.907 31.148 34.939 31.212 ;
			RECT	35.075 31.148 35.107 31.212 ;
			RECT	35.243 31.148 35.275 31.212 ;
			RECT	35.411 31.148 35.443 31.212 ;
			RECT	35.579 31.148 35.611 31.212 ;
			RECT	35.747 31.148 35.779 31.212 ;
			RECT	35.915 31.148 35.947 31.212 ;
			RECT	36.083 31.148 36.115 31.212 ;
			RECT	36.251 31.148 36.283 31.212 ;
			RECT	36.419 31.148 36.451 31.212 ;
			RECT	36.587 31.148 36.619 31.212 ;
			RECT	36.755 31.148 36.787 31.212 ;
			RECT	36.923 31.148 36.955 31.212 ;
			RECT	37.091 31.148 37.123 31.212 ;
			RECT	37.259 31.148 37.291 31.212 ;
			RECT	37.427 31.148 37.459 31.212 ;
			RECT	37.595 31.148 37.627 31.212 ;
			RECT	37.763 31.148 37.795 31.212 ;
			RECT	37.931 31.148 37.963 31.212 ;
			RECT	38.099 31.148 38.131 31.212 ;
			RECT	38.267 31.148 38.299 31.212 ;
			RECT	38.435 31.148 38.467 31.212 ;
			RECT	38.603 31.148 38.635 31.212 ;
			RECT	38.771 31.148 38.803 31.212 ;
			RECT	38.939 31.148 38.971 31.212 ;
			RECT	39.107 31.148 39.139 31.212 ;
			RECT	39.275 31.148 39.307 31.212 ;
			RECT	39.443 31.148 39.475 31.212 ;
			RECT	39.611 31.148 39.643 31.212 ;
			RECT	39.779 31.148 39.811 31.212 ;
			RECT	39.947 31.148 39.979 31.212 ;
			RECT	40.115 31.148 40.147 31.212 ;
			RECT	40.283 31.148 40.315 31.212 ;
			RECT	40.451 31.148 40.483 31.212 ;
			RECT	40.619 31.148 40.651 31.212 ;
			RECT	40.787 31.148 40.819 31.212 ;
			RECT	40.955 31.148 40.987 31.212 ;
			RECT	41.123 31.148 41.155 31.212 ;
			RECT	41.291 31.148 41.323 31.212 ;
			RECT	41.459 31.148 41.491 31.212 ;
			RECT	41.627 31.148 41.659 31.212 ;
			RECT	41.795 31.148 41.827 31.212 ;
			RECT	41.963 31.148 41.995 31.212 ;
			RECT	42.131 31.148 42.163 31.212 ;
			RECT	42.299 31.148 42.331 31.212 ;
			RECT	42.467 31.148 42.499 31.212 ;
			RECT	42.635 31.148 42.667 31.212 ;
			RECT	42.803 31.148 42.835 31.212 ;
			RECT	42.971 31.148 43.003 31.212 ;
			RECT	43.139 31.148 43.171 31.212 ;
			RECT	43.307 31.148 43.339 31.212 ;
			RECT	43.475 31.148 43.507 31.212 ;
			RECT	43.643 31.148 43.675 31.212 ;
			RECT	43.811 31.148 43.843 31.212 ;
			RECT	43.979 31.148 44.011 31.212 ;
			RECT	44.147 31.148 44.179 31.212 ;
			RECT	44.315 31.148 44.347 31.212 ;
			RECT	44.483 31.148 44.515 31.212 ;
			RECT	44.651 31.148 44.683 31.212 ;
			RECT	44.819 31.148 44.851 31.212 ;
			RECT	44.987 31.148 45.019 31.212 ;
			RECT	45.155 31.148 45.187 31.212 ;
			RECT	45.323 31.148 45.355 31.212 ;
			RECT	45.491 31.148 45.523 31.212 ;
			RECT	45.659 31.148 45.691 31.212 ;
			RECT	45.827 31.148 45.859 31.212 ;
			RECT	45.995 31.148 46.027 31.212 ;
			RECT	46.163 31.148 46.195 31.212 ;
			RECT	46.331 31.148 46.363 31.212 ;
			RECT	46.499 31.148 46.531 31.212 ;
			RECT	46.667 31.148 46.699 31.212 ;
			RECT	46.835 31.148 46.867 31.212 ;
			RECT	47.003 31.148 47.035 31.212 ;
			RECT	47.171 31.148 47.203 31.212 ;
			RECT	47.339 31.148 47.371 31.212 ;
			RECT	47.507 31.148 47.539 31.212 ;
			RECT	47.675 31.148 47.707 31.212 ;
			RECT	47.843 31.148 47.875 31.212 ;
			RECT	48.011 31.148 48.043 31.212 ;
			RECT	48.179 31.148 48.211 31.212 ;
			RECT	48.347 31.148 48.379 31.212 ;
			RECT	48.515 31.148 48.547 31.212 ;
			RECT	48.683 31.148 48.715 31.212 ;
			RECT	48.851 31.148 48.883 31.212 ;
			RECT	49.019 31.148 49.051 31.212 ;
			RECT	49.187 31.148 49.219 31.212 ;
			RECT	49.318 31.164 49.35 31.196 ;
			RECT	49.439 31.164 49.471 31.196 ;
			RECT	49.569 31.148 49.601 31.212 ;
			RECT	51.881 31.148 51.913 31.212 ;
			RECT	53.132 31.148 53.196 31.212 ;
			RECT	53.812 31.148 53.844 31.212 ;
			RECT	54.251 31.148 54.283 31.212 ;
			RECT	55.562 31.148 55.626 31.212 ;
			RECT	58.603 31.148 58.635 31.212 ;
			RECT	58.733 31.164 58.765 31.196 ;
			RECT	58.854 31.164 58.886 31.196 ;
			RECT	58.985 31.148 59.017 31.212 ;
			RECT	59.153 31.148 59.185 31.212 ;
			RECT	59.321 31.148 59.353 31.212 ;
			RECT	59.489 31.148 59.521 31.212 ;
			RECT	59.657 31.148 59.689 31.212 ;
			RECT	59.825 31.148 59.857 31.212 ;
			RECT	59.993 31.148 60.025 31.212 ;
			RECT	60.161 31.148 60.193 31.212 ;
			RECT	60.329 31.148 60.361 31.212 ;
			RECT	60.497 31.148 60.529 31.212 ;
			RECT	60.665 31.148 60.697 31.212 ;
			RECT	60.833 31.148 60.865 31.212 ;
			RECT	61.001 31.148 61.033 31.212 ;
			RECT	61.169 31.148 61.201 31.212 ;
			RECT	61.337 31.148 61.369 31.212 ;
			RECT	61.505 31.148 61.537 31.212 ;
			RECT	61.673 31.148 61.705 31.212 ;
			RECT	61.841 31.148 61.873 31.212 ;
			RECT	62.009 31.148 62.041 31.212 ;
			RECT	62.177 31.148 62.209 31.212 ;
			RECT	62.345 31.148 62.377 31.212 ;
			RECT	62.513 31.148 62.545 31.212 ;
			RECT	62.681 31.148 62.713 31.212 ;
			RECT	62.849 31.148 62.881 31.212 ;
			RECT	63.017 31.148 63.049 31.212 ;
			RECT	63.185 31.148 63.217 31.212 ;
			RECT	63.353 31.148 63.385 31.212 ;
			RECT	63.521 31.148 63.553 31.212 ;
			RECT	63.689 31.148 63.721 31.212 ;
			RECT	63.857 31.148 63.889 31.212 ;
			RECT	64.025 31.148 64.057 31.212 ;
			RECT	64.193 31.148 64.225 31.212 ;
			RECT	64.361 31.148 64.393 31.212 ;
			RECT	64.529 31.148 64.561 31.212 ;
			RECT	64.697 31.148 64.729 31.212 ;
			RECT	64.865 31.148 64.897 31.212 ;
			RECT	65.033 31.148 65.065 31.212 ;
			RECT	65.201 31.148 65.233 31.212 ;
			RECT	65.369 31.148 65.401 31.212 ;
			RECT	65.537 31.148 65.569 31.212 ;
			RECT	65.705 31.148 65.737 31.212 ;
			RECT	65.873 31.148 65.905 31.212 ;
			RECT	66.041 31.148 66.073 31.212 ;
			RECT	66.209 31.148 66.241 31.212 ;
			RECT	66.377 31.148 66.409 31.212 ;
			RECT	66.545 31.148 66.577 31.212 ;
			RECT	66.713 31.148 66.745 31.212 ;
			RECT	66.881 31.148 66.913 31.212 ;
			RECT	67.049 31.148 67.081 31.212 ;
			RECT	67.217 31.148 67.249 31.212 ;
			RECT	67.385 31.148 67.417 31.212 ;
			RECT	67.553 31.148 67.585 31.212 ;
			RECT	67.721 31.148 67.753 31.212 ;
			RECT	67.889 31.148 67.921 31.212 ;
			RECT	68.057 31.148 68.089 31.212 ;
			RECT	68.225 31.148 68.257 31.212 ;
			RECT	68.393 31.148 68.425 31.212 ;
			RECT	68.561 31.148 68.593 31.212 ;
			RECT	68.729 31.148 68.761 31.212 ;
			RECT	68.897 31.148 68.929 31.212 ;
			RECT	69.065 31.148 69.097 31.212 ;
			RECT	69.233 31.148 69.265 31.212 ;
			RECT	69.401 31.148 69.433 31.212 ;
			RECT	69.569 31.148 69.601 31.212 ;
			RECT	69.737 31.148 69.769 31.212 ;
			RECT	69.905 31.148 69.937 31.212 ;
			RECT	70.073 31.148 70.105 31.212 ;
			RECT	70.241 31.148 70.273 31.212 ;
			RECT	70.409 31.148 70.441 31.212 ;
			RECT	70.577 31.148 70.609 31.212 ;
			RECT	70.745 31.148 70.777 31.212 ;
			RECT	70.913 31.148 70.945 31.212 ;
			RECT	71.081 31.148 71.113 31.212 ;
			RECT	71.249 31.148 71.281 31.212 ;
			RECT	71.417 31.148 71.449 31.212 ;
			RECT	71.585 31.148 71.617 31.212 ;
			RECT	71.753 31.148 71.785 31.212 ;
			RECT	71.921 31.148 71.953 31.212 ;
			RECT	72.089 31.148 72.121 31.212 ;
			RECT	72.257 31.148 72.289 31.212 ;
			RECT	72.425 31.148 72.457 31.212 ;
			RECT	72.593 31.148 72.625 31.212 ;
			RECT	72.761 31.148 72.793 31.212 ;
			RECT	72.929 31.148 72.961 31.212 ;
			RECT	73.097 31.148 73.129 31.212 ;
			RECT	73.265 31.148 73.297 31.212 ;
			RECT	73.433 31.148 73.465 31.212 ;
			RECT	73.601 31.148 73.633 31.212 ;
			RECT	73.769 31.148 73.801 31.212 ;
			RECT	73.937 31.148 73.969 31.212 ;
			RECT	74.105 31.148 74.137 31.212 ;
			RECT	74.273 31.148 74.305 31.212 ;
			RECT	74.441 31.148 74.473 31.212 ;
			RECT	74.609 31.148 74.641 31.212 ;
			RECT	74.777 31.148 74.809 31.212 ;
			RECT	74.945 31.148 74.977 31.212 ;
			RECT	75.113 31.148 75.145 31.212 ;
			RECT	75.281 31.148 75.313 31.212 ;
			RECT	75.449 31.148 75.481 31.212 ;
			RECT	75.617 31.148 75.649 31.212 ;
			RECT	75.785 31.148 75.817 31.212 ;
			RECT	75.953 31.148 75.985 31.212 ;
			RECT	76.121 31.148 76.153 31.212 ;
			RECT	76.289 31.148 76.321 31.212 ;
			RECT	76.457 31.148 76.489 31.212 ;
			RECT	76.625 31.148 76.657 31.212 ;
			RECT	76.793 31.148 76.825 31.212 ;
			RECT	76.961 31.148 76.993 31.212 ;
			RECT	77.129 31.148 77.161 31.212 ;
			RECT	77.297 31.148 77.329 31.212 ;
			RECT	77.465 31.148 77.497 31.212 ;
			RECT	77.633 31.148 77.665 31.212 ;
			RECT	77.801 31.148 77.833 31.212 ;
			RECT	77.969 31.148 78.001 31.212 ;
			RECT	78.137 31.148 78.169 31.212 ;
			RECT	78.305 31.148 78.337 31.212 ;
			RECT	78.473 31.148 78.505 31.212 ;
			RECT	78.641 31.148 78.673 31.212 ;
			RECT	78.809 31.148 78.841 31.212 ;
			RECT	78.977 31.148 79.009 31.212 ;
			RECT	79.145 31.148 79.177 31.212 ;
			RECT	79.313 31.148 79.345 31.212 ;
			RECT	79.481 31.148 79.513 31.212 ;
			RECT	79.649 31.148 79.681 31.212 ;
			RECT	79.817 31.148 79.849 31.212 ;
			RECT	79.985 31.148 80.017 31.212 ;
			RECT	80.153 31.148 80.185 31.212 ;
			RECT	80.321 31.148 80.353 31.212 ;
			RECT	80.489 31.148 80.521 31.212 ;
			RECT	80.657 31.148 80.689 31.212 ;
			RECT	80.825 31.148 80.857 31.212 ;
			RECT	80.993 31.148 81.025 31.212 ;
			RECT	81.161 31.148 81.193 31.212 ;
			RECT	81.329 31.148 81.361 31.212 ;
			RECT	81.497 31.148 81.529 31.212 ;
			RECT	81.665 31.148 81.697 31.212 ;
			RECT	81.833 31.148 81.865 31.212 ;
			RECT	82.001 31.148 82.033 31.212 ;
			RECT	82.169 31.148 82.201 31.212 ;
			RECT	82.337 31.148 82.369 31.212 ;
			RECT	82.505 31.148 82.537 31.212 ;
			RECT	82.673 31.148 82.705 31.212 ;
			RECT	82.841 31.148 82.873 31.212 ;
			RECT	83.009 31.148 83.041 31.212 ;
			RECT	83.177 31.148 83.209 31.212 ;
			RECT	83.345 31.148 83.377 31.212 ;
			RECT	83.513 31.148 83.545 31.212 ;
			RECT	83.681 31.148 83.713 31.212 ;
			RECT	83.849 31.148 83.881 31.212 ;
			RECT	84.017 31.148 84.049 31.212 ;
			RECT	84.185 31.148 84.217 31.212 ;
			RECT	84.353 31.148 84.385 31.212 ;
			RECT	84.521 31.148 84.553 31.212 ;
			RECT	84.689 31.148 84.721 31.212 ;
			RECT	84.857 31.148 84.889 31.212 ;
			RECT	85.025 31.148 85.057 31.212 ;
			RECT	85.193 31.148 85.225 31.212 ;
			RECT	85.361 31.148 85.393 31.212 ;
			RECT	85.529 31.148 85.561 31.212 ;
			RECT	85.697 31.148 85.729 31.212 ;
			RECT	85.865 31.148 85.897 31.212 ;
			RECT	86.033 31.148 86.065 31.212 ;
			RECT	86.201 31.148 86.233 31.212 ;
			RECT	86.369 31.148 86.401 31.212 ;
			RECT	86.537 31.148 86.569 31.212 ;
			RECT	86.705 31.148 86.737 31.212 ;
			RECT	86.873 31.148 86.905 31.212 ;
			RECT	87.041 31.148 87.073 31.212 ;
			RECT	87.209 31.148 87.241 31.212 ;
			RECT	87.377 31.148 87.409 31.212 ;
			RECT	87.545 31.148 87.577 31.212 ;
			RECT	87.713 31.148 87.745 31.212 ;
			RECT	87.881 31.148 87.913 31.212 ;
			RECT	88.049 31.148 88.081 31.212 ;
			RECT	88.217 31.148 88.249 31.212 ;
			RECT	88.385 31.148 88.417 31.212 ;
			RECT	88.553 31.148 88.585 31.212 ;
			RECT	88.721 31.148 88.753 31.212 ;
			RECT	88.889 31.148 88.921 31.212 ;
			RECT	89.057 31.148 89.089 31.212 ;
			RECT	89.225 31.148 89.257 31.212 ;
			RECT	89.393 31.148 89.425 31.212 ;
			RECT	89.561 31.148 89.593 31.212 ;
			RECT	89.729 31.148 89.761 31.212 ;
			RECT	89.897 31.148 89.929 31.212 ;
			RECT	90.065 31.148 90.097 31.212 ;
			RECT	90.233 31.148 90.265 31.212 ;
			RECT	90.401 31.148 90.433 31.212 ;
			RECT	90.569 31.148 90.601 31.212 ;
			RECT	90.737 31.148 90.769 31.212 ;
			RECT	90.905 31.148 90.937 31.212 ;
			RECT	91.073 31.148 91.105 31.212 ;
			RECT	91.241 31.148 91.273 31.212 ;
			RECT	91.409 31.148 91.441 31.212 ;
			RECT	91.577 31.148 91.609 31.212 ;
			RECT	91.745 31.148 91.777 31.212 ;
			RECT	91.913 31.148 91.945 31.212 ;
			RECT	92.081 31.148 92.113 31.212 ;
			RECT	92.249 31.148 92.281 31.212 ;
			RECT	92.417 31.148 92.449 31.212 ;
			RECT	92.585 31.148 92.617 31.212 ;
			RECT	92.753 31.148 92.785 31.212 ;
			RECT	92.921 31.148 92.953 31.212 ;
			RECT	93.089 31.148 93.121 31.212 ;
			RECT	93.257 31.148 93.289 31.212 ;
			RECT	93.425 31.148 93.457 31.212 ;
			RECT	93.593 31.148 93.625 31.212 ;
			RECT	93.761 31.148 93.793 31.212 ;
			RECT	93.929 31.148 93.961 31.212 ;
			RECT	94.097 31.148 94.129 31.212 ;
			RECT	94.265 31.148 94.297 31.212 ;
			RECT	94.433 31.148 94.465 31.212 ;
			RECT	94.601 31.148 94.633 31.212 ;
			RECT	94.769 31.148 94.801 31.212 ;
			RECT	94.937 31.148 94.969 31.212 ;
			RECT	95.105 31.148 95.137 31.212 ;
			RECT	95.273 31.148 95.305 31.212 ;
			RECT	95.441 31.148 95.473 31.212 ;
			RECT	95.609 31.148 95.641 31.212 ;
			RECT	95.777 31.148 95.809 31.212 ;
			RECT	95.945 31.148 95.977 31.212 ;
			RECT	96.113 31.148 96.145 31.212 ;
			RECT	96.281 31.148 96.313 31.212 ;
			RECT	96.449 31.148 96.481 31.212 ;
			RECT	96.617 31.148 96.649 31.212 ;
			RECT	96.785 31.148 96.817 31.212 ;
			RECT	96.953 31.148 96.985 31.212 ;
			RECT	97.121 31.148 97.153 31.212 ;
			RECT	97.289 31.148 97.321 31.212 ;
			RECT	97.457 31.148 97.489 31.212 ;
			RECT	97.625 31.148 97.657 31.212 ;
			RECT	97.793 31.148 97.825 31.212 ;
			RECT	97.961 31.148 97.993 31.212 ;
			RECT	98.129 31.148 98.161 31.212 ;
			RECT	98.297 31.148 98.329 31.212 ;
			RECT	98.465 31.148 98.497 31.212 ;
			RECT	98.633 31.148 98.665 31.212 ;
			RECT	98.801 31.148 98.833 31.212 ;
			RECT	98.969 31.148 99.001 31.212 ;
			RECT	99.137 31.148 99.169 31.212 ;
			RECT	99.305 31.148 99.337 31.212 ;
			RECT	99.473 31.148 99.505 31.212 ;
			RECT	99.641 31.148 99.673 31.212 ;
			RECT	99.809 31.148 99.841 31.212 ;
			RECT	99.977 31.148 100.009 31.212 ;
			RECT	100.145 31.148 100.177 31.212 ;
			RECT	100.313 31.148 100.345 31.212 ;
			RECT	100.481 31.148 100.513 31.212 ;
			RECT	100.649 31.148 100.681 31.212 ;
			RECT	100.817 31.148 100.849 31.212 ;
			RECT	100.985 31.148 101.017 31.212 ;
			RECT	101.153 31.148 101.185 31.212 ;
			RECT	101.321 31.148 101.353 31.212 ;
			RECT	101.489 31.148 101.521 31.212 ;
			RECT	101.657 31.148 101.689 31.212 ;
			RECT	101.825 31.148 101.857 31.212 ;
			RECT	101.993 31.148 102.025 31.212 ;
			RECT	102.123 31.164 102.155 31.196 ;
			RECT	102.245 31.169 102.277 31.201 ;
			RECT	102.375 31.148 102.407 31.212 ;
			RECT	103.795 31.148 103.827 31.212 ;
			RECT	103.925 31.169 103.957 31.201 ;
			RECT	104.047 31.164 104.079 31.196 ;
			RECT	104.177 31.148 104.209 31.212 ;
			RECT	104.345 31.148 104.377 31.212 ;
			RECT	104.513 31.148 104.545 31.212 ;
			RECT	104.681 31.148 104.713 31.212 ;
			RECT	104.849 31.148 104.881 31.212 ;
			RECT	105.017 31.148 105.049 31.212 ;
			RECT	105.185 31.148 105.217 31.212 ;
			RECT	105.353 31.148 105.385 31.212 ;
			RECT	105.521 31.148 105.553 31.212 ;
			RECT	105.689 31.148 105.721 31.212 ;
			RECT	105.857 31.148 105.889 31.212 ;
			RECT	106.025 31.148 106.057 31.212 ;
			RECT	106.193 31.148 106.225 31.212 ;
			RECT	106.361 31.148 106.393 31.212 ;
			RECT	106.529 31.148 106.561 31.212 ;
			RECT	106.697 31.148 106.729 31.212 ;
			RECT	106.865 31.148 106.897 31.212 ;
			RECT	107.033 31.148 107.065 31.212 ;
			RECT	107.201 31.148 107.233 31.212 ;
			RECT	107.369 31.148 107.401 31.212 ;
			RECT	107.537 31.148 107.569 31.212 ;
			RECT	107.705 31.148 107.737 31.212 ;
			RECT	107.873 31.148 107.905 31.212 ;
			RECT	108.041 31.148 108.073 31.212 ;
			RECT	108.209 31.148 108.241 31.212 ;
			RECT	108.377 31.148 108.409 31.212 ;
			RECT	108.545 31.148 108.577 31.212 ;
			RECT	108.713 31.148 108.745 31.212 ;
			RECT	108.881 31.148 108.913 31.212 ;
			RECT	109.049 31.148 109.081 31.212 ;
			RECT	109.217 31.148 109.249 31.212 ;
			RECT	109.385 31.148 109.417 31.212 ;
			RECT	109.553 31.148 109.585 31.212 ;
			RECT	109.721 31.148 109.753 31.212 ;
			RECT	109.889 31.148 109.921 31.212 ;
			RECT	110.057 31.148 110.089 31.212 ;
			RECT	110.225 31.148 110.257 31.212 ;
			RECT	110.393 31.148 110.425 31.212 ;
			RECT	110.561 31.148 110.593 31.212 ;
			RECT	110.729 31.148 110.761 31.212 ;
			RECT	110.897 31.148 110.929 31.212 ;
			RECT	111.065 31.148 111.097 31.212 ;
			RECT	111.233 31.148 111.265 31.212 ;
			RECT	111.401 31.148 111.433 31.212 ;
			RECT	111.569 31.148 111.601 31.212 ;
			RECT	111.737 31.148 111.769 31.212 ;
			RECT	111.905 31.148 111.937 31.212 ;
			RECT	112.073 31.148 112.105 31.212 ;
			RECT	112.241 31.148 112.273 31.212 ;
			RECT	112.409 31.148 112.441 31.212 ;
			RECT	112.577 31.148 112.609 31.212 ;
			RECT	112.745 31.148 112.777 31.212 ;
			RECT	112.913 31.148 112.945 31.212 ;
			RECT	113.081 31.148 113.113 31.212 ;
			RECT	113.249 31.148 113.281 31.212 ;
			RECT	113.417 31.148 113.449 31.212 ;
			RECT	113.585 31.148 113.617 31.212 ;
			RECT	113.753 31.148 113.785 31.212 ;
			RECT	113.921 31.148 113.953 31.212 ;
			RECT	114.089 31.148 114.121 31.212 ;
			RECT	114.257 31.148 114.289 31.212 ;
			RECT	114.425 31.148 114.457 31.212 ;
			RECT	114.593 31.148 114.625 31.212 ;
			RECT	114.761 31.148 114.793 31.212 ;
			RECT	114.929 31.148 114.961 31.212 ;
			RECT	115.097 31.148 115.129 31.212 ;
			RECT	115.265 31.148 115.297 31.212 ;
			RECT	115.433 31.148 115.465 31.212 ;
			RECT	115.601 31.148 115.633 31.212 ;
			RECT	115.769 31.148 115.801 31.212 ;
			RECT	115.937 31.148 115.969 31.212 ;
			RECT	116.105 31.148 116.137 31.212 ;
			RECT	116.273 31.148 116.305 31.212 ;
			RECT	116.441 31.148 116.473 31.212 ;
			RECT	116.609 31.148 116.641 31.212 ;
			RECT	116.777 31.148 116.809 31.212 ;
			RECT	116.945 31.148 116.977 31.212 ;
			RECT	117.113 31.148 117.145 31.212 ;
			RECT	117.281 31.148 117.313 31.212 ;
			RECT	117.449 31.148 117.481 31.212 ;
			RECT	117.617 31.148 117.649 31.212 ;
			RECT	117.785 31.148 117.817 31.212 ;
			RECT	117.953 31.148 117.985 31.212 ;
			RECT	118.121 31.148 118.153 31.212 ;
			RECT	118.289 31.148 118.321 31.212 ;
			RECT	118.457 31.148 118.489 31.212 ;
			RECT	118.625 31.148 118.657 31.212 ;
			RECT	118.793 31.148 118.825 31.212 ;
			RECT	118.961 31.148 118.993 31.212 ;
			RECT	119.129 31.148 119.161 31.212 ;
			RECT	119.297 31.148 119.329 31.212 ;
			RECT	119.465 31.148 119.497 31.212 ;
			RECT	119.633 31.148 119.665 31.212 ;
			RECT	119.801 31.148 119.833 31.212 ;
			RECT	119.969 31.148 120.001 31.212 ;
			RECT	120.137 31.148 120.169 31.212 ;
			RECT	120.305 31.148 120.337 31.212 ;
			RECT	120.473 31.148 120.505 31.212 ;
			RECT	120.641 31.148 120.673 31.212 ;
			RECT	120.809 31.148 120.841 31.212 ;
			RECT	120.977 31.148 121.009 31.212 ;
			RECT	121.145 31.148 121.177 31.212 ;
			RECT	121.313 31.148 121.345 31.212 ;
			RECT	121.481 31.148 121.513 31.212 ;
			RECT	121.649 31.148 121.681 31.212 ;
			RECT	121.817 31.148 121.849 31.212 ;
			RECT	121.985 31.148 122.017 31.212 ;
			RECT	122.153 31.148 122.185 31.212 ;
			RECT	122.321 31.148 122.353 31.212 ;
			RECT	122.489 31.148 122.521 31.212 ;
			RECT	122.657 31.148 122.689 31.212 ;
			RECT	122.825 31.148 122.857 31.212 ;
			RECT	122.993 31.148 123.025 31.212 ;
			RECT	123.161 31.148 123.193 31.212 ;
			RECT	123.329 31.148 123.361 31.212 ;
			RECT	123.497 31.148 123.529 31.212 ;
			RECT	123.665 31.148 123.697 31.212 ;
			RECT	123.833 31.148 123.865 31.212 ;
			RECT	124.001 31.148 124.033 31.212 ;
			RECT	124.169 31.148 124.201 31.212 ;
			RECT	124.337 31.148 124.369 31.212 ;
			RECT	124.505 31.148 124.537 31.212 ;
			RECT	124.673 31.148 124.705 31.212 ;
			RECT	124.841 31.148 124.873 31.212 ;
			RECT	125.009 31.148 125.041 31.212 ;
			RECT	125.177 31.148 125.209 31.212 ;
			RECT	125.345 31.148 125.377 31.212 ;
			RECT	125.513 31.148 125.545 31.212 ;
			RECT	125.681 31.148 125.713 31.212 ;
			RECT	125.849 31.148 125.881 31.212 ;
			RECT	126.017 31.148 126.049 31.212 ;
			RECT	126.185 31.148 126.217 31.212 ;
			RECT	126.353 31.148 126.385 31.212 ;
			RECT	126.521 31.148 126.553 31.212 ;
			RECT	126.689 31.148 126.721 31.212 ;
			RECT	126.857 31.148 126.889 31.212 ;
			RECT	127.025 31.148 127.057 31.212 ;
			RECT	127.193 31.148 127.225 31.212 ;
			RECT	127.361 31.148 127.393 31.212 ;
			RECT	127.529 31.148 127.561 31.212 ;
			RECT	127.697 31.148 127.729 31.212 ;
			RECT	127.865 31.148 127.897 31.212 ;
			RECT	128.033 31.148 128.065 31.212 ;
			RECT	128.201 31.148 128.233 31.212 ;
			RECT	128.369 31.148 128.401 31.212 ;
			RECT	128.537 31.148 128.569 31.212 ;
			RECT	128.705 31.148 128.737 31.212 ;
			RECT	128.873 31.148 128.905 31.212 ;
			RECT	129.041 31.148 129.073 31.212 ;
			RECT	129.209 31.148 129.241 31.212 ;
			RECT	129.377 31.148 129.409 31.212 ;
			RECT	129.545 31.148 129.577 31.212 ;
			RECT	129.713 31.148 129.745 31.212 ;
			RECT	129.881 31.148 129.913 31.212 ;
			RECT	130.049 31.148 130.081 31.212 ;
			RECT	130.217 31.148 130.249 31.212 ;
			RECT	130.385 31.148 130.417 31.212 ;
			RECT	130.553 31.148 130.585 31.212 ;
			RECT	130.721 31.148 130.753 31.212 ;
			RECT	130.889 31.148 130.921 31.212 ;
			RECT	131.057 31.148 131.089 31.212 ;
			RECT	131.225 31.148 131.257 31.212 ;
			RECT	131.393 31.148 131.425 31.212 ;
			RECT	131.561 31.148 131.593 31.212 ;
			RECT	131.729 31.148 131.761 31.212 ;
			RECT	131.897 31.148 131.929 31.212 ;
			RECT	132.065 31.148 132.097 31.212 ;
			RECT	132.233 31.148 132.265 31.212 ;
			RECT	132.401 31.148 132.433 31.212 ;
			RECT	132.569 31.148 132.601 31.212 ;
			RECT	132.737 31.148 132.769 31.212 ;
			RECT	132.905 31.148 132.937 31.212 ;
			RECT	133.073 31.148 133.105 31.212 ;
			RECT	133.241 31.148 133.273 31.212 ;
			RECT	133.409 31.148 133.441 31.212 ;
			RECT	133.577 31.148 133.609 31.212 ;
			RECT	133.745 31.148 133.777 31.212 ;
			RECT	133.913 31.148 133.945 31.212 ;
			RECT	134.081 31.148 134.113 31.212 ;
			RECT	134.249 31.148 134.281 31.212 ;
			RECT	134.417 31.148 134.449 31.212 ;
			RECT	134.585 31.148 134.617 31.212 ;
			RECT	134.753 31.148 134.785 31.212 ;
			RECT	134.921 31.148 134.953 31.212 ;
			RECT	135.089 31.148 135.121 31.212 ;
			RECT	135.257 31.148 135.289 31.212 ;
			RECT	135.425 31.148 135.457 31.212 ;
			RECT	135.593 31.148 135.625 31.212 ;
			RECT	135.761 31.148 135.793 31.212 ;
			RECT	135.929 31.148 135.961 31.212 ;
			RECT	136.097 31.148 136.129 31.212 ;
			RECT	136.265 31.148 136.297 31.212 ;
			RECT	136.433 31.148 136.465 31.212 ;
			RECT	136.601 31.148 136.633 31.212 ;
			RECT	136.769 31.148 136.801 31.212 ;
			RECT	136.937 31.148 136.969 31.212 ;
			RECT	137.105 31.148 137.137 31.212 ;
			RECT	137.273 31.148 137.305 31.212 ;
			RECT	137.441 31.148 137.473 31.212 ;
			RECT	137.609 31.148 137.641 31.212 ;
			RECT	137.777 31.148 137.809 31.212 ;
			RECT	137.945 31.148 137.977 31.212 ;
			RECT	138.113 31.148 138.145 31.212 ;
			RECT	138.281 31.148 138.313 31.212 ;
			RECT	138.449 31.148 138.481 31.212 ;
			RECT	138.617 31.148 138.649 31.212 ;
			RECT	138.785 31.148 138.817 31.212 ;
			RECT	138.953 31.148 138.985 31.212 ;
			RECT	139.121 31.148 139.153 31.212 ;
			RECT	139.289 31.148 139.321 31.212 ;
			RECT	139.457 31.148 139.489 31.212 ;
			RECT	139.625 31.148 139.657 31.212 ;
			RECT	139.793 31.148 139.825 31.212 ;
			RECT	139.961 31.148 139.993 31.212 ;
			RECT	140.129 31.148 140.161 31.212 ;
			RECT	140.297 31.148 140.329 31.212 ;
			RECT	140.465 31.148 140.497 31.212 ;
			RECT	140.633 31.148 140.665 31.212 ;
			RECT	140.801 31.148 140.833 31.212 ;
			RECT	140.969 31.148 141.001 31.212 ;
			RECT	141.137 31.148 141.169 31.212 ;
			RECT	141.305 31.148 141.337 31.212 ;
			RECT	141.473 31.148 141.505 31.212 ;
			RECT	141.641 31.148 141.673 31.212 ;
			RECT	141.809 31.148 141.841 31.212 ;
			RECT	141.977 31.148 142.009 31.212 ;
			RECT	142.145 31.148 142.177 31.212 ;
			RECT	142.313 31.148 142.345 31.212 ;
			RECT	142.481 31.148 142.513 31.212 ;
			RECT	142.649 31.148 142.681 31.212 ;
			RECT	142.817 31.148 142.849 31.212 ;
			RECT	142.985 31.148 143.017 31.212 ;
			RECT	143.153 31.148 143.185 31.212 ;
			RECT	143.321 31.148 143.353 31.212 ;
			RECT	143.489 31.148 143.521 31.212 ;
			RECT	143.657 31.148 143.689 31.212 ;
			RECT	143.825 31.148 143.857 31.212 ;
			RECT	143.993 31.148 144.025 31.212 ;
			RECT	144.161 31.148 144.193 31.212 ;
			RECT	144.329 31.148 144.361 31.212 ;
			RECT	144.497 31.148 144.529 31.212 ;
			RECT	144.665 31.148 144.697 31.212 ;
			RECT	144.833 31.148 144.865 31.212 ;
			RECT	145.001 31.148 145.033 31.212 ;
			RECT	145.169 31.148 145.201 31.212 ;
			RECT	145.337 31.148 145.369 31.212 ;
			RECT	145.505 31.148 145.537 31.212 ;
			RECT	145.673 31.148 145.705 31.212 ;
			RECT	145.841 31.148 145.873 31.212 ;
			RECT	146.009 31.148 146.041 31.212 ;
			RECT	146.177 31.148 146.209 31.212 ;
			RECT	146.345 31.148 146.377 31.212 ;
			RECT	146.513 31.148 146.545 31.212 ;
			RECT	146.681 31.148 146.713 31.212 ;
			RECT	146.849 31.148 146.881 31.212 ;
			RECT	147.017 31.148 147.049 31.212 ;
			RECT	147.185 31.148 147.217 31.212 ;
			RECT	147.316 31.164 147.348 31.196 ;
			RECT	147.437 31.164 147.469 31.196 ;
			RECT	147.567 31.148 147.599 31.212 ;
			RECT	149.879 31.148 149.911 31.212 ;
			RECT	151.13 31.148 151.194 31.212 ;
			RECT	151.81 31.148 151.842 31.212 ;
			RECT	152.249 31.148 152.281 31.212 ;
			RECT	153.56 31.148 153.624 31.212 ;
			RECT	156.601 31.148 156.633 31.212 ;
			RECT	156.731 31.164 156.763 31.196 ;
			RECT	156.852 31.164 156.884 31.196 ;
			RECT	156.983 31.148 157.015 31.212 ;
			RECT	157.151 31.148 157.183 31.212 ;
			RECT	157.319 31.148 157.351 31.212 ;
			RECT	157.487 31.148 157.519 31.212 ;
			RECT	157.655 31.148 157.687 31.212 ;
			RECT	157.823 31.148 157.855 31.212 ;
			RECT	157.991 31.148 158.023 31.212 ;
			RECT	158.159 31.148 158.191 31.212 ;
			RECT	158.327 31.148 158.359 31.212 ;
			RECT	158.495 31.148 158.527 31.212 ;
			RECT	158.663 31.148 158.695 31.212 ;
			RECT	158.831 31.148 158.863 31.212 ;
			RECT	158.999 31.148 159.031 31.212 ;
			RECT	159.167 31.148 159.199 31.212 ;
			RECT	159.335 31.148 159.367 31.212 ;
			RECT	159.503 31.148 159.535 31.212 ;
			RECT	159.671 31.148 159.703 31.212 ;
			RECT	159.839 31.148 159.871 31.212 ;
			RECT	160.007 31.148 160.039 31.212 ;
			RECT	160.175 31.148 160.207 31.212 ;
			RECT	160.343 31.148 160.375 31.212 ;
			RECT	160.511 31.148 160.543 31.212 ;
			RECT	160.679 31.148 160.711 31.212 ;
			RECT	160.847 31.148 160.879 31.212 ;
			RECT	161.015 31.148 161.047 31.212 ;
			RECT	161.183 31.148 161.215 31.212 ;
			RECT	161.351 31.148 161.383 31.212 ;
			RECT	161.519 31.148 161.551 31.212 ;
			RECT	161.687 31.148 161.719 31.212 ;
			RECT	161.855 31.148 161.887 31.212 ;
			RECT	162.023 31.148 162.055 31.212 ;
			RECT	162.191 31.148 162.223 31.212 ;
			RECT	162.359 31.148 162.391 31.212 ;
			RECT	162.527 31.148 162.559 31.212 ;
			RECT	162.695 31.148 162.727 31.212 ;
			RECT	162.863 31.148 162.895 31.212 ;
			RECT	163.031 31.148 163.063 31.212 ;
			RECT	163.199 31.148 163.231 31.212 ;
			RECT	163.367 31.148 163.399 31.212 ;
			RECT	163.535 31.148 163.567 31.212 ;
			RECT	163.703 31.148 163.735 31.212 ;
			RECT	163.871 31.148 163.903 31.212 ;
			RECT	164.039 31.148 164.071 31.212 ;
			RECT	164.207 31.148 164.239 31.212 ;
			RECT	164.375 31.148 164.407 31.212 ;
			RECT	164.543 31.148 164.575 31.212 ;
			RECT	164.711 31.148 164.743 31.212 ;
			RECT	164.879 31.148 164.911 31.212 ;
			RECT	165.047 31.148 165.079 31.212 ;
			RECT	165.215 31.148 165.247 31.212 ;
			RECT	165.383 31.148 165.415 31.212 ;
			RECT	165.551 31.148 165.583 31.212 ;
			RECT	165.719 31.148 165.751 31.212 ;
			RECT	165.887 31.148 165.919 31.212 ;
			RECT	166.055 31.148 166.087 31.212 ;
			RECT	166.223 31.148 166.255 31.212 ;
			RECT	166.391 31.148 166.423 31.212 ;
			RECT	166.559 31.148 166.591 31.212 ;
			RECT	166.727 31.148 166.759 31.212 ;
			RECT	166.895 31.148 166.927 31.212 ;
			RECT	167.063 31.148 167.095 31.212 ;
			RECT	167.231 31.148 167.263 31.212 ;
			RECT	167.399 31.148 167.431 31.212 ;
			RECT	167.567 31.148 167.599 31.212 ;
			RECT	167.735 31.148 167.767 31.212 ;
			RECT	167.903 31.148 167.935 31.212 ;
			RECT	168.071 31.148 168.103 31.212 ;
			RECT	168.239 31.148 168.271 31.212 ;
			RECT	168.407 31.148 168.439 31.212 ;
			RECT	168.575 31.148 168.607 31.212 ;
			RECT	168.743 31.148 168.775 31.212 ;
			RECT	168.911 31.148 168.943 31.212 ;
			RECT	169.079 31.148 169.111 31.212 ;
			RECT	169.247 31.148 169.279 31.212 ;
			RECT	169.415 31.148 169.447 31.212 ;
			RECT	169.583 31.148 169.615 31.212 ;
			RECT	169.751 31.148 169.783 31.212 ;
			RECT	169.919 31.148 169.951 31.212 ;
			RECT	170.087 31.148 170.119 31.212 ;
			RECT	170.255 31.148 170.287 31.212 ;
			RECT	170.423 31.148 170.455 31.212 ;
			RECT	170.591 31.148 170.623 31.212 ;
			RECT	170.759 31.148 170.791 31.212 ;
			RECT	170.927 31.148 170.959 31.212 ;
			RECT	171.095 31.148 171.127 31.212 ;
			RECT	171.263 31.148 171.295 31.212 ;
			RECT	171.431 31.148 171.463 31.212 ;
			RECT	171.599 31.148 171.631 31.212 ;
			RECT	171.767 31.148 171.799 31.212 ;
			RECT	171.935 31.148 171.967 31.212 ;
			RECT	172.103 31.148 172.135 31.212 ;
			RECT	172.271 31.148 172.303 31.212 ;
			RECT	172.439 31.148 172.471 31.212 ;
			RECT	172.607 31.148 172.639 31.212 ;
			RECT	172.775 31.148 172.807 31.212 ;
			RECT	172.943 31.148 172.975 31.212 ;
			RECT	173.111 31.148 173.143 31.212 ;
			RECT	173.279 31.148 173.311 31.212 ;
			RECT	173.447 31.148 173.479 31.212 ;
			RECT	173.615 31.148 173.647 31.212 ;
			RECT	173.783 31.148 173.815 31.212 ;
			RECT	173.951 31.148 173.983 31.212 ;
			RECT	174.119 31.148 174.151 31.212 ;
			RECT	174.287 31.148 174.319 31.212 ;
			RECT	174.455 31.148 174.487 31.212 ;
			RECT	174.623 31.148 174.655 31.212 ;
			RECT	174.791 31.148 174.823 31.212 ;
			RECT	174.959 31.148 174.991 31.212 ;
			RECT	175.127 31.148 175.159 31.212 ;
			RECT	175.295 31.148 175.327 31.212 ;
			RECT	175.463 31.148 175.495 31.212 ;
			RECT	175.631 31.148 175.663 31.212 ;
			RECT	175.799 31.148 175.831 31.212 ;
			RECT	175.967 31.148 175.999 31.212 ;
			RECT	176.135 31.148 176.167 31.212 ;
			RECT	176.303 31.148 176.335 31.212 ;
			RECT	176.471 31.148 176.503 31.212 ;
			RECT	176.639 31.148 176.671 31.212 ;
			RECT	176.807 31.148 176.839 31.212 ;
			RECT	176.975 31.148 177.007 31.212 ;
			RECT	177.143 31.148 177.175 31.212 ;
			RECT	177.311 31.148 177.343 31.212 ;
			RECT	177.479 31.148 177.511 31.212 ;
			RECT	177.647 31.148 177.679 31.212 ;
			RECT	177.815 31.148 177.847 31.212 ;
			RECT	177.983 31.148 178.015 31.212 ;
			RECT	178.151 31.148 178.183 31.212 ;
			RECT	178.319 31.148 178.351 31.212 ;
			RECT	178.487 31.148 178.519 31.212 ;
			RECT	178.655 31.148 178.687 31.212 ;
			RECT	178.823 31.148 178.855 31.212 ;
			RECT	178.991 31.148 179.023 31.212 ;
			RECT	179.159 31.148 179.191 31.212 ;
			RECT	179.327 31.148 179.359 31.212 ;
			RECT	179.495 31.148 179.527 31.212 ;
			RECT	179.663 31.148 179.695 31.212 ;
			RECT	179.831 31.148 179.863 31.212 ;
			RECT	179.999 31.148 180.031 31.212 ;
			RECT	180.167 31.148 180.199 31.212 ;
			RECT	180.335 31.148 180.367 31.212 ;
			RECT	180.503 31.148 180.535 31.212 ;
			RECT	180.671 31.148 180.703 31.212 ;
			RECT	180.839 31.148 180.871 31.212 ;
			RECT	181.007 31.148 181.039 31.212 ;
			RECT	181.175 31.148 181.207 31.212 ;
			RECT	181.343 31.148 181.375 31.212 ;
			RECT	181.511 31.148 181.543 31.212 ;
			RECT	181.679 31.148 181.711 31.212 ;
			RECT	181.847 31.148 181.879 31.212 ;
			RECT	182.015 31.148 182.047 31.212 ;
			RECT	182.183 31.148 182.215 31.212 ;
			RECT	182.351 31.148 182.383 31.212 ;
			RECT	182.519 31.148 182.551 31.212 ;
			RECT	182.687 31.148 182.719 31.212 ;
			RECT	182.855 31.148 182.887 31.212 ;
			RECT	183.023 31.148 183.055 31.212 ;
			RECT	183.191 31.148 183.223 31.212 ;
			RECT	183.359 31.148 183.391 31.212 ;
			RECT	183.527 31.148 183.559 31.212 ;
			RECT	183.695 31.148 183.727 31.212 ;
			RECT	183.863 31.148 183.895 31.212 ;
			RECT	184.031 31.148 184.063 31.212 ;
			RECT	184.199 31.148 184.231 31.212 ;
			RECT	184.367 31.148 184.399 31.212 ;
			RECT	184.535 31.148 184.567 31.212 ;
			RECT	184.703 31.148 184.735 31.212 ;
			RECT	184.871 31.148 184.903 31.212 ;
			RECT	185.039 31.148 185.071 31.212 ;
			RECT	185.207 31.148 185.239 31.212 ;
			RECT	185.375 31.148 185.407 31.212 ;
			RECT	185.543 31.148 185.575 31.212 ;
			RECT	185.711 31.148 185.743 31.212 ;
			RECT	185.879 31.148 185.911 31.212 ;
			RECT	186.047 31.148 186.079 31.212 ;
			RECT	186.215 31.148 186.247 31.212 ;
			RECT	186.383 31.148 186.415 31.212 ;
			RECT	186.551 31.148 186.583 31.212 ;
			RECT	186.719 31.148 186.751 31.212 ;
			RECT	186.887 31.148 186.919 31.212 ;
			RECT	187.055 31.148 187.087 31.212 ;
			RECT	187.223 31.148 187.255 31.212 ;
			RECT	187.391 31.148 187.423 31.212 ;
			RECT	187.559 31.148 187.591 31.212 ;
			RECT	187.727 31.148 187.759 31.212 ;
			RECT	187.895 31.148 187.927 31.212 ;
			RECT	188.063 31.148 188.095 31.212 ;
			RECT	188.231 31.148 188.263 31.212 ;
			RECT	188.399 31.148 188.431 31.212 ;
			RECT	188.567 31.148 188.599 31.212 ;
			RECT	188.735 31.148 188.767 31.212 ;
			RECT	188.903 31.148 188.935 31.212 ;
			RECT	189.071 31.148 189.103 31.212 ;
			RECT	189.239 31.148 189.271 31.212 ;
			RECT	189.407 31.148 189.439 31.212 ;
			RECT	189.575 31.148 189.607 31.212 ;
			RECT	189.743 31.148 189.775 31.212 ;
			RECT	189.911 31.148 189.943 31.212 ;
			RECT	190.079 31.148 190.111 31.212 ;
			RECT	190.247 31.148 190.279 31.212 ;
			RECT	190.415 31.148 190.447 31.212 ;
			RECT	190.583 31.148 190.615 31.212 ;
			RECT	190.751 31.148 190.783 31.212 ;
			RECT	190.919 31.148 190.951 31.212 ;
			RECT	191.087 31.148 191.119 31.212 ;
			RECT	191.255 31.148 191.287 31.212 ;
			RECT	191.423 31.148 191.455 31.212 ;
			RECT	191.591 31.148 191.623 31.212 ;
			RECT	191.759 31.148 191.791 31.212 ;
			RECT	191.927 31.148 191.959 31.212 ;
			RECT	192.095 31.148 192.127 31.212 ;
			RECT	192.263 31.148 192.295 31.212 ;
			RECT	192.431 31.148 192.463 31.212 ;
			RECT	192.599 31.148 192.631 31.212 ;
			RECT	192.767 31.148 192.799 31.212 ;
			RECT	192.935 31.148 192.967 31.212 ;
			RECT	193.103 31.148 193.135 31.212 ;
			RECT	193.271 31.148 193.303 31.212 ;
			RECT	193.439 31.148 193.471 31.212 ;
			RECT	193.607 31.148 193.639 31.212 ;
			RECT	193.775 31.148 193.807 31.212 ;
			RECT	193.943 31.148 193.975 31.212 ;
			RECT	194.111 31.148 194.143 31.212 ;
			RECT	194.279 31.148 194.311 31.212 ;
			RECT	194.447 31.148 194.479 31.212 ;
			RECT	194.615 31.148 194.647 31.212 ;
			RECT	194.783 31.148 194.815 31.212 ;
			RECT	194.951 31.148 194.983 31.212 ;
			RECT	195.119 31.148 195.151 31.212 ;
			RECT	195.287 31.148 195.319 31.212 ;
			RECT	195.455 31.148 195.487 31.212 ;
			RECT	195.623 31.148 195.655 31.212 ;
			RECT	195.791 31.148 195.823 31.212 ;
			RECT	195.959 31.148 195.991 31.212 ;
			RECT	196.127 31.148 196.159 31.212 ;
			RECT	196.295 31.148 196.327 31.212 ;
			RECT	196.463 31.148 196.495 31.212 ;
			RECT	196.631 31.148 196.663 31.212 ;
			RECT	196.799 31.148 196.831 31.212 ;
			RECT	196.967 31.148 196.999 31.212 ;
			RECT	197.135 31.148 197.167 31.212 ;
			RECT	197.303 31.148 197.335 31.212 ;
			RECT	197.471 31.148 197.503 31.212 ;
			RECT	197.639 31.148 197.671 31.212 ;
			RECT	197.807 31.148 197.839 31.212 ;
			RECT	197.975 31.148 198.007 31.212 ;
			RECT	198.143 31.148 198.175 31.212 ;
			RECT	198.311 31.148 198.343 31.212 ;
			RECT	198.479 31.148 198.511 31.212 ;
			RECT	198.647 31.148 198.679 31.212 ;
			RECT	198.815 31.148 198.847 31.212 ;
			RECT	198.983 31.148 199.015 31.212 ;
			RECT	199.151 31.148 199.183 31.212 ;
			RECT	199.319 31.148 199.351 31.212 ;
			RECT	199.487 31.148 199.519 31.212 ;
			RECT	199.655 31.148 199.687 31.212 ;
			RECT	199.823 31.148 199.855 31.212 ;
			RECT	199.991 31.148 200.023 31.212 ;
			RECT	200.121 31.164 200.153 31.196 ;
			RECT	200.243 31.169 200.275 31.201 ;
			RECT	200.373 31.148 200.405 31.212 ;
			RECT	200.9 31.148 200.932 31.212 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 29.2 201.665 29.32 ;
			LAYER	J3 ;
			RECT	0.755 29.228 0.787 29.292 ;
			RECT	1.645 29.228 1.709 29.292 ;
			RECT	2.323 29.228 2.387 29.292 ;
			RECT	3.438 29.228 3.47 29.292 ;
			RECT	3.585 29.228 3.617 29.292 ;
			RECT	4.195 29.228 4.227 29.292 ;
			RECT	4.72 29.228 4.752 29.292 ;
			RECT	4.944 29.228 5.008 29.292 ;
			RECT	5.267 29.228 5.299 29.292 ;
			RECT	5.797 29.228 5.829 29.292 ;
			RECT	5.927 29.249 5.959 29.281 ;
			RECT	6.049 29.244 6.081 29.276 ;
			RECT	6.179 29.228 6.211 29.292 ;
			RECT	6.347 29.228 6.379 29.292 ;
			RECT	6.515 29.228 6.547 29.292 ;
			RECT	6.683 29.228 6.715 29.292 ;
			RECT	6.851 29.228 6.883 29.292 ;
			RECT	7.019 29.228 7.051 29.292 ;
			RECT	7.187 29.228 7.219 29.292 ;
			RECT	7.355 29.228 7.387 29.292 ;
			RECT	7.523 29.228 7.555 29.292 ;
			RECT	7.691 29.228 7.723 29.292 ;
			RECT	7.859 29.228 7.891 29.292 ;
			RECT	8.027 29.228 8.059 29.292 ;
			RECT	8.195 29.228 8.227 29.292 ;
			RECT	8.363 29.228 8.395 29.292 ;
			RECT	8.531 29.228 8.563 29.292 ;
			RECT	8.699 29.228 8.731 29.292 ;
			RECT	8.867 29.228 8.899 29.292 ;
			RECT	9.035 29.228 9.067 29.292 ;
			RECT	9.203 29.228 9.235 29.292 ;
			RECT	9.371 29.228 9.403 29.292 ;
			RECT	9.539 29.228 9.571 29.292 ;
			RECT	9.707 29.228 9.739 29.292 ;
			RECT	9.875 29.228 9.907 29.292 ;
			RECT	10.043 29.228 10.075 29.292 ;
			RECT	10.211 29.228 10.243 29.292 ;
			RECT	10.379 29.228 10.411 29.292 ;
			RECT	10.547 29.228 10.579 29.292 ;
			RECT	10.715 29.228 10.747 29.292 ;
			RECT	10.883 29.228 10.915 29.292 ;
			RECT	11.051 29.228 11.083 29.292 ;
			RECT	11.219 29.228 11.251 29.292 ;
			RECT	11.387 29.228 11.419 29.292 ;
			RECT	11.555 29.228 11.587 29.292 ;
			RECT	11.723 29.228 11.755 29.292 ;
			RECT	11.891 29.228 11.923 29.292 ;
			RECT	12.059 29.228 12.091 29.292 ;
			RECT	12.227 29.228 12.259 29.292 ;
			RECT	12.395 29.228 12.427 29.292 ;
			RECT	12.563 29.228 12.595 29.292 ;
			RECT	12.731 29.228 12.763 29.292 ;
			RECT	12.899 29.228 12.931 29.292 ;
			RECT	13.067 29.228 13.099 29.292 ;
			RECT	13.235 29.228 13.267 29.292 ;
			RECT	13.403 29.228 13.435 29.292 ;
			RECT	13.571 29.228 13.603 29.292 ;
			RECT	13.739 29.228 13.771 29.292 ;
			RECT	13.907 29.228 13.939 29.292 ;
			RECT	14.075 29.228 14.107 29.292 ;
			RECT	14.243 29.228 14.275 29.292 ;
			RECT	14.411 29.228 14.443 29.292 ;
			RECT	14.579 29.228 14.611 29.292 ;
			RECT	14.747 29.228 14.779 29.292 ;
			RECT	14.915 29.228 14.947 29.292 ;
			RECT	15.083 29.228 15.115 29.292 ;
			RECT	15.251 29.228 15.283 29.292 ;
			RECT	15.419 29.228 15.451 29.292 ;
			RECT	15.587 29.228 15.619 29.292 ;
			RECT	15.755 29.228 15.787 29.292 ;
			RECT	15.923 29.228 15.955 29.292 ;
			RECT	16.091 29.228 16.123 29.292 ;
			RECT	16.259 29.228 16.291 29.292 ;
			RECT	16.427 29.228 16.459 29.292 ;
			RECT	16.595 29.228 16.627 29.292 ;
			RECT	16.763 29.228 16.795 29.292 ;
			RECT	16.931 29.228 16.963 29.292 ;
			RECT	17.099 29.228 17.131 29.292 ;
			RECT	17.267 29.228 17.299 29.292 ;
			RECT	17.435 29.228 17.467 29.292 ;
			RECT	17.603 29.228 17.635 29.292 ;
			RECT	17.771 29.228 17.803 29.292 ;
			RECT	17.939 29.228 17.971 29.292 ;
			RECT	18.107 29.228 18.139 29.292 ;
			RECT	18.275 29.228 18.307 29.292 ;
			RECT	18.443 29.228 18.475 29.292 ;
			RECT	18.611 29.228 18.643 29.292 ;
			RECT	18.779 29.228 18.811 29.292 ;
			RECT	18.947 29.228 18.979 29.292 ;
			RECT	19.115 29.228 19.147 29.292 ;
			RECT	19.283 29.228 19.315 29.292 ;
			RECT	19.451 29.228 19.483 29.292 ;
			RECT	19.619 29.228 19.651 29.292 ;
			RECT	19.787 29.228 19.819 29.292 ;
			RECT	19.955 29.228 19.987 29.292 ;
			RECT	20.123 29.228 20.155 29.292 ;
			RECT	20.291 29.228 20.323 29.292 ;
			RECT	20.459 29.228 20.491 29.292 ;
			RECT	20.627 29.228 20.659 29.292 ;
			RECT	20.795 29.228 20.827 29.292 ;
			RECT	20.963 29.228 20.995 29.292 ;
			RECT	21.131 29.228 21.163 29.292 ;
			RECT	21.299 29.228 21.331 29.292 ;
			RECT	21.467 29.228 21.499 29.292 ;
			RECT	21.635 29.228 21.667 29.292 ;
			RECT	21.803 29.228 21.835 29.292 ;
			RECT	21.971 29.228 22.003 29.292 ;
			RECT	22.139 29.228 22.171 29.292 ;
			RECT	22.307 29.228 22.339 29.292 ;
			RECT	22.475 29.228 22.507 29.292 ;
			RECT	22.643 29.228 22.675 29.292 ;
			RECT	22.811 29.228 22.843 29.292 ;
			RECT	22.979 29.228 23.011 29.292 ;
			RECT	23.147 29.228 23.179 29.292 ;
			RECT	23.315 29.228 23.347 29.292 ;
			RECT	23.483 29.228 23.515 29.292 ;
			RECT	23.651 29.228 23.683 29.292 ;
			RECT	23.819 29.228 23.851 29.292 ;
			RECT	23.987 29.228 24.019 29.292 ;
			RECT	24.155 29.228 24.187 29.292 ;
			RECT	24.323 29.228 24.355 29.292 ;
			RECT	24.491 29.228 24.523 29.292 ;
			RECT	24.659 29.228 24.691 29.292 ;
			RECT	24.827 29.228 24.859 29.292 ;
			RECT	24.995 29.228 25.027 29.292 ;
			RECT	25.163 29.228 25.195 29.292 ;
			RECT	25.331 29.228 25.363 29.292 ;
			RECT	25.499 29.228 25.531 29.292 ;
			RECT	25.667 29.228 25.699 29.292 ;
			RECT	25.835 29.228 25.867 29.292 ;
			RECT	26.003 29.228 26.035 29.292 ;
			RECT	26.171 29.228 26.203 29.292 ;
			RECT	26.339 29.228 26.371 29.292 ;
			RECT	26.507 29.228 26.539 29.292 ;
			RECT	26.675 29.228 26.707 29.292 ;
			RECT	26.843 29.228 26.875 29.292 ;
			RECT	27.011 29.228 27.043 29.292 ;
			RECT	27.179 29.228 27.211 29.292 ;
			RECT	27.347 29.228 27.379 29.292 ;
			RECT	27.515 29.228 27.547 29.292 ;
			RECT	27.683 29.228 27.715 29.292 ;
			RECT	27.851 29.228 27.883 29.292 ;
			RECT	28.019 29.228 28.051 29.292 ;
			RECT	28.187 29.228 28.219 29.292 ;
			RECT	28.355 29.228 28.387 29.292 ;
			RECT	28.523 29.228 28.555 29.292 ;
			RECT	28.691 29.228 28.723 29.292 ;
			RECT	28.859 29.228 28.891 29.292 ;
			RECT	29.027 29.228 29.059 29.292 ;
			RECT	29.195 29.228 29.227 29.292 ;
			RECT	29.363 29.228 29.395 29.292 ;
			RECT	29.531 29.228 29.563 29.292 ;
			RECT	29.699 29.228 29.731 29.292 ;
			RECT	29.867 29.228 29.899 29.292 ;
			RECT	30.035 29.228 30.067 29.292 ;
			RECT	30.203 29.228 30.235 29.292 ;
			RECT	30.371 29.228 30.403 29.292 ;
			RECT	30.539 29.228 30.571 29.292 ;
			RECT	30.707 29.228 30.739 29.292 ;
			RECT	30.875 29.228 30.907 29.292 ;
			RECT	31.043 29.228 31.075 29.292 ;
			RECT	31.211 29.228 31.243 29.292 ;
			RECT	31.379 29.228 31.411 29.292 ;
			RECT	31.547 29.228 31.579 29.292 ;
			RECT	31.715 29.228 31.747 29.292 ;
			RECT	31.883 29.228 31.915 29.292 ;
			RECT	32.051 29.228 32.083 29.292 ;
			RECT	32.219 29.228 32.251 29.292 ;
			RECT	32.387 29.228 32.419 29.292 ;
			RECT	32.555 29.228 32.587 29.292 ;
			RECT	32.723 29.228 32.755 29.292 ;
			RECT	32.891 29.228 32.923 29.292 ;
			RECT	33.059 29.228 33.091 29.292 ;
			RECT	33.227 29.228 33.259 29.292 ;
			RECT	33.395 29.228 33.427 29.292 ;
			RECT	33.563 29.228 33.595 29.292 ;
			RECT	33.731 29.228 33.763 29.292 ;
			RECT	33.899 29.228 33.931 29.292 ;
			RECT	34.067 29.228 34.099 29.292 ;
			RECT	34.235 29.228 34.267 29.292 ;
			RECT	34.403 29.228 34.435 29.292 ;
			RECT	34.571 29.228 34.603 29.292 ;
			RECT	34.739 29.228 34.771 29.292 ;
			RECT	34.907 29.228 34.939 29.292 ;
			RECT	35.075 29.228 35.107 29.292 ;
			RECT	35.243 29.228 35.275 29.292 ;
			RECT	35.411 29.228 35.443 29.292 ;
			RECT	35.579 29.228 35.611 29.292 ;
			RECT	35.747 29.228 35.779 29.292 ;
			RECT	35.915 29.228 35.947 29.292 ;
			RECT	36.083 29.228 36.115 29.292 ;
			RECT	36.251 29.228 36.283 29.292 ;
			RECT	36.419 29.228 36.451 29.292 ;
			RECT	36.587 29.228 36.619 29.292 ;
			RECT	36.755 29.228 36.787 29.292 ;
			RECT	36.923 29.228 36.955 29.292 ;
			RECT	37.091 29.228 37.123 29.292 ;
			RECT	37.259 29.228 37.291 29.292 ;
			RECT	37.427 29.228 37.459 29.292 ;
			RECT	37.595 29.228 37.627 29.292 ;
			RECT	37.763 29.228 37.795 29.292 ;
			RECT	37.931 29.228 37.963 29.292 ;
			RECT	38.099 29.228 38.131 29.292 ;
			RECT	38.267 29.228 38.299 29.292 ;
			RECT	38.435 29.228 38.467 29.292 ;
			RECT	38.603 29.228 38.635 29.292 ;
			RECT	38.771 29.228 38.803 29.292 ;
			RECT	38.939 29.228 38.971 29.292 ;
			RECT	39.107 29.228 39.139 29.292 ;
			RECT	39.275 29.228 39.307 29.292 ;
			RECT	39.443 29.228 39.475 29.292 ;
			RECT	39.611 29.228 39.643 29.292 ;
			RECT	39.779 29.228 39.811 29.292 ;
			RECT	39.947 29.228 39.979 29.292 ;
			RECT	40.115 29.228 40.147 29.292 ;
			RECT	40.283 29.228 40.315 29.292 ;
			RECT	40.451 29.228 40.483 29.292 ;
			RECT	40.619 29.228 40.651 29.292 ;
			RECT	40.787 29.228 40.819 29.292 ;
			RECT	40.955 29.228 40.987 29.292 ;
			RECT	41.123 29.228 41.155 29.292 ;
			RECT	41.291 29.228 41.323 29.292 ;
			RECT	41.459 29.228 41.491 29.292 ;
			RECT	41.627 29.228 41.659 29.292 ;
			RECT	41.795 29.228 41.827 29.292 ;
			RECT	41.963 29.228 41.995 29.292 ;
			RECT	42.131 29.228 42.163 29.292 ;
			RECT	42.299 29.228 42.331 29.292 ;
			RECT	42.467 29.228 42.499 29.292 ;
			RECT	42.635 29.228 42.667 29.292 ;
			RECT	42.803 29.228 42.835 29.292 ;
			RECT	42.971 29.228 43.003 29.292 ;
			RECT	43.139 29.228 43.171 29.292 ;
			RECT	43.307 29.228 43.339 29.292 ;
			RECT	43.475 29.228 43.507 29.292 ;
			RECT	43.643 29.228 43.675 29.292 ;
			RECT	43.811 29.228 43.843 29.292 ;
			RECT	43.979 29.228 44.011 29.292 ;
			RECT	44.147 29.228 44.179 29.292 ;
			RECT	44.315 29.228 44.347 29.292 ;
			RECT	44.483 29.228 44.515 29.292 ;
			RECT	44.651 29.228 44.683 29.292 ;
			RECT	44.819 29.228 44.851 29.292 ;
			RECT	44.987 29.228 45.019 29.292 ;
			RECT	45.155 29.228 45.187 29.292 ;
			RECT	45.323 29.228 45.355 29.292 ;
			RECT	45.491 29.228 45.523 29.292 ;
			RECT	45.659 29.228 45.691 29.292 ;
			RECT	45.827 29.228 45.859 29.292 ;
			RECT	45.995 29.228 46.027 29.292 ;
			RECT	46.163 29.228 46.195 29.292 ;
			RECT	46.331 29.228 46.363 29.292 ;
			RECT	46.499 29.228 46.531 29.292 ;
			RECT	46.667 29.228 46.699 29.292 ;
			RECT	46.835 29.228 46.867 29.292 ;
			RECT	47.003 29.228 47.035 29.292 ;
			RECT	47.171 29.228 47.203 29.292 ;
			RECT	47.339 29.228 47.371 29.292 ;
			RECT	47.507 29.228 47.539 29.292 ;
			RECT	47.675 29.228 47.707 29.292 ;
			RECT	47.843 29.228 47.875 29.292 ;
			RECT	48.011 29.228 48.043 29.292 ;
			RECT	48.179 29.228 48.211 29.292 ;
			RECT	48.347 29.228 48.379 29.292 ;
			RECT	48.515 29.228 48.547 29.292 ;
			RECT	48.683 29.228 48.715 29.292 ;
			RECT	48.851 29.228 48.883 29.292 ;
			RECT	49.019 29.228 49.051 29.292 ;
			RECT	49.187 29.228 49.219 29.292 ;
			RECT	49.318 29.244 49.35 29.276 ;
			RECT	49.439 29.244 49.471 29.276 ;
			RECT	49.569 29.228 49.601 29.292 ;
			RECT	51.881 29.228 51.913 29.292 ;
			RECT	53.132 29.228 53.196 29.292 ;
			RECT	53.812 29.228 53.844 29.292 ;
			RECT	54.251 29.228 54.283 29.292 ;
			RECT	55.562 29.228 55.626 29.292 ;
			RECT	58.603 29.228 58.635 29.292 ;
			RECT	58.733 29.244 58.765 29.276 ;
			RECT	58.854 29.244 58.886 29.276 ;
			RECT	58.985 29.228 59.017 29.292 ;
			RECT	59.153 29.228 59.185 29.292 ;
			RECT	59.321 29.228 59.353 29.292 ;
			RECT	59.489 29.228 59.521 29.292 ;
			RECT	59.657 29.228 59.689 29.292 ;
			RECT	59.825 29.228 59.857 29.292 ;
			RECT	59.993 29.228 60.025 29.292 ;
			RECT	60.161 29.228 60.193 29.292 ;
			RECT	60.329 29.228 60.361 29.292 ;
			RECT	60.497 29.228 60.529 29.292 ;
			RECT	60.665 29.228 60.697 29.292 ;
			RECT	60.833 29.228 60.865 29.292 ;
			RECT	61.001 29.228 61.033 29.292 ;
			RECT	61.169 29.228 61.201 29.292 ;
			RECT	61.337 29.228 61.369 29.292 ;
			RECT	61.505 29.228 61.537 29.292 ;
			RECT	61.673 29.228 61.705 29.292 ;
			RECT	61.841 29.228 61.873 29.292 ;
			RECT	62.009 29.228 62.041 29.292 ;
			RECT	62.177 29.228 62.209 29.292 ;
			RECT	62.345 29.228 62.377 29.292 ;
			RECT	62.513 29.228 62.545 29.292 ;
			RECT	62.681 29.228 62.713 29.292 ;
			RECT	62.849 29.228 62.881 29.292 ;
			RECT	63.017 29.228 63.049 29.292 ;
			RECT	63.185 29.228 63.217 29.292 ;
			RECT	63.353 29.228 63.385 29.292 ;
			RECT	63.521 29.228 63.553 29.292 ;
			RECT	63.689 29.228 63.721 29.292 ;
			RECT	63.857 29.228 63.889 29.292 ;
			RECT	64.025 29.228 64.057 29.292 ;
			RECT	64.193 29.228 64.225 29.292 ;
			RECT	64.361 29.228 64.393 29.292 ;
			RECT	64.529 29.228 64.561 29.292 ;
			RECT	64.697 29.228 64.729 29.292 ;
			RECT	64.865 29.228 64.897 29.292 ;
			RECT	65.033 29.228 65.065 29.292 ;
			RECT	65.201 29.228 65.233 29.292 ;
			RECT	65.369 29.228 65.401 29.292 ;
			RECT	65.537 29.228 65.569 29.292 ;
			RECT	65.705 29.228 65.737 29.292 ;
			RECT	65.873 29.228 65.905 29.292 ;
			RECT	66.041 29.228 66.073 29.292 ;
			RECT	66.209 29.228 66.241 29.292 ;
			RECT	66.377 29.228 66.409 29.292 ;
			RECT	66.545 29.228 66.577 29.292 ;
			RECT	66.713 29.228 66.745 29.292 ;
			RECT	66.881 29.228 66.913 29.292 ;
			RECT	67.049 29.228 67.081 29.292 ;
			RECT	67.217 29.228 67.249 29.292 ;
			RECT	67.385 29.228 67.417 29.292 ;
			RECT	67.553 29.228 67.585 29.292 ;
			RECT	67.721 29.228 67.753 29.292 ;
			RECT	67.889 29.228 67.921 29.292 ;
			RECT	68.057 29.228 68.089 29.292 ;
			RECT	68.225 29.228 68.257 29.292 ;
			RECT	68.393 29.228 68.425 29.292 ;
			RECT	68.561 29.228 68.593 29.292 ;
			RECT	68.729 29.228 68.761 29.292 ;
			RECT	68.897 29.228 68.929 29.292 ;
			RECT	69.065 29.228 69.097 29.292 ;
			RECT	69.233 29.228 69.265 29.292 ;
			RECT	69.401 29.228 69.433 29.292 ;
			RECT	69.569 29.228 69.601 29.292 ;
			RECT	69.737 29.228 69.769 29.292 ;
			RECT	69.905 29.228 69.937 29.292 ;
			RECT	70.073 29.228 70.105 29.292 ;
			RECT	70.241 29.228 70.273 29.292 ;
			RECT	70.409 29.228 70.441 29.292 ;
			RECT	70.577 29.228 70.609 29.292 ;
			RECT	70.745 29.228 70.777 29.292 ;
			RECT	70.913 29.228 70.945 29.292 ;
			RECT	71.081 29.228 71.113 29.292 ;
			RECT	71.249 29.228 71.281 29.292 ;
			RECT	71.417 29.228 71.449 29.292 ;
			RECT	71.585 29.228 71.617 29.292 ;
			RECT	71.753 29.228 71.785 29.292 ;
			RECT	71.921 29.228 71.953 29.292 ;
			RECT	72.089 29.228 72.121 29.292 ;
			RECT	72.257 29.228 72.289 29.292 ;
			RECT	72.425 29.228 72.457 29.292 ;
			RECT	72.593 29.228 72.625 29.292 ;
			RECT	72.761 29.228 72.793 29.292 ;
			RECT	72.929 29.228 72.961 29.292 ;
			RECT	73.097 29.228 73.129 29.292 ;
			RECT	73.265 29.228 73.297 29.292 ;
			RECT	73.433 29.228 73.465 29.292 ;
			RECT	73.601 29.228 73.633 29.292 ;
			RECT	73.769 29.228 73.801 29.292 ;
			RECT	73.937 29.228 73.969 29.292 ;
			RECT	74.105 29.228 74.137 29.292 ;
			RECT	74.273 29.228 74.305 29.292 ;
			RECT	74.441 29.228 74.473 29.292 ;
			RECT	74.609 29.228 74.641 29.292 ;
			RECT	74.777 29.228 74.809 29.292 ;
			RECT	74.945 29.228 74.977 29.292 ;
			RECT	75.113 29.228 75.145 29.292 ;
			RECT	75.281 29.228 75.313 29.292 ;
			RECT	75.449 29.228 75.481 29.292 ;
			RECT	75.617 29.228 75.649 29.292 ;
			RECT	75.785 29.228 75.817 29.292 ;
			RECT	75.953 29.228 75.985 29.292 ;
			RECT	76.121 29.228 76.153 29.292 ;
			RECT	76.289 29.228 76.321 29.292 ;
			RECT	76.457 29.228 76.489 29.292 ;
			RECT	76.625 29.228 76.657 29.292 ;
			RECT	76.793 29.228 76.825 29.292 ;
			RECT	76.961 29.228 76.993 29.292 ;
			RECT	77.129 29.228 77.161 29.292 ;
			RECT	77.297 29.228 77.329 29.292 ;
			RECT	77.465 29.228 77.497 29.292 ;
			RECT	77.633 29.228 77.665 29.292 ;
			RECT	77.801 29.228 77.833 29.292 ;
			RECT	77.969 29.228 78.001 29.292 ;
			RECT	78.137 29.228 78.169 29.292 ;
			RECT	78.305 29.228 78.337 29.292 ;
			RECT	78.473 29.228 78.505 29.292 ;
			RECT	78.641 29.228 78.673 29.292 ;
			RECT	78.809 29.228 78.841 29.292 ;
			RECT	78.977 29.228 79.009 29.292 ;
			RECT	79.145 29.228 79.177 29.292 ;
			RECT	79.313 29.228 79.345 29.292 ;
			RECT	79.481 29.228 79.513 29.292 ;
			RECT	79.649 29.228 79.681 29.292 ;
			RECT	79.817 29.228 79.849 29.292 ;
			RECT	79.985 29.228 80.017 29.292 ;
			RECT	80.153 29.228 80.185 29.292 ;
			RECT	80.321 29.228 80.353 29.292 ;
			RECT	80.489 29.228 80.521 29.292 ;
			RECT	80.657 29.228 80.689 29.292 ;
			RECT	80.825 29.228 80.857 29.292 ;
			RECT	80.993 29.228 81.025 29.292 ;
			RECT	81.161 29.228 81.193 29.292 ;
			RECT	81.329 29.228 81.361 29.292 ;
			RECT	81.497 29.228 81.529 29.292 ;
			RECT	81.665 29.228 81.697 29.292 ;
			RECT	81.833 29.228 81.865 29.292 ;
			RECT	82.001 29.228 82.033 29.292 ;
			RECT	82.169 29.228 82.201 29.292 ;
			RECT	82.337 29.228 82.369 29.292 ;
			RECT	82.505 29.228 82.537 29.292 ;
			RECT	82.673 29.228 82.705 29.292 ;
			RECT	82.841 29.228 82.873 29.292 ;
			RECT	83.009 29.228 83.041 29.292 ;
			RECT	83.177 29.228 83.209 29.292 ;
			RECT	83.345 29.228 83.377 29.292 ;
			RECT	83.513 29.228 83.545 29.292 ;
			RECT	83.681 29.228 83.713 29.292 ;
			RECT	83.849 29.228 83.881 29.292 ;
			RECT	84.017 29.228 84.049 29.292 ;
			RECT	84.185 29.228 84.217 29.292 ;
			RECT	84.353 29.228 84.385 29.292 ;
			RECT	84.521 29.228 84.553 29.292 ;
			RECT	84.689 29.228 84.721 29.292 ;
			RECT	84.857 29.228 84.889 29.292 ;
			RECT	85.025 29.228 85.057 29.292 ;
			RECT	85.193 29.228 85.225 29.292 ;
			RECT	85.361 29.228 85.393 29.292 ;
			RECT	85.529 29.228 85.561 29.292 ;
			RECT	85.697 29.228 85.729 29.292 ;
			RECT	85.865 29.228 85.897 29.292 ;
			RECT	86.033 29.228 86.065 29.292 ;
			RECT	86.201 29.228 86.233 29.292 ;
			RECT	86.369 29.228 86.401 29.292 ;
			RECT	86.537 29.228 86.569 29.292 ;
			RECT	86.705 29.228 86.737 29.292 ;
			RECT	86.873 29.228 86.905 29.292 ;
			RECT	87.041 29.228 87.073 29.292 ;
			RECT	87.209 29.228 87.241 29.292 ;
			RECT	87.377 29.228 87.409 29.292 ;
			RECT	87.545 29.228 87.577 29.292 ;
			RECT	87.713 29.228 87.745 29.292 ;
			RECT	87.881 29.228 87.913 29.292 ;
			RECT	88.049 29.228 88.081 29.292 ;
			RECT	88.217 29.228 88.249 29.292 ;
			RECT	88.385 29.228 88.417 29.292 ;
			RECT	88.553 29.228 88.585 29.292 ;
			RECT	88.721 29.228 88.753 29.292 ;
			RECT	88.889 29.228 88.921 29.292 ;
			RECT	89.057 29.228 89.089 29.292 ;
			RECT	89.225 29.228 89.257 29.292 ;
			RECT	89.393 29.228 89.425 29.292 ;
			RECT	89.561 29.228 89.593 29.292 ;
			RECT	89.729 29.228 89.761 29.292 ;
			RECT	89.897 29.228 89.929 29.292 ;
			RECT	90.065 29.228 90.097 29.292 ;
			RECT	90.233 29.228 90.265 29.292 ;
			RECT	90.401 29.228 90.433 29.292 ;
			RECT	90.569 29.228 90.601 29.292 ;
			RECT	90.737 29.228 90.769 29.292 ;
			RECT	90.905 29.228 90.937 29.292 ;
			RECT	91.073 29.228 91.105 29.292 ;
			RECT	91.241 29.228 91.273 29.292 ;
			RECT	91.409 29.228 91.441 29.292 ;
			RECT	91.577 29.228 91.609 29.292 ;
			RECT	91.745 29.228 91.777 29.292 ;
			RECT	91.913 29.228 91.945 29.292 ;
			RECT	92.081 29.228 92.113 29.292 ;
			RECT	92.249 29.228 92.281 29.292 ;
			RECT	92.417 29.228 92.449 29.292 ;
			RECT	92.585 29.228 92.617 29.292 ;
			RECT	92.753 29.228 92.785 29.292 ;
			RECT	92.921 29.228 92.953 29.292 ;
			RECT	93.089 29.228 93.121 29.292 ;
			RECT	93.257 29.228 93.289 29.292 ;
			RECT	93.425 29.228 93.457 29.292 ;
			RECT	93.593 29.228 93.625 29.292 ;
			RECT	93.761 29.228 93.793 29.292 ;
			RECT	93.929 29.228 93.961 29.292 ;
			RECT	94.097 29.228 94.129 29.292 ;
			RECT	94.265 29.228 94.297 29.292 ;
			RECT	94.433 29.228 94.465 29.292 ;
			RECT	94.601 29.228 94.633 29.292 ;
			RECT	94.769 29.228 94.801 29.292 ;
			RECT	94.937 29.228 94.969 29.292 ;
			RECT	95.105 29.228 95.137 29.292 ;
			RECT	95.273 29.228 95.305 29.292 ;
			RECT	95.441 29.228 95.473 29.292 ;
			RECT	95.609 29.228 95.641 29.292 ;
			RECT	95.777 29.228 95.809 29.292 ;
			RECT	95.945 29.228 95.977 29.292 ;
			RECT	96.113 29.228 96.145 29.292 ;
			RECT	96.281 29.228 96.313 29.292 ;
			RECT	96.449 29.228 96.481 29.292 ;
			RECT	96.617 29.228 96.649 29.292 ;
			RECT	96.785 29.228 96.817 29.292 ;
			RECT	96.953 29.228 96.985 29.292 ;
			RECT	97.121 29.228 97.153 29.292 ;
			RECT	97.289 29.228 97.321 29.292 ;
			RECT	97.457 29.228 97.489 29.292 ;
			RECT	97.625 29.228 97.657 29.292 ;
			RECT	97.793 29.228 97.825 29.292 ;
			RECT	97.961 29.228 97.993 29.292 ;
			RECT	98.129 29.228 98.161 29.292 ;
			RECT	98.297 29.228 98.329 29.292 ;
			RECT	98.465 29.228 98.497 29.292 ;
			RECT	98.633 29.228 98.665 29.292 ;
			RECT	98.801 29.228 98.833 29.292 ;
			RECT	98.969 29.228 99.001 29.292 ;
			RECT	99.137 29.228 99.169 29.292 ;
			RECT	99.305 29.228 99.337 29.292 ;
			RECT	99.473 29.228 99.505 29.292 ;
			RECT	99.641 29.228 99.673 29.292 ;
			RECT	99.809 29.228 99.841 29.292 ;
			RECT	99.977 29.228 100.009 29.292 ;
			RECT	100.145 29.228 100.177 29.292 ;
			RECT	100.313 29.228 100.345 29.292 ;
			RECT	100.481 29.228 100.513 29.292 ;
			RECT	100.649 29.228 100.681 29.292 ;
			RECT	100.817 29.228 100.849 29.292 ;
			RECT	100.985 29.228 101.017 29.292 ;
			RECT	101.153 29.228 101.185 29.292 ;
			RECT	101.321 29.228 101.353 29.292 ;
			RECT	101.489 29.228 101.521 29.292 ;
			RECT	101.657 29.228 101.689 29.292 ;
			RECT	101.825 29.228 101.857 29.292 ;
			RECT	101.993 29.228 102.025 29.292 ;
			RECT	102.123 29.244 102.155 29.276 ;
			RECT	102.245 29.249 102.277 29.281 ;
			RECT	102.375 29.228 102.407 29.292 ;
			RECT	103.795 29.228 103.827 29.292 ;
			RECT	103.925 29.249 103.957 29.281 ;
			RECT	104.047 29.244 104.079 29.276 ;
			RECT	104.177 29.228 104.209 29.292 ;
			RECT	104.345 29.228 104.377 29.292 ;
			RECT	104.513 29.228 104.545 29.292 ;
			RECT	104.681 29.228 104.713 29.292 ;
			RECT	104.849 29.228 104.881 29.292 ;
			RECT	105.017 29.228 105.049 29.292 ;
			RECT	105.185 29.228 105.217 29.292 ;
			RECT	105.353 29.228 105.385 29.292 ;
			RECT	105.521 29.228 105.553 29.292 ;
			RECT	105.689 29.228 105.721 29.292 ;
			RECT	105.857 29.228 105.889 29.292 ;
			RECT	106.025 29.228 106.057 29.292 ;
			RECT	106.193 29.228 106.225 29.292 ;
			RECT	106.361 29.228 106.393 29.292 ;
			RECT	106.529 29.228 106.561 29.292 ;
			RECT	106.697 29.228 106.729 29.292 ;
			RECT	106.865 29.228 106.897 29.292 ;
			RECT	107.033 29.228 107.065 29.292 ;
			RECT	107.201 29.228 107.233 29.292 ;
			RECT	107.369 29.228 107.401 29.292 ;
			RECT	107.537 29.228 107.569 29.292 ;
			RECT	107.705 29.228 107.737 29.292 ;
			RECT	107.873 29.228 107.905 29.292 ;
			RECT	108.041 29.228 108.073 29.292 ;
			RECT	108.209 29.228 108.241 29.292 ;
			RECT	108.377 29.228 108.409 29.292 ;
			RECT	108.545 29.228 108.577 29.292 ;
			RECT	108.713 29.228 108.745 29.292 ;
			RECT	108.881 29.228 108.913 29.292 ;
			RECT	109.049 29.228 109.081 29.292 ;
			RECT	109.217 29.228 109.249 29.292 ;
			RECT	109.385 29.228 109.417 29.292 ;
			RECT	109.553 29.228 109.585 29.292 ;
			RECT	109.721 29.228 109.753 29.292 ;
			RECT	109.889 29.228 109.921 29.292 ;
			RECT	110.057 29.228 110.089 29.292 ;
			RECT	110.225 29.228 110.257 29.292 ;
			RECT	110.393 29.228 110.425 29.292 ;
			RECT	110.561 29.228 110.593 29.292 ;
			RECT	110.729 29.228 110.761 29.292 ;
			RECT	110.897 29.228 110.929 29.292 ;
			RECT	111.065 29.228 111.097 29.292 ;
			RECT	111.233 29.228 111.265 29.292 ;
			RECT	111.401 29.228 111.433 29.292 ;
			RECT	111.569 29.228 111.601 29.292 ;
			RECT	111.737 29.228 111.769 29.292 ;
			RECT	111.905 29.228 111.937 29.292 ;
			RECT	112.073 29.228 112.105 29.292 ;
			RECT	112.241 29.228 112.273 29.292 ;
			RECT	112.409 29.228 112.441 29.292 ;
			RECT	112.577 29.228 112.609 29.292 ;
			RECT	112.745 29.228 112.777 29.292 ;
			RECT	112.913 29.228 112.945 29.292 ;
			RECT	113.081 29.228 113.113 29.292 ;
			RECT	113.249 29.228 113.281 29.292 ;
			RECT	113.417 29.228 113.449 29.292 ;
			RECT	113.585 29.228 113.617 29.292 ;
			RECT	113.753 29.228 113.785 29.292 ;
			RECT	113.921 29.228 113.953 29.292 ;
			RECT	114.089 29.228 114.121 29.292 ;
			RECT	114.257 29.228 114.289 29.292 ;
			RECT	114.425 29.228 114.457 29.292 ;
			RECT	114.593 29.228 114.625 29.292 ;
			RECT	114.761 29.228 114.793 29.292 ;
			RECT	114.929 29.228 114.961 29.292 ;
			RECT	115.097 29.228 115.129 29.292 ;
			RECT	115.265 29.228 115.297 29.292 ;
			RECT	115.433 29.228 115.465 29.292 ;
			RECT	115.601 29.228 115.633 29.292 ;
			RECT	115.769 29.228 115.801 29.292 ;
			RECT	115.937 29.228 115.969 29.292 ;
			RECT	116.105 29.228 116.137 29.292 ;
			RECT	116.273 29.228 116.305 29.292 ;
			RECT	116.441 29.228 116.473 29.292 ;
			RECT	116.609 29.228 116.641 29.292 ;
			RECT	116.777 29.228 116.809 29.292 ;
			RECT	116.945 29.228 116.977 29.292 ;
			RECT	117.113 29.228 117.145 29.292 ;
			RECT	117.281 29.228 117.313 29.292 ;
			RECT	117.449 29.228 117.481 29.292 ;
			RECT	117.617 29.228 117.649 29.292 ;
			RECT	117.785 29.228 117.817 29.292 ;
			RECT	117.953 29.228 117.985 29.292 ;
			RECT	118.121 29.228 118.153 29.292 ;
			RECT	118.289 29.228 118.321 29.292 ;
			RECT	118.457 29.228 118.489 29.292 ;
			RECT	118.625 29.228 118.657 29.292 ;
			RECT	118.793 29.228 118.825 29.292 ;
			RECT	118.961 29.228 118.993 29.292 ;
			RECT	119.129 29.228 119.161 29.292 ;
			RECT	119.297 29.228 119.329 29.292 ;
			RECT	119.465 29.228 119.497 29.292 ;
			RECT	119.633 29.228 119.665 29.292 ;
			RECT	119.801 29.228 119.833 29.292 ;
			RECT	119.969 29.228 120.001 29.292 ;
			RECT	120.137 29.228 120.169 29.292 ;
			RECT	120.305 29.228 120.337 29.292 ;
			RECT	120.473 29.228 120.505 29.292 ;
			RECT	120.641 29.228 120.673 29.292 ;
			RECT	120.809 29.228 120.841 29.292 ;
			RECT	120.977 29.228 121.009 29.292 ;
			RECT	121.145 29.228 121.177 29.292 ;
			RECT	121.313 29.228 121.345 29.292 ;
			RECT	121.481 29.228 121.513 29.292 ;
			RECT	121.649 29.228 121.681 29.292 ;
			RECT	121.817 29.228 121.849 29.292 ;
			RECT	121.985 29.228 122.017 29.292 ;
			RECT	122.153 29.228 122.185 29.292 ;
			RECT	122.321 29.228 122.353 29.292 ;
			RECT	122.489 29.228 122.521 29.292 ;
			RECT	122.657 29.228 122.689 29.292 ;
			RECT	122.825 29.228 122.857 29.292 ;
			RECT	122.993 29.228 123.025 29.292 ;
			RECT	123.161 29.228 123.193 29.292 ;
			RECT	123.329 29.228 123.361 29.292 ;
			RECT	123.497 29.228 123.529 29.292 ;
			RECT	123.665 29.228 123.697 29.292 ;
			RECT	123.833 29.228 123.865 29.292 ;
			RECT	124.001 29.228 124.033 29.292 ;
			RECT	124.169 29.228 124.201 29.292 ;
			RECT	124.337 29.228 124.369 29.292 ;
			RECT	124.505 29.228 124.537 29.292 ;
			RECT	124.673 29.228 124.705 29.292 ;
			RECT	124.841 29.228 124.873 29.292 ;
			RECT	125.009 29.228 125.041 29.292 ;
			RECT	125.177 29.228 125.209 29.292 ;
			RECT	125.345 29.228 125.377 29.292 ;
			RECT	125.513 29.228 125.545 29.292 ;
			RECT	125.681 29.228 125.713 29.292 ;
			RECT	125.849 29.228 125.881 29.292 ;
			RECT	126.017 29.228 126.049 29.292 ;
			RECT	126.185 29.228 126.217 29.292 ;
			RECT	126.353 29.228 126.385 29.292 ;
			RECT	126.521 29.228 126.553 29.292 ;
			RECT	126.689 29.228 126.721 29.292 ;
			RECT	126.857 29.228 126.889 29.292 ;
			RECT	127.025 29.228 127.057 29.292 ;
			RECT	127.193 29.228 127.225 29.292 ;
			RECT	127.361 29.228 127.393 29.292 ;
			RECT	127.529 29.228 127.561 29.292 ;
			RECT	127.697 29.228 127.729 29.292 ;
			RECT	127.865 29.228 127.897 29.292 ;
			RECT	128.033 29.228 128.065 29.292 ;
			RECT	128.201 29.228 128.233 29.292 ;
			RECT	128.369 29.228 128.401 29.292 ;
			RECT	128.537 29.228 128.569 29.292 ;
			RECT	128.705 29.228 128.737 29.292 ;
			RECT	128.873 29.228 128.905 29.292 ;
			RECT	129.041 29.228 129.073 29.292 ;
			RECT	129.209 29.228 129.241 29.292 ;
			RECT	129.377 29.228 129.409 29.292 ;
			RECT	129.545 29.228 129.577 29.292 ;
			RECT	129.713 29.228 129.745 29.292 ;
			RECT	129.881 29.228 129.913 29.292 ;
			RECT	130.049 29.228 130.081 29.292 ;
			RECT	130.217 29.228 130.249 29.292 ;
			RECT	130.385 29.228 130.417 29.292 ;
			RECT	130.553 29.228 130.585 29.292 ;
			RECT	130.721 29.228 130.753 29.292 ;
			RECT	130.889 29.228 130.921 29.292 ;
			RECT	131.057 29.228 131.089 29.292 ;
			RECT	131.225 29.228 131.257 29.292 ;
			RECT	131.393 29.228 131.425 29.292 ;
			RECT	131.561 29.228 131.593 29.292 ;
			RECT	131.729 29.228 131.761 29.292 ;
			RECT	131.897 29.228 131.929 29.292 ;
			RECT	132.065 29.228 132.097 29.292 ;
			RECT	132.233 29.228 132.265 29.292 ;
			RECT	132.401 29.228 132.433 29.292 ;
			RECT	132.569 29.228 132.601 29.292 ;
			RECT	132.737 29.228 132.769 29.292 ;
			RECT	132.905 29.228 132.937 29.292 ;
			RECT	133.073 29.228 133.105 29.292 ;
			RECT	133.241 29.228 133.273 29.292 ;
			RECT	133.409 29.228 133.441 29.292 ;
			RECT	133.577 29.228 133.609 29.292 ;
			RECT	133.745 29.228 133.777 29.292 ;
			RECT	133.913 29.228 133.945 29.292 ;
			RECT	134.081 29.228 134.113 29.292 ;
			RECT	134.249 29.228 134.281 29.292 ;
			RECT	134.417 29.228 134.449 29.292 ;
			RECT	134.585 29.228 134.617 29.292 ;
			RECT	134.753 29.228 134.785 29.292 ;
			RECT	134.921 29.228 134.953 29.292 ;
			RECT	135.089 29.228 135.121 29.292 ;
			RECT	135.257 29.228 135.289 29.292 ;
			RECT	135.425 29.228 135.457 29.292 ;
			RECT	135.593 29.228 135.625 29.292 ;
			RECT	135.761 29.228 135.793 29.292 ;
			RECT	135.929 29.228 135.961 29.292 ;
			RECT	136.097 29.228 136.129 29.292 ;
			RECT	136.265 29.228 136.297 29.292 ;
			RECT	136.433 29.228 136.465 29.292 ;
			RECT	136.601 29.228 136.633 29.292 ;
			RECT	136.769 29.228 136.801 29.292 ;
			RECT	136.937 29.228 136.969 29.292 ;
			RECT	137.105 29.228 137.137 29.292 ;
			RECT	137.273 29.228 137.305 29.292 ;
			RECT	137.441 29.228 137.473 29.292 ;
			RECT	137.609 29.228 137.641 29.292 ;
			RECT	137.777 29.228 137.809 29.292 ;
			RECT	137.945 29.228 137.977 29.292 ;
			RECT	138.113 29.228 138.145 29.292 ;
			RECT	138.281 29.228 138.313 29.292 ;
			RECT	138.449 29.228 138.481 29.292 ;
			RECT	138.617 29.228 138.649 29.292 ;
			RECT	138.785 29.228 138.817 29.292 ;
			RECT	138.953 29.228 138.985 29.292 ;
			RECT	139.121 29.228 139.153 29.292 ;
			RECT	139.289 29.228 139.321 29.292 ;
			RECT	139.457 29.228 139.489 29.292 ;
			RECT	139.625 29.228 139.657 29.292 ;
			RECT	139.793 29.228 139.825 29.292 ;
			RECT	139.961 29.228 139.993 29.292 ;
			RECT	140.129 29.228 140.161 29.292 ;
			RECT	140.297 29.228 140.329 29.292 ;
			RECT	140.465 29.228 140.497 29.292 ;
			RECT	140.633 29.228 140.665 29.292 ;
			RECT	140.801 29.228 140.833 29.292 ;
			RECT	140.969 29.228 141.001 29.292 ;
			RECT	141.137 29.228 141.169 29.292 ;
			RECT	141.305 29.228 141.337 29.292 ;
			RECT	141.473 29.228 141.505 29.292 ;
			RECT	141.641 29.228 141.673 29.292 ;
			RECT	141.809 29.228 141.841 29.292 ;
			RECT	141.977 29.228 142.009 29.292 ;
			RECT	142.145 29.228 142.177 29.292 ;
			RECT	142.313 29.228 142.345 29.292 ;
			RECT	142.481 29.228 142.513 29.292 ;
			RECT	142.649 29.228 142.681 29.292 ;
			RECT	142.817 29.228 142.849 29.292 ;
			RECT	142.985 29.228 143.017 29.292 ;
			RECT	143.153 29.228 143.185 29.292 ;
			RECT	143.321 29.228 143.353 29.292 ;
			RECT	143.489 29.228 143.521 29.292 ;
			RECT	143.657 29.228 143.689 29.292 ;
			RECT	143.825 29.228 143.857 29.292 ;
			RECT	143.993 29.228 144.025 29.292 ;
			RECT	144.161 29.228 144.193 29.292 ;
			RECT	144.329 29.228 144.361 29.292 ;
			RECT	144.497 29.228 144.529 29.292 ;
			RECT	144.665 29.228 144.697 29.292 ;
			RECT	144.833 29.228 144.865 29.292 ;
			RECT	145.001 29.228 145.033 29.292 ;
			RECT	145.169 29.228 145.201 29.292 ;
			RECT	145.337 29.228 145.369 29.292 ;
			RECT	145.505 29.228 145.537 29.292 ;
			RECT	145.673 29.228 145.705 29.292 ;
			RECT	145.841 29.228 145.873 29.292 ;
			RECT	146.009 29.228 146.041 29.292 ;
			RECT	146.177 29.228 146.209 29.292 ;
			RECT	146.345 29.228 146.377 29.292 ;
			RECT	146.513 29.228 146.545 29.292 ;
			RECT	146.681 29.228 146.713 29.292 ;
			RECT	146.849 29.228 146.881 29.292 ;
			RECT	147.017 29.228 147.049 29.292 ;
			RECT	147.185 29.228 147.217 29.292 ;
			RECT	147.316 29.244 147.348 29.276 ;
			RECT	147.437 29.244 147.469 29.276 ;
			RECT	147.567 29.228 147.599 29.292 ;
			RECT	149.879 29.228 149.911 29.292 ;
			RECT	151.13 29.228 151.194 29.292 ;
			RECT	151.81 29.228 151.842 29.292 ;
			RECT	152.249 29.228 152.281 29.292 ;
			RECT	153.56 29.228 153.624 29.292 ;
			RECT	156.601 29.228 156.633 29.292 ;
			RECT	156.731 29.244 156.763 29.276 ;
			RECT	156.852 29.244 156.884 29.276 ;
			RECT	156.983 29.228 157.015 29.292 ;
			RECT	157.151 29.228 157.183 29.292 ;
			RECT	157.319 29.228 157.351 29.292 ;
			RECT	157.487 29.228 157.519 29.292 ;
			RECT	157.655 29.228 157.687 29.292 ;
			RECT	157.823 29.228 157.855 29.292 ;
			RECT	157.991 29.228 158.023 29.292 ;
			RECT	158.159 29.228 158.191 29.292 ;
			RECT	158.327 29.228 158.359 29.292 ;
			RECT	158.495 29.228 158.527 29.292 ;
			RECT	158.663 29.228 158.695 29.292 ;
			RECT	158.831 29.228 158.863 29.292 ;
			RECT	158.999 29.228 159.031 29.292 ;
			RECT	159.167 29.228 159.199 29.292 ;
			RECT	159.335 29.228 159.367 29.292 ;
			RECT	159.503 29.228 159.535 29.292 ;
			RECT	159.671 29.228 159.703 29.292 ;
			RECT	159.839 29.228 159.871 29.292 ;
			RECT	160.007 29.228 160.039 29.292 ;
			RECT	160.175 29.228 160.207 29.292 ;
			RECT	160.343 29.228 160.375 29.292 ;
			RECT	160.511 29.228 160.543 29.292 ;
			RECT	160.679 29.228 160.711 29.292 ;
			RECT	160.847 29.228 160.879 29.292 ;
			RECT	161.015 29.228 161.047 29.292 ;
			RECT	161.183 29.228 161.215 29.292 ;
			RECT	161.351 29.228 161.383 29.292 ;
			RECT	161.519 29.228 161.551 29.292 ;
			RECT	161.687 29.228 161.719 29.292 ;
			RECT	161.855 29.228 161.887 29.292 ;
			RECT	162.023 29.228 162.055 29.292 ;
			RECT	162.191 29.228 162.223 29.292 ;
			RECT	162.359 29.228 162.391 29.292 ;
			RECT	162.527 29.228 162.559 29.292 ;
			RECT	162.695 29.228 162.727 29.292 ;
			RECT	162.863 29.228 162.895 29.292 ;
			RECT	163.031 29.228 163.063 29.292 ;
			RECT	163.199 29.228 163.231 29.292 ;
			RECT	163.367 29.228 163.399 29.292 ;
			RECT	163.535 29.228 163.567 29.292 ;
			RECT	163.703 29.228 163.735 29.292 ;
			RECT	163.871 29.228 163.903 29.292 ;
			RECT	164.039 29.228 164.071 29.292 ;
			RECT	164.207 29.228 164.239 29.292 ;
			RECT	164.375 29.228 164.407 29.292 ;
			RECT	164.543 29.228 164.575 29.292 ;
			RECT	164.711 29.228 164.743 29.292 ;
			RECT	164.879 29.228 164.911 29.292 ;
			RECT	165.047 29.228 165.079 29.292 ;
			RECT	165.215 29.228 165.247 29.292 ;
			RECT	165.383 29.228 165.415 29.292 ;
			RECT	165.551 29.228 165.583 29.292 ;
			RECT	165.719 29.228 165.751 29.292 ;
			RECT	165.887 29.228 165.919 29.292 ;
			RECT	166.055 29.228 166.087 29.292 ;
			RECT	166.223 29.228 166.255 29.292 ;
			RECT	166.391 29.228 166.423 29.292 ;
			RECT	166.559 29.228 166.591 29.292 ;
			RECT	166.727 29.228 166.759 29.292 ;
			RECT	166.895 29.228 166.927 29.292 ;
			RECT	167.063 29.228 167.095 29.292 ;
			RECT	167.231 29.228 167.263 29.292 ;
			RECT	167.399 29.228 167.431 29.292 ;
			RECT	167.567 29.228 167.599 29.292 ;
			RECT	167.735 29.228 167.767 29.292 ;
			RECT	167.903 29.228 167.935 29.292 ;
			RECT	168.071 29.228 168.103 29.292 ;
			RECT	168.239 29.228 168.271 29.292 ;
			RECT	168.407 29.228 168.439 29.292 ;
			RECT	168.575 29.228 168.607 29.292 ;
			RECT	168.743 29.228 168.775 29.292 ;
			RECT	168.911 29.228 168.943 29.292 ;
			RECT	169.079 29.228 169.111 29.292 ;
			RECT	169.247 29.228 169.279 29.292 ;
			RECT	169.415 29.228 169.447 29.292 ;
			RECT	169.583 29.228 169.615 29.292 ;
			RECT	169.751 29.228 169.783 29.292 ;
			RECT	169.919 29.228 169.951 29.292 ;
			RECT	170.087 29.228 170.119 29.292 ;
			RECT	170.255 29.228 170.287 29.292 ;
			RECT	170.423 29.228 170.455 29.292 ;
			RECT	170.591 29.228 170.623 29.292 ;
			RECT	170.759 29.228 170.791 29.292 ;
			RECT	170.927 29.228 170.959 29.292 ;
			RECT	171.095 29.228 171.127 29.292 ;
			RECT	171.263 29.228 171.295 29.292 ;
			RECT	171.431 29.228 171.463 29.292 ;
			RECT	171.599 29.228 171.631 29.292 ;
			RECT	171.767 29.228 171.799 29.292 ;
			RECT	171.935 29.228 171.967 29.292 ;
			RECT	172.103 29.228 172.135 29.292 ;
			RECT	172.271 29.228 172.303 29.292 ;
			RECT	172.439 29.228 172.471 29.292 ;
			RECT	172.607 29.228 172.639 29.292 ;
			RECT	172.775 29.228 172.807 29.292 ;
			RECT	172.943 29.228 172.975 29.292 ;
			RECT	173.111 29.228 173.143 29.292 ;
			RECT	173.279 29.228 173.311 29.292 ;
			RECT	173.447 29.228 173.479 29.292 ;
			RECT	173.615 29.228 173.647 29.292 ;
			RECT	173.783 29.228 173.815 29.292 ;
			RECT	173.951 29.228 173.983 29.292 ;
			RECT	174.119 29.228 174.151 29.292 ;
			RECT	174.287 29.228 174.319 29.292 ;
			RECT	174.455 29.228 174.487 29.292 ;
			RECT	174.623 29.228 174.655 29.292 ;
			RECT	174.791 29.228 174.823 29.292 ;
			RECT	174.959 29.228 174.991 29.292 ;
			RECT	175.127 29.228 175.159 29.292 ;
			RECT	175.295 29.228 175.327 29.292 ;
			RECT	175.463 29.228 175.495 29.292 ;
			RECT	175.631 29.228 175.663 29.292 ;
			RECT	175.799 29.228 175.831 29.292 ;
			RECT	175.967 29.228 175.999 29.292 ;
			RECT	176.135 29.228 176.167 29.292 ;
			RECT	176.303 29.228 176.335 29.292 ;
			RECT	176.471 29.228 176.503 29.292 ;
			RECT	176.639 29.228 176.671 29.292 ;
			RECT	176.807 29.228 176.839 29.292 ;
			RECT	176.975 29.228 177.007 29.292 ;
			RECT	177.143 29.228 177.175 29.292 ;
			RECT	177.311 29.228 177.343 29.292 ;
			RECT	177.479 29.228 177.511 29.292 ;
			RECT	177.647 29.228 177.679 29.292 ;
			RECT	177.815 29.228 177.847 29.292 ;
			RECT	177.983 29.228 178.015 29.292 ;
			RECT	178.151 29.228 178.183 29.292 ;
			RECT	178.319 29.228 178.351 29.292 ;
			RECT	178.487 29.228 178.519 29.292 ;
			RECT	178.655 29.228 178.687 29.292 ;
			RECT	178.823 29.228 178.855 29.292 ;
			RECT	178.991 29.228 179.023 29.292 ;
			RECT	179.159 29.228 179.191 29.292 ;
			RECT	179.327 29.228 179.359 29.292 ;
			RECT	179.495 29.228 179.527 29.292 ;
			RECT	179.663 29.228 179.695 29.292 ;
			RECT	179.831 29.228 179.863 29.292 ;
			RECT	179.999 29.228 180.031 29.292 ;
			RECT	180.167 29.228 180.199 29.292 ;
			RECT	180.335 29.228 180.367 29.292 ;
			RECT	180.503 29.228 180.535 29.292 ;
			RECT	180.671 29.228 180.703 29.292 ;
			RECT	180.839 29.228 180.871 29.292 ;
			RECT	181.007 29.228 181.039 29.292 ;
			RECT	181.175 29.228 181.207 29.292 ;
			RECT	181.343 29.228 181.375 29.292 ;
			RECT	181.511 29.228 181.543 29.292 ;
			RECT	181.679 29.228 181.711 29.292 ;
			RECT	181.847 29.228 181.879 29.292 ;
			RECT	182.015 29.228 182.047 29.292 ;
			RECT	182.183 29.228 182.215 29.292 ;
			RECT	182.351 29.228 182.383 29.292 ;
			RECT	182.519 29.228 182.551 29.292 ;
			RECT	182.687 29.228 182.719 29.292 ;
			RECT	182.855 29.228 182.887 29.292 ;
			RECT	183.023 29.228 183.055 29.292 ;
			RECT	183.191 29.228 183.223 29.292 ;
			RECT	183.359 29.228 183.391 29.292 ;
			RECT	183.527 29.228 183.559 29.292 ;
			RECT	183.695 29.228 183.727 29.292 ;
			RECT	183.863 29.228 183.895 29.292 ;
			RECT	184.031 29.228 184.063 29.292 ;
			RECT	184.199 29.228 184.231 29.292 ;
			RECT	184.367 29.228 184.399 29.292 ;
			RECT	184.535 29.228 184.567 29.292 ;
			RECT	184.703 29.228 184.735 29.292 ;
			RECT	184.871 29.228 184.903 29.292 ;
			RECT	185.039 29.228 185.071 29.292 ;
			RECT	185.207 29.228 185.239 29.292 ;
			RECT	185.375 29.228 185.407 29.292 ;
			RECT	185.543 29.228 185.575 29.292 ;
			RECT	185.711 29.228 185.743 29.292 ;
			RECT	185.879 29.228 185.911 29.292 ;
			RECT	186.047 29.228 186.079 29.292 ;
			RECT	186.215 29.228 186.247 29.292 ;
			RECT	186.383 29.228 186.415 29.292 ;
			RECT	186.551 29.228 186.583 29.292 ;
			RECT	186.719 29.228 186.751 29.292 ;
			RECT	186.887 29.228 186.919 29.292 ;
			RECT	187.055 29.228 187.087 29.292 ;
			RECT	187.223 29.228 187.255 29.292 ;
			RECT	187.391 29.228 187.423 29.292 ;
			RECT	187.559 29.228 187.591 29.292 ;
			RECT	187.727 29.228 187.759 29.292 ;
			RECT	187.895 29.228 187.927 29.292 ;
			RECT	188.063 29.228 188.095 29.292 ;
			RECT	188.231 29.228 188.263 29.292 ;
			RECT	188.399 29.228 188.431 29.292 ;
			RECT	188.567 29.228 188.599 29.292 ;
			RECT	188.735 29.228 188.767 29.292 ;
			RECT	188.903 29.228 188.935 29.292 ;
			RECT	189.071 29.228 189.103 29.292 ;
			RECT	189.239 29.228 189.271 29.292 ;
			RECT	189.407 29.228 189.439 29.292 ;
			RECT	189.575 29.228 189.607 29.292 ;
			RECT	189.743 29.228 189.775 29.292 ;
			RECT	189.911 29.228 189.943 29.292 ;
			RECT	190.079 29.228 190.111 29.292 ;
			RECT	190.247 29.228 190.279 29.292 ;
			RECT	190.415 29.228 190.447 29.292 ;
			RECT	190.583 29.228 190.615 29.292 ;
			RECT	190.751 29.228 190.783 29.292 ;
			RECT	190.919 29.228 190.951 29.292 ;
			RECT	191.087 29.228 191.119 29.292 ;
			RECT	191.255 29.228 191.287 29.292 ;
			RECT	191.423 29.228 191.455 29.292 ;
			RECT	191.591 29.228 191.623 29.292 ;
			RECT	191.759 29.228 191.791 29.292 ;
			RECT	191.927 29.228 191.959 29.292 ;
			RECT	192.095 29.228 192.127 29.292 ;
			RECT	192.263 29.228 192.295 29.292 ;
			RECT	192.431 29.228 192.463 29.292 ;
			RECT	192.599 29.228 192.631 29.292 ;
			RECT	192.767 29.228 192.799 29.292 ;
			RECT	192.935 29.228 192.967 29.292 ;
			RECT	193.103 29.228 193.135 29.292 ;
			RECT	193.271 29.228 193.303 29.292 ;
			RECT	193.439 29.228 193.471 29.292 ;
			RECT	193.607 29.228 193.639 29.292 ;
			RECT	193.775 29.228 193.807 29.292 ;
			RECT	193.943 29.228 193.975 29.292 ;
			RECT	194.111 29.228 194.143 29.292 ;
			RECT	194.279 29.228 194.311 29.292 ;
			RECT	194.447 29.228 194.479 29.292 ;
			RECT	194.615 29.228 194.647 29.292 ;
			RECT	194.783 29.228 194.815 29.292 ;
			RECT	194.951 29.228 194.983 29.292 ;
			RECT	195.119 29.228 195.151 29.292 ;
			RECT	195.287 29.228 195.319 29.292 ;
			RECT	195.455 29.228 195.487 29.292 ;
			RECT	195.623 29.228 195.655 29.292 ;
			RECT	195.791 29.228 195.823 29.292 ;
			RECT	195.959 29.228 195.991 29.292 ;
			RECT	196.127 29.228 196.159 29.292 ;
			RECT	196.295 29.228 196.327 29.292 ;
			RECT	196.463 29.228 196.495 29.292 ;
			RECT	196.631 29.228 196.663 29.292 ;
			RECT	196.799 29.228 196.831 29.292 ;
			RECT	196.967 29.228 196.999 29.292 ;
			RECT	197.135 29.228 197.167 29.292 ;
			RECT	197.303 29.228 197.335 29.292 ;
			RECT	197.471 29.228 197.503 29.292 ;
			RECT	197.639 29.228 197.671 29.292 ;
			RECT	197.807 29.228 197.839 29.292 ;
			RECT	197.975 29.228 198.007 29.292 ;
			RECT	198.143 29.228 198.175 29.292 ;
			RECT	198.311 29.228 198.343 29.292 ;
			RECT	198.479 29.228 198.511 29.292 ;
			RECT	198.647 29.228 198.679 29.292 ;
			RECT	198.815 29.228 198.847 29.292 ;
			RECT	198.983 29.228 199.015 29.292 ;
			RECT	199.151 29.228 199.183 29.292 ;
			RECT	199.319 29.228 199.351 29.292 ;
			RECT	199.487 29.228 199.519 29.292 ;
			RECT	199.655 29.228 199.687 29.292 ;
			RECT	199.823 29.228 199.855 29.292 ;
			RECT	199.991 29.228 200.023 29.292 ;
			RECT	200.121 29.244 200.153 29.276 ;
			RECT	200.243 29.249 200.275 29.281 ;
			RECT	200.373 29.228 200.405 29.292 ;
			RECT	200.9 29.228 200.932 29.292 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 75.896 201.665 76.016 ;
			LAYER	J3 ;
			RECT	0.755 75.924 0.787 75.988 ;
			RECT	1.645 75.924 1.709 75.988 ;
			RECT	2.323 75.924 2.387 75.988 ;
			RECT	3.438 75.924 3.47 75.988 ;
			RECT	3.585 75.924 3.617 75.988 ;
			RECT	4.195 75.924 4.227 75.988 ;
			RECT	4.72 75.924 4.752 75.988 ;
			RECT	4.944 75.924 5.008 75.988 ;
			RECT	5.267 75.924 5.299 75.988 ;
			RECT	5.797 75.924 5.829 75.988 ;
			RECT	5.927 75.935 5.959 75.967 ;
			RECT	6.049 75.94 6.081 75.972 ;
			RECT	6.179 75.924 6.211 75.988 ;
			RECT	6.347 75.924 6.379 75.988 ;
			RECT	6.515 75.924 6.547 75.988 ;
			RECT	6.683 75.924 6.715 75.988 ;
			RECT	6.851 75.924 6.883 75.988 ;
			RECT	7.019 75.924 7.051 75.988 ;
			RECT	7.187 75.924 7.219 75.988 ;
			RECT	7.355 75.924 7.387 75.988 ;
			RECT	7.523 75.924 7.555 75.988 ;
			RECT	7.691 75.924 7.723 75.988 ;
			RECT	7.859 75.924 7.891 75.988 ;
			RECT	8.027 75.924 8.059 75.988 ;
			RECT	8.195 75.924 8.227 75.988 ;
			RECT	8.363 75.924 8.395 75.988 ;
			RECT	8.531 75.924 8.563 75.988 ;
			RECT	8.699 75.924 8.731 75.988 ;
			RECT	8.867 75.924 8.899 75.988 ;
			RECT	9.035 75.924 9.067 75.988 ;
			RECT	9.203 75.924 9.235 75.988 ;
			RECT	9.371 75.924 9.403 75.988 ;
			RECT	9.539 75.924 9.571 75.988 ;
			RECT	9.707 75.924 9.739 75.988 ;
			RECT	9.875 75.924 9.907 75.988 ;
			RECT	10.043 75.924 10.075 75.988 ;
			RECT	10.211 75.924 10.243 75.988 ;
			RECT	10.379 75.924 10.411 75.988 ;
			RECT	10.547 75.924 10.579 75.988 ;
			RECT	10.715 75.924 10.747 75.988 ;
			RECT	10.883 75.924 10.915 75.988 ;
			RECT	11.051 75.924 11.083 75.988 ;
			RECT	11.219 75.924 11.251 75.988 ;
			RECT	11.387 75.924 11.419 75.988 ;
			RECT	11.555 75.924 11.587 75.988 ;
			RECT	11.723 75.924 11.755 75.988 ;
			RECT	11.891 75.924 11.923 75.988 ;
			RECT	12.059 75.924 12.091 75.988 ;
			RECT	12.227 75.924 12.259 75.988 ;
			RECT	12.395 75.924 12.427 75.988 ;
			RECT	12.563 75.924 12.595 75.988 ;
			RECT	12.731 75.924 12.763 75.988 ;
			RECT	12.899 75.924 12.931 75.988 ;
			RECT	13.067 75.924 13.099 75.988 ;
			RECT	13.235 75.924 13.267 75.988 ;
			RECT	13.403 75.924 13.435 75.988 ;
			RECT	13.571 75.924 13.603 75.988 ;
			RECT	13.739 75.924 13.771 75.988 ;
			RECT	13.907 75.924 13.939 75.988 ;
			RECT	14.075 75.924 14.107 75.988 ;
			RECT	14.243 75.924 14.275 75.988 ;
			RECT	14.411 75.924 14.443 75.988 ;
			RECT	14.579 75.924 14.611 75.988 ;
			RECT	14.747 75.924 14.779 75.988 ;
			RECT	14.915 75.924 14.947 75.988 ;
			RECT	15.083 75.924 15.115 75.988 ;
			RECT	15.251 75.924 15.283 75.988 ;
			RECT	15.419 75.924 15.451 75.988 ;
			RECT	15.587 75.924 15.619 75.988 ;
			RECT	15.755 75.924 15.787 75.988 ;
			RECT	15.923 75.924 15.955 75.988 ;
			RECT	16.091 75.924 16.123 75.988 ;
			RECT	16.259 75.924 16.291 75.988 ;
			RECT	16.427 75.924 16.459 75.988 ;
			RECT	16.595 75.924 16.627 75.988 ;
			RECT	16.763 75.924 16.795 75.988 ;
			RECT	16.931 75.924 16.963 75.988 ;
			RECT	17.099 75.924 17.131 75.988 ;
			RECT	17.267 75.924 17.299 75.988 ;
			RECT	17.435 75.924 17.467 75.988 ;
			RECT	17.603 75.924 17.635 75.988 ;
			RECT	17.771 75.924 17.803 75.988 ;
			RECT	17.939 75.924 17.971 75.988 ;
			RECT	18.107 75.924 18.139 75.988 ;
			RECT	18.275 75.924 18.307 75.988 ;
			RECT	18.443 75.924 18.475 75.988 ;
			RECT	18.611 75.924 18.643 75.988 ;
			RECT	18.779 75.924 18.811 75.988 ;
			RECT	18.947 75.924 18.979 75.988 ;
			RECT	19.115 75.924 19.147 75.988 ;
			RECT	19.283 75.924 19.315 75.988 ;
			RECT	19.451 75.924 19.483 75.988 ;
			RECT	19.619 75.924 19.651 75.988 ;
			RECT	19.787 75.924 19.819 75.988 ;
			RECT	19.955 75.924 19.987 75.988 ;
			RECT	20.123 75.924 20.155 75.988 ;
			RECT	20.291 75.924 20.323 75.988 ;
			RECT	20.459 75.924 20.491 75.988 ;
			RECT	20.627 75.924 20.659 75.988 ;
			RECT	20.795 75.924 20.827 75.988 ;
			RECT	20.963 75.924 20.995 75.988 ;
			RECT	21.131 75.924 21.163 75.988 ;
			RECT	21.299 75.924 21.331 75.988 ;
			RECT	21.467 75.924 21.499 75.988 ;
			RECT	21.635 75.924 21.667 75.988 ;
			RECT	21.803 75.924 21.835 75.988 ;
			RECT	21.971 75.924 22.003 75.988 ;
			RECT	22.139 75.924 22.171 75.988 ;
			RECT	22.307 75.924 22.339 75.988 ;
			RECT	22.475 75.924 22.507 75.988 ;
			RECT	22.643 75.924 22.675 75.988 ;
			RECT	22.811 75.924 22.843 75.988 ;
			RECT	22.979 75.924 23.011 75.988 ;
			RECT	23.147 75.924 23.179 75.988 ;
			RECT	23.315 75.924 23.347 75.988 ;
			RECT	23.483 75.924 23.515 75.988 ;
			RECT	23.651 75.924 23.683 75.988 ;
			RECT	23.819 75.924 23.851 75.988 ;
			RECT	23.987 75.924 24.019 75.988 ;
			RECT	24.155 75.924 24.187 75.988 ;
			RECT	24.323 75.924 24.355 75.988 ;
			RECT	24.491 75.924 24.523 75.988 ;
			RECT	24.659 75.924 24.691 75.988 ;
			RECT	24.827 75.924 24.859 75.988 ;
			RECT	24.995 75.924 25.027 75.988 ;
			RECT	25.163 75.924 25.195 75.988 ;
			RECT	25.331 75.924 25.363 75.988 ;
			RECT	25.499 75.924 25.531 75.988 ;
			RECT	25.667 75.924 25.699 75.988 ;
			RECT	25.835 75.924 25.867 75.988 ;
			RECT	26.003 75.924 26.035 75.988 ;
			RECT	26.171 75.924 26.203 75.988 ;
			RECT	26.339 75.924 26.371 75.988 ;
			RECT	26.507 75.924 26.539 75.988 ;
			RECT	26.675 75.924 26.707 75.988 ;
			RECT	26.843 75.924 26.875 75.988 ;
			RECT	27.011 75.924 27.043 75.988 ;
			RECT	27.179 75.924 27.211 75.988 ;
			RECT	27.347 75.924 27.379 75.988 ;
			RECT	27.515 75.924 27.547 75.988 ;
			RECT	27.683 75.924 27.715 75.988 ;
			RECT	27.851 75.924 27.883 75.988 ;
			RECT	28.019 75.924 28.051 75.988 ;
			RECT	28.187 75.924 28.219 75.988 ;
			RECT	28.355 75.924 28.387 75.988 ;
			RECT	28.523 75.924 28.555 75.988 ;
			RECT	28.691 75.924 28.723 75.988 ;
			RECT	28.859 75.924 28.891 75.988 ;
			RECT	29.027 75.924 29.059 75.988 ;
			RECT	29.195 75.924 29.227 75.988 ;
			RECT	29.363 75.924 29.395 75.988 ;
			RECT	29.531 75.924 29.563 75.988 ;
			RECT	29.699 75.924 29.731 75.988 ;
			RECT	29.867 75.924 29.899 75.988 ;
			RECT	30.035 75.924 30.067 75.988 ;
			RECT	30.203 75.924 30.235 75.988 ;
			RECT	30.371 75.924 30.403 75.988 ;
			RECT	30.539 75.924 30.571 75.988 ;
			RECT	30.707 75.924 30.739 75.988 ;
			RECT	30.875 75.924 30.907 75.988 ;
			RECT	31.043 75.924 31.075 75.988 ;
			RECT	31.211 75.924 31.243 75.988 ;
			RECT	31.379 75.924 31.411 75.988 ;
			RECT	31.547 75.924 31.579 75.988 ;
			RECT	31.715 75.924 31.747 75.988 ;
			RECT	31.883 75.924 31.915 75.988 ;
			RECT	32.051 75.924 32.083 75.988 ;
			RECT	32.219 75.924 32.251 75.988 ;
			RECT	32.387 75.924 32.419 75.988 ;
			RECT	32.555 75.924 32.587 75.988 ;
			RECT	32.723 75.924 32.755 75.988 ;
			RECT	32.891 75.924 32.923 75.988 ;
			RECT	33.059 75.924 33.091 75.988 ;
			RECT	33.227 75.924 33.259 75.988 ;
			RECT	33.395 75.924 33.427 75.988 ;
			RECT	33.563 75.924 33.595 75.988 ;
			RECT	33.731 75.924 33.763 75.988 ;
			RECT	33.899 75.924 33.931 75.988 ;
			RECT	34.067 75.924 34.099 75.988 ;
			RECT	34.235 75.924 34.267 75.988 ;
			RECT	34.403 75.924 34.435 75.988 ;
			RECT	34.571 75.924 34.603 75.988 ;
			RECT	34.739 75.924 34.771 75.988 ;
			RECT	34.907 75.924 34.939 75.988 ;
			RECT	35.075 75.924 35.107 75.988 ;
			RECT	35.243 75.924 35.275 75.988 ;
			RECT	35.411 75.924 35.443 75.988 ;
			RECT	35.579 75.924 35.611 75.988 ;
			RECT	35.747 75.924 35.779 75.988 ;
			RECT	35.915 75.924 35.947 75.988 ;
			RECT	36.083 75.924 36.115 75.988 ;
			RECT	36.251 75.924 36.283 75.988 ;
			RECT	36.419 75.924 36.451 75.988 ;
			RECT	36.587 75.924 36.619 75.988 ;
			RECT	36.755 75.924 36.787 75.988 ;
			RECT	36.923 75.924 36.955 75.988 ;
			RECT	37.091 75.924 37.123 75.988 ;
			RECT	37.259 75.924 37.291 75.988 ;
			RECT	37.427 75.924 37.459 75.988 ;
			RECT	37.595 75.924 37.627 75.988 ;
			RECT	37.763 75.924 37.795 75.988 ;
			RECT	37.931 75.924 37.963 75.988 ;
			RECT	38.099 75.924 38.131 75.988 ;
			RECT	38.267 75.924 38.299 75.988 ;
			RECT	38.435 75.924 38.467 75.988 ;
			RECT	38.603 75.924 38.635 75.988 ;
			RECT	38.771 75.924 38.803 75.988 ;
			RECT	38.939 75.924 38.971 75.988 ;
			RECT	39.107 75.924 39.139 75.988 ;
			RECT	39.275 75.924 39.307 75.988 ;
			RECT	39.443 75.924 39.475 75.988 ;
			RECT	39.611 75.924 39.643 75.988 ;
			RECT	39.779 75.924 39.811 75.988 ;
			RECT	39.947 75.924 39.979 75.988 ;
			RECT	40.115 75.924 40.147 75.988 ;
			RECT	40.283 75.924 40.315 75.988 ;
			RECT	40.451 75.924 40.483 75.988 ;
			RECT	40.619 75.924 40.651 75.988 ;
			RECT	40.787 75.924 40.819 75.988 ;
			RECT	40.955 75.924 40.987 75.988 ;
			RECT	41.123 75.924 41.155 75.988 ;
			RECT	41.291 75.924 41.323 75.988 ;
			RECT	41.459 75.924 41.491 75.988 ;
			RECT	41.627 75.924 41.659 75.988 ;
			RECT	41.795 75.924 41.827 75.988 ;
			RECT	41.963 75.924 41.995 75.988 ;
			RECT	42.131 75.924 42.163 75.988 ;
			RECT	42.299 75.924 42.331 75.988 ;
			RECT	42.467 75.924 42.499 75.988 ;
			RECT	42.635 75.924 42.667 75.988 ;
			RECT	42.803 75.924 42.835 75.988 ;
			RECT	42.971 75.924 43.003 75.988 ;
			RECT	43.139 75.924 43.171 75.988 ;
			RECT	43.307 75.924 43.339 75.988 ;
			RECT	43.475 75.924 43.507 75.988 ;
			RECT	43.643 75.924 43.675 75.988 ;
			RECT	43.811 75.924 43.843 75.988 ;
			RECT	43.979 75.924 44.011 75.988 ;
			RECT	44.147 75.924 44.179 75.988 ;
			RECT	44.315 75.924 44.347 75.988 ;
			RECT	44.483 75.924 44.515 75.988 ;
			RECT	44.651 75.924 44.683 75.988 ;
			RECT	44.819 75.924 44.851 75.988 ;
			RECT	44.987 75.924 45.019 75.988 ;
			RECT	45.155 75.924 45.187 75.988 ;
			RECT	45.323 75.924 45.355 75.988 ;
			RECT	45.491 75.924 45.523 75.988 ;
			RECT	45.659 75.924 45.691 75.988 ;
			RECT	45.827 75.924 45.859 75.988 ;
			RECT	45.995 75.924 46.027 75.988 ;
			RECT	46.163 75.924 46.195 75.988 ;
			RECT	46.331 75.924 46.363 75.988 ;
			RECT	46.499 75.924 46.531 75.988 ;
			RECT	46.667 75.924 46.699 75.988 ;
			RECT	46.835 75.924 46.867 75.988 ;
			RECT	47.003 75.924 47.035 75.988 ;
			RECT	47.171 75.924 47.203 75.988 ;
			RECT	47.339 75.924 47.371 75.988 ;
			RECT	47.507 75.924 47.539 75.988 ;
			RECT	47.675 75.924 47.707 75.988 ;
			RECT	47.843 75.924 47.875 75.988 ;
			RECT	48.011 75.924 48.043 75.988 ;
			RECT	48.179 75.924 48.211 75.988 ;
			RECT	48.347 75.924 48.379 75.988 ;
			RECT	48.515 75.924 48.547 75.988 ;
			RECT	48.683 75.924 48.715 75.988 ;
			RECT	48.851 75.924 48.883 75.988 ;
			RECT	49.019 75.924 49.051 75.988 ;
			RECT	49.187 75.924 49.219 75.988 ;
			RECT	49.318 75.94 49.35 75.972 ;
			RECT	49.439 75.94 49.471 75.972 ;
			RECT	49.569 75.924 49.601 75.988 ;
			RECT	51.881 75.924 51.913 75.988 ;
			RECT	53.132 75.924 53.196 75.988 ;
			RECT	53.812 75.924 53.844 75.988 ;
			RECT	54.251 75.924 54.283 75.988 ;
			RECT	55.562 75.924 55.626 75.988 ;
			RECT	58.603 75.924 58.635 75.988 ;
			RECT	58.733 75.94 58.765 75.972 ;
			RECT	58.854 75.94 58.886 75.972 ;
			RECT	58.985 75.924 59.017 75.988 ;
			RECT	59.153 75.924 59.185 75.988 ;
			RECT	59.321 75.924 59.353 75.988 ;
			RECT	59.489 75.924 59.521 75.988 ;
			RECT	59.657 75.924 59.689 75.988 ;
			RECT	59.825 75.924 59.857 75.988 ;
			RECT	59.993 75.924 60.025 75.988 ;
			RECT	60.161 75.924 60.193 75.988 ;
			RECT	60.329 75.924 60.361 75.988 ;
			RECT	60.497 75.924 60.529 75.988 ;
			RECT	60.665 75.924 60.697 75.988 ;
			RECT	60.833 75.924 60.865 75.988 ;
			RECT	61.001 75.924 61.033 75.988 ;
			RECT	61.169 75.924 61.201 75.988 ;
			RECT	61.337 75.924 61.369 75.988 ;
			RECT	61.505 75.924 61.537 75.988 ;
			RECT	61.673 75.924 61.705 75.988 ;
			RECT	61.841 75.924 61.873 75.988 ;
			RECT	62.009 75.924 62.041 75.988 ;
			RECT	62.177 75.924 62.209 75.988 ;
			RECT	62.345 75.924 62.377 75.988 ;
			RECT	62.513 75.924 62.545 75.988 ;
			RECT	62.681 75.924 62.713 75.988 ;
			RECT	62.849 75.924 62.881 75.988 ;
			RECT	63.017 75.924 63.049 75.988 ;
			RECT	63.185 75.924 63.217 75.988 ;
			RECT	63.353 75.924 63.385 75.988 ;
			RECT	63.521 75.924 63.553 75.988 ;
			RECT	63.689 75.924 63.721 75.988 ;
			RECT	63.857 75.924 63.889 75.988 ;
			RECT	64.025 75.924 64.057 75.988 ;
			RECT	64.193 75.924 64.225 75.988 ;
			RECT	64.361 75.924 64.393 75.988 ;
			RECT	64.529 75.924 64.561 75.988 ;
			RECT	64.697 75.924 64.729 75.988 ;
			RECT	64.865 75.924 64.897 75.988 ;
			RECT	65.033 75.924 65.065 75.988 ;
			RECT	65.201 75.924 65.233 75.988 ;
			RECT	65.369 75.924 65.401 75.988 ;
			RECT	65.537 75.924 65.569 75.988 ;
			RECT	65.705 75.924 65.737 75.988 ;
			RECT	65.873 75.924 65.905 75.988 ;
			RECT	66.041 75.924 66.073 75.988 ;
			RECT	66.209 75.924 66.241 75.988 ;
			RECT	66.377 75.924 66.409 75.988 ;
			RECT	66.545 75.924 66.577 75.988 ;
			RECT	66.713 75.924 66.745 75.988 ;
			RECT	66.881 75.924 66.913 75.988 ;
			RECT	67.049 75.924 67.081 75.988 ;
			RECT	67.217 75.924 67.249 75.988 ;
			RECT	67.385 75.924 67.417 75.988 ;
			RECT	67.553 75.924 67.585 75.988 ;
			RECT	67.721 75.924 67.753 75.988 ;
			RECT	67.889 75.924 67.921 75.988 ;
			RECT	68.057 75.924 68.089 75.988 ;
			RECT	68.225 75.924 68.257 75.988 ;
			RECT	68.393 75.924 68.425 75.988 ;
			RECT	68.561 75.924 68.593 75.988 ;
			RECT	68.729 75.924 68.761 75.988 ;
			RECT	68.897 75.924 68.929 75.988 ;
			RECT	69.065 75.924 69.097 75.988 ;
			RECT	69.233 75.924 69.265 75.988 ;
			RECT	69.401 75.924 69.433 75.988 ;
			RECT	69.569 75.924 69.601 75.988 ;
			RECT	69.737 75.924 69.769 75.988 ;
			RECT	69.905 75.924 69.937 75.988 ;
			RECT	70.073 75.924 70.105 75.988 ;
			RECT	70.241 75.924 70.273 75.988 ;
			RECT	70.409 75.924 70.441 75.988 ;
			RECT	70.577 75.924 70.609 75.988 ;
			RECT	70.745 75.924 70.777 75.988 ;
			RECT	70.913 75.924 70.945 75.988 ;
			RECT	71.081 75.924 71.113 75.988 ;
			RECT	71.249 75.924 71.281 75.988 ;
			RECT	71.417 75.924 71.449 75.988 ;
			RECT	71.585 75.924 71.617 75.988 ;
			RECT	71.753 75.924 71.785 75.988 ;
			RECT	71.921 75.924 71.953 75.988 ;
			RECT	72.089 75.924 72.121 75.988 ;
			RECT	72.257 75.924 72.289 75.988 ;
			RECT	72.425 75.924 72.457 75.988 ;
			RECT	72.593 75.924 72.625 75.988 ;
			RECT	72.761 75.924 72.793 75.988 ;
			RECT	72.929 75.924 72.961 75.988 ;
			RECT	73.097 75.924 73.129 75.988 ;
			RECT	73.265 75.924 73.297 75.988 ;
			RECT	73.433 75.924 73.465 75.988 ;
			RECT	73.601 75.924 73.633 75.988 ;
			RECT	73.769 75.924 73.801 75.988 ;
			RECT	73.937 75.924 73.969 75.988 ;
			RECT	74.105 75.924 74.137 75.988 ;
			RECT	74.273 75.924 74.305 75.988 ;
			RECT	74.441 75.924 74.473 75.988 ;
			RECT	74.609 75.924 74.641 75.988 ;
			RECT	74.777 75.924 74.809 75.988 ;
			RECT	74.945 75.924 74.977 75.988 ;
			RECT	75.113 75.924 75.145 75.988 ;
			RECT	75.281 75.924 75.313 75.988 ;
			RECT	75.449 75.924 75.481 75.988 ;
			RECT	75.617 75.924 75.649 75.988 ;
			RECT	75.785 75.924 75.817 75.988 ;
			RECT	75.953 75.924 75.985 75.988 ;
			RECT	76.121 75.924 76.153 75.988 ;
			RECT	76.289 75.924 76.321 75.988 ;
			RECT	76.457 75.924 76.489 75.988 ;
			RECT	76.625 75.924 76.657 75.988 ;
			RECT	76.793 75.924 76.825 75.988 ;
			RECT	76.961 75.924 76.993 75.988 ;
			RECT	77.129 75.924 77.161 75.988 ;
			RECT	77.297 75.924 77.329 75.988 ;
			RECT	77.465 75.924 77.497 75.988 ;
			RECT	77.633 75.924 77.665 75.988 ;
			RECT	77.801 75.924 77.833 75.988 ;
			RECT	77.969 75.924 78.001 75.988 ;
			RECT	78.137 75.924 78.169 75.988 ;
			RECT	78.305 75.924 78.337 75.988 ;
			RECT	78.473 75.924 78.505 75.988 ;
			RECT	78.641 75.924 78.673 75.988 ;
			RECT	78.809 75.924 78.841 75.988 ;
			RECT	78.977 75.924 79.009 75.988 ;
			RECT	79.145 75.924 79.177 75.988 ;
			RECT	79.313 75.924 79.345 75.988 ;
			RECT	79.481 75.924 79.513 75.988 ;
			RECT	79.649 75.924 79.681 75.988 ;
			RECT	79.817 75.924 79.849 75.988 ;
			RECT	79.985 75.924 80.017 75.988 ;
			RECT	80.153 75.924 80.185 75.988 ;
			RECT	80.321 75.924 80.353 75.988 ;
			RECT	80.489 75.924 80.521 75.988 ;
			RECT	80.657 75.924 80.689 75.988 ;
			RECT	80.825 75.924 80.857 75.988 ;
			RECT	80.993 75.924 81.025 75.988 ;
			RECT	81.161 75.924 81.193 75.988 ;
			RECT	81.329 75.924 81.361 75.988 ;
			RECT	81.497 75.924 81.529 75.988 ;
			RECT	81.665 75.924 81.697 75.988 ;
			RECT	81.833 75.924 81.865 75.988 ;
			RECT	82.001 75.924 82.033 75.988 ;
			RECT	82.169 75.924 82.201 75.988 ;
			RECT	82.337 75.924 82.369 75.988 ;
			RECT	82.505 75.924 82.537 75.988 ;
			RECT	82.673 75.924 82.705 75.988 ;
			RECT	82.841 75.924 82.873 75.988 ;
			RECT	83.009 75.924 83.041 75.988 ;
			RECT	83.177 75.924 83.209 75.988 ;
			RECT	83.345 75.924 83.377 75.988 ;
			RECT	83.513 75.924 83.545 75.988 ;
			RECT	83.681 75.924 83.713 75.988 ;
			RECT	83.849 75.924 83.881 75.988 ;
			RECT	84.017 75.924 84.049 75.988 ;
			RECT	84.185 75.924 84.217 75.988 ;
			RECT	84.353 75.924 84.385 75.988 ;
			RECT	84.521 75.924 84.553 75.988 ;
			RECT	84.689 75.924 84.721 75.988 ;
			RECT	84.857 75.924 84.889 75.988 ;
			RECT	85.025 75.924 85.057 75.988 ;
			RECT	85.193 75.924 85.225 75.988 ;
			RECT	85.361 75.924 85.393 75.988 ;
			RECT	85.529 75.924 85.561 75.988 ;
			RECT	85.697 75.924 85.729 75.988 ;
			RECT	85.865 75.924 85.897 75.988 ;
			RECT	86.033 75.924 86.065 75.988 ;
			RECT	86.201 75.924 86.233 75.988 ;
			RECT	86.369 75.924 86.401 75.988 ;
			RECT	86.537 75.924 86.569 75.988 ;
			RECT	86.705 75.924 86.737 75.988 ;
			RECT	86.873 75.924 86.905 75.988 ;
			RECT	87.041 75.924 87.073 75.988 ;
			RECT	87.209 75.924 87.241 75.988 ;
			RECT	87.377 75.924 87.409 75.988 ;
			RECT	87.545 75.924 87.577 75.988 ;
			RECT	87.713 75.924 87.745 75.988 ;
			RECT	87.881 75.924 87.913 75.988 ;
			RECT	88.049 75.924 88.081 75.988 ;
			RECT	88.217 75.924 88.249 75.988 ;
			RECT	88.385 75.924 88.417 75.988 ;
			RECT	88.553 75.924 88.585 75.988 ;
			RECT	88.721 75.924 88.753 75.988 ;
			RECT	88.889 75.924 88.921 75.988 ;
			RECT	89.057 75.924 89.089 75.988 ;
			RECT	89.225 75.924 89.257 75.988 ;
			RECT	89.393 75.924 89.425 75.988 ;
			RECT	89.561 75.924 89.593 75.988 ;
			RECT	89.729 75.924 89.761 75.988 ;
			RECT	89.897 75.924 89.929 75.988 ;
			RECT	90.065 75.924 90.097 75.988 ;
			RECT	90.233 75.924 90.265 75.988 ;
			RECT	90.401 75.924 90.433 75.988 ;
			RECT	90.569 75.924 90.601 75.988 ;
			RECT	90.737 75.924 90.769 75.988 ;
			RECT	90.905 75.924 90.937 75.988 ;
			RECT	91.073 75.924 91.105 75.988 ;
			RECT	91.241 75.924 91.273 75.988 ;
			RECT	91.409 75.924 91.441 75.988 ;
			RECT	91.577 75.924 91.609 75.988 ;
			RECT	91.745 75.924 91.777 75.988 ;
			RECT	91.913 75.924 91.945 75.988 ;
			RECT	92.081 75.924 92.113 75.988 ;
			RECT	92.249 75.924 92.281 75.988 ;
			RECT	92.417 75.924 92.449 75.988 ;
			RECT	92.585 75.924 92.617 75.988 ;
			RECT	92.753 75.924 92.785 75.988 ;
			RECT	92.921 75.924 92.953 75.988 ;
			RECT	93.089 75.924 93.121 75.988 ;
			RECT	93.257 75.924 93.289 75.988 ;
			RECT	93.425 75.924 93.457 75.988 ;
			RECT	93.593 75.924 93.625 75.988 ;
			RECT	93.761 75.924 93.793 75.988 ;
			RECT	93.929 75.924 93.961 75.988 ;
			RECT	94.097 75.924 94.129 75.988 ;
			RECT	94.265 75.924 94.297 75.988 ;
			RECT	94.433 75.924 94.465 75.988 ;
			RECT	94.601 75.924 94.633 75.988 ;
			RECT	94.769 75.924 94.801 75.988 ;
			RECT	94.937 75.924 94.969 75.988 ;
			RECT	95.105 75.924 95.137 75.988 ;
			RECT	95.273 75.924 95.305 75.988 ;
			RECT	95.441 75.924 95.473 75.988 ;
			RECT	95.609 75.924 95.641 75.988 ;
			RECT	95.777 75.924 95.809 75.988 ;
			RECT	95.945 75.924 95.977 75.988 ;
			RECT	96.113 75.924 96.145 75.988 ;
			RECT	96.281 75.924 96.313 75.988 ;
			RECT	96.449 75.924 96.481 75.988 ;
			RECT	96.617 75.924 96.649 75.988 ;
			RECT	96.785 75.924 96.817 75.988 ;
			RECT	96.953 75.924 96.985 75.988 ;
			RECT	97.121 75.924 97.153 75.988 ;
			RECT	97.289 75.924 97.321 75.988 ;
			RECT	97.457 75.924 97.489 75.988 ;
			RECT	97.625 75.924 97.657 75.988 ;
			RECT	97.793 75.924 97.825 75.988 ;
			RECT	97.961 75.924 97.993 75.988 ;
			RECT	98.129 75.924 98.161 75.988 ;
			RECT	98.297 75.924 98.329 75.988 ;
			RECT	98.465 75.924 98.497 75.988 ;
			RECT	98.633 75.924 98.665 75.988 ;
			RECT	98.801 75.924 98.833 75.988 ;
			RECT	98.969 75.924 99.001 75.988 ;
			RECT	99.137 75.924 99.169 75.988 ;
			RECT	99.305 75.924 99.337 75.988 ;
			RECT	99.473 75.924 99.505 75.988 ;
			RECT	99.641 75.924 99.673 75.988 ;
			RECT	99.809 75.924 99.841 75.988 ;
			RECT	99.977 75.924 100.009 75.988 ;
			RECT	100.145 75.924 100.177 75.988 ;
			RECT	100.313 75.924 100.345 75.988 ;
			RECT	100.481 75.924 100.513 75.988 ;
			RECT	100.649 75.924 100.681 75.988 ;
			RECT	100.817 75.924 100.849 75.988 ;
			RECT	100.985 75.924 101.017 75.988 ;
			RECT	101.153 75.924 101.185 75.988 ;
			RECT	101.321 75.924 101.353 75.988 ;
			RECT	101.489 75.924 101.521 75.988 ;
			RECT	101.657 75.924 101.689 75.988 ;
			RECT	101.825 75.924 101.857 75.988 ;
			RECT	101.993 75.924 102.025 75.988 ;
			RECT	102.123 75.94 102.155 75.972 ;
			RECT	102.245 75.935 102.277 75.967 ;
			RECT	102.375 75.924 102.407 75.988 ;
			RECT	103.795 75.924 103.827 75.988 ;
			RECT	103.925 75.935 103.957 75.967 ;
			RECT	104.047 75.94 104.079 75.972 ;
			RECT	104.177 75.924 104.209 75.988 ;
			RECT	104.345 75.924 104.377 75.988 ;
			RECT	104.513 75.924 104.545 75.988 ;
			RECT	104.681 75.924 104.713 75.988 ;
			RECT	104.849 75.924 104.881 75.988 ;
			RECT	105.017 75.924 105.049 75.988 ;
			RECT	105.185 75.924 105.217 75.988 ;
			RECT	105.353 75.924 105.385 75.988 ;
			RECT	105.521 75.924 105.553 75.988 ;
			RECT	105.689 75.924 105.721 75.988 ;
			RECT	105.857 75.924 105.889 75.988 ;
			RECT	106.025 75.924 106.057 75.988 ;
			RECT	106.193 75.924 106.225 75.988 ;
			RECT	106.361 75.924 106.393 75.988 ;
			RECT	106.529 75.924 106.561 75.988 ;
			RECT	106.697 75.924 106.729 75.988 ;
			RECT	106.865 75.924 106.897 75.988 ;
			RECT	107.033 75.924 107.065 75.988 ;
			RECT	107.201 75.924 107.233 75.988 ;
			RECT	107.369 75.924 107.401 75.988 ;
			RECT	107.537 75.924 107.569 75.988 ;
			RECT	107.705 75.924 107.737 75.988 ;
			RECT	107.873 75.924 107.905 75.988 ;
			RECT	108.041 75.924 108.073 75.988 ;
			RECT	108.209 75.924 108.241 75.988 ;
			RECT	108.377 75.924 108.409 75.988 ;
			RECT	108.545 75.924 108.577 75.988 ;
			RECT	108.713 75.924 108.745 75.988 ;
			RECT	108.881 75.924 108.913 75.988 ;
			RECT	109.049 75.924 109.081 75.988 ;
			RECT	109.217 75.924 109.249 75.988 ;
			RECT	109.385 75.924 109.417 75.988 ;
			RECT	109.553 75.924 109.585 75.988 ;
			RECT	109.721 75.924 109.753 75.988 ;
			RECT	109.889 75.924 109.921 75.988 ;
			RECT	110.057 75.924 110.089 75.988 ;
			RECT	110.225 75.924 110.257 75.988 ;
			RECT	110.393 75.924 110.425 75.988 ;
			RECT	110.561 75.924 110.593 75.988 ;
			RECT	110.729 75.924 110.761 75.988 ;
			RECT	110.897 75.924 110.929 75.988 ;
			RECT	111.065 75.924 111.097 75.988 ;
			RECT	111.233 75.924 111.265 75.988 ;
			RECT	111.401 75.924 111.433 75.988 ;
			RECT	111.569 75.924 111.601 75.988 ;
			RECT	111.737 75.924 111.769 75.988 ;
			RECT	111.905 75.924 111.937 75.988 ;
			RECT	112.073 75.924 112.105 75.988 ;
			RECT	112.241 75.924 112.273 75.988 ;
			RECT	112.409 75.924 112.441 75.988 ;
			RECT	112.577 75.924 112.609 75.988 ;
			RECT	112.745 75.924 112.777 75.988 ;
			RECT	112.913 75.924 112.945 75.988 ;
			RECT	113.081 75.924 113.113 75.988 ;
			RECT	113.249 75.924 113.281 75.988 ;
			RECT	113.417 75.924 113.449 75.988 ;
			RECT	113.585 75.924 113.617 75.988 ;
			RECT	113.753 75.924 113.785 75.988 ;
			RECT	113.921 75.924 113.953 75.988 ;
			RECT	114.089 75.924 114.121 75.988 ;
			RECT	114.257 75.924 114.289 75.988 ;
			RECT	114.425 75.924 114.457 75.988 ;
			RECT	114.593 75.924 114.625 75.988 ;
			RECT	114.761 75.924 114.793 75.988 ;
			RECT	114.929 75.924 114.961 75.988 ;
			RECT	115.097 75.924 115.129 75.988 ;
			RECT	115.265 75.924 115.297 75.988 ;
			RECT	115.433 75.924 115.465 75.988 ;
			RECT	115.601 75.924 115.633 75.988 ;
			RECT	115.769 75.924 115.801 75.988 ;
			RECT	115.937 75.924 115.969 75.988 ;
			RECT	116.105 75.924 116.137 75.988 ;
			RECT	116.273 75.924 116.305 75.988 ;
			RECT	116.441 75.924 116.473 75.988 ;
			RECT	116.609 75.924 116.641 75.988 ;
			RECT	116.777 75.924 116.809 75.988 ;
			RECT	116.945 75.924 116.977 75.988 ;
			RECT	117.113 75.924 117.145 75.988 ;
			RECT	117.281 75.924 117.313 75.988 ;
			RECT	117.449 75.924 117.481 75.988 ;
			RECT	117.617 75.924 117.649 75.988 ;
			RECT	117.785 75.924 117.817 75.988 ;
			RECT	117.953 75.924 117.985 75.988 ;
			RECT	118.121 75.924 118.153 75.988 ;
			RECT	118.289 75.924 118.321 75.988 ;
			RECT	118.457 75.924 118.489 75.988 ;
			RECT	118.625 75.924 118.657 75.988 ;
			RECT	118.793 75.924 118.825 75.988 ;
			RECT	118.961 75.924 118.993 75.988 ;
			RECT	119.129 75.924 119.161 75.988 ;
			RECT	119.297 75.924 119.329 75.988 ;
			RECT	119.465 75.924 119.497 75.988 ;
			RECT	119.633 75.924 119.665 75.988 ;
			RECT	119.801 75.924 119.833 75.988 ;
			RECT	119.969 75.924 120.001 75.988 ;
			RECT	120.137 75.924 120.169 75.988 ;
			RECT	120.305 75.924 120.337 75.988 ;
			RECT	120.473 75.924 120.505 75.988 ;
			RECT	120.641 75.924 120.673 75.988 ;
			RECT	120.809 75.924 120.841 75.988 ;
			RECT	120.977 75.924 121.009 75.988 ;
			RECT	121.145 75.924 121.177 75.988 ;
			RECT	121.313 75.924 121.345 75.988 ;
			RECT	121.481 75.924 121.513 75.988 ;
			RECT	121.649 75.924 121.681 75.988 ;
			RECT	121.817 75.924 121.849 75.988 ;
			RECT	121.985 75.924 122.017 75.988 ;
			RECT	122.153 75.924 122.185 75.988 ;
			RECT	122.321 75.924 122.353 75.988 ;
			RECT	122.489 75.924 122.521 75.988 ;
			RECT	122.657 75.924 122.689 75.988 ;
			RECT	122.825 75.924 122.857 75.988 ;
			RECT	122.993 75.924 123.025 75.988 ;
			RECT	123.161 75.924 123.193 75.988 ;
			RECT	123.329 75.924 123.361 75.988 ;
			RECT	123.497 75.924 123.529 75.988 ;
			RECT	123.665 75.924 123.697 75.988 ;
			RECT	123.833 75.924 123.865 75.988 ;
			RECT	124.001 75.924 124.033 75.988 ;
			RECT	124.169 75.924 124.201 75.988 ;
			RECT	124.337 75.924 124.369 75.988 ;
			RECT	124.505 75.924 124.537 75.988 ;
			RECT	124.673 75.924 124.705 75.988 ;
			RECT	124.841 75.924 124.873 75.988 ;
			RECT	125.009 75.924 125.041 75.988 ;
			RECT	125.177 75.924 125.209 75.988 ;
			RECT	125.345 75.924 125.377 75.988 ;
			RECT	125.513 75.924 125.545 75.988 ;
			RECT	125.681 75.924 125.713 75.988 ;
			RECT	125.849 75.924 125.881 75.988 ;
			RECT	126.017 75.924 126.049 75.988 ;
			RECT	126.185 75.924 126.217 75.988 ;
			RECT	126.353 75.924 126.385 75.988 ;
			RECT	126.521 75.924 126.553 75.988 ;
			RECT	126.689 75.924 126.721 75.988 ;
			RECT	126.857 75.924 126.889 75.988 ;
			RECT	127.025 75.924 127.057 75.988 ;
			RECT	127.193 75.924 127.225 75.988 ;
			RECT	127.361 75.924 127.393 75.988 ;
			RECT	127.529 75.924 127.561 75.988 ;
			RECT	127.697 75.924 127.729 75.988 ;
			RECT	127.865 75.924 127.897 75.988 ;
			RECT	128.033 75.924 128.065 75.988 ;
			RECT	128.201 75.924 128.233 75.988 ;
			RECT	128.369 75.924 128.401 75.988 ;
			RECT	128.537 75.924 128.569 75.988 ;
			RECT	128.705 75.924 128.737 75.988 ;
			RECT	128.873 75.924 128.905 75.988 ;
			RECT	129.041 75.924 129.073 75.988 ;
			RECT	129.209 75.924 129.241 75.988 ;
			RECT	129.377 75.924 129.409 75.988 ;
			RECT	129.545 75.924 129.577 75.988 ;
			RECT	129.713 75.924 129.745 75.988 ;
			RECT	129.881 75.924 129.913 75.988 ;
			RECT	130.049 75.924 130.081 75.988 ;
			RECT	130.217 75.924 130.249 75.988 ;
			RECT	130.385 75.924 130.417 75.988 ;
			RECT	130.553 75.924 130.585 75.988 ;
			RECT	130.721 75.924 130.753 75.988 ;
			RECT	130.889 75.924 130.921 75.988 ;
			RECT	131.057 75.924 131.089 75.988 ;
			RECT	131.225 75.924 131.257 75.988 ;
			RECT	131.393 75.924 131.425 75.988 ;
			RECT	131.561 75.924 131.593 75.988 ;
			RECT	131.729 75.924 131.761 75.988 ;
			RECT	131.897 75.924 131.929 75.988 ;
			RECT	132.065 75.924 132.097 75.988 ;
			RECT	132.233 75.924 132.265 75.988 ;
			RECT	132.401 75.924 132.433 75.988 ;
			RECT	132.569 75.924 132.601 75.988 ;
			RECT	132.737 75.924 132.769 75.988 ;
			RECT	132.905 75.924 132.937 75.988 ;
			RECT	133.073 75.924 133.105 75.988 ;
			RECT	133.241 75.924 133.273 75.988 ;
			RECT	133.409 75.924 133.441 75.988 ;
			RECT	133.577 75.924 133.609 75.988 ;
			RECT	133.745 75.924 133.777 75.988 ;
			RECT	133.913 75.924 133.945 75.988 ;
			RECT	134.081 75.924 134.113 75.988 ;
			RECT	134.249 75.924 134.281 75.988 ;
			RECT	134.417 75.924 134.449 75.988 ;
			RECT	134.585 75.924 134.617 75.988 ;
			RECT	134.753 75.924 134.785 75.988 ;
			RECT	134.921 75.924 134.953 75.988 ;
			RECT	135.089 75.924 135.121 75.988 ;
			RECT	135.257 75.924 135.289 75.988 ;
			RECT	135.425 75.924 135.457 75.988 ;
			RECT	135.593 75.924 135.625 75.988 ;
			RECT	135.761 75.924 135.793 75.988 ;
			RECT	135.929 75.924 135.961 75.988 ;
			RECT	136.097 75.924 136.129 75.988 ;
			RECT	136.265 75.924 136.297 75.988 ;
			RECT	136.433 75.924 136.465 75.988 ;
			RECT	136.601 75.924 136.633 75.988 ;
			RECT	136.769 75.924 136.801 75.988 ;
			RECT	136.937 75.924 136.969 75.988 ;
			RECT	137.105 75.924 137.137 75.988 ;
			RECT	137.273 75.924 137.305 75.988 ;
			RECT	137.441 75.924 137.473 75.988 ;
			RECT	137.609 75.924 137.641 75.988 ;
			RECT	137.777 75.924 137.809 75.988 ;
			RECT	137.945 75.924 137.977 75.988 ;
			RECT	138.113 75.924 138.145 75.988 ;
			RECT	138.281 75.924 138.313 75.988 ;
			RECT	138.449 75.924 138.481 75.988 ;
			RECT	138.617 75.924 138.649 75.988 ;
			RECT	138.785 75.924 138.817 75.988 ;
			RECT	138.953 75.924 138.985 75.988 ;
			RECT	139.121 75.924 139.153 75.988 ;
			RECT	139.289 75.924 139.321 75.988 ;
			RECT	139.457 75.924 139.489 75.988 ;
			RECT	139.625 75.924 139.657 75.988 ;
			RECT	139.793 75.924 139.825 75.988 ;
			RECT	139.961 75.924 139.993 75.988 ;
			RECT	140.129 75.924 140.161 75.988 ;
			RECT	140.297 75.924 140.329 75.988 ;
			RECT	140.465 75.924 140.497 75.988 ;
			RECT	140.633 75.924 140.665 75.988 ;
			RECT	140.801 75.924 140.833 75.988 ;
			RECT	140.969 75.924 141.001 75.988 ;
			RECT	141.137 75.924 141.169 75.988 ;
			RECT	141.305 75.924 141.337 75.988 ;
			RECT	141.473 75.924 141.505 75.988 ;
			RECT	141.641 75.924 141.673 75.988 ;
			RECT	141.809 75.924 141.841 75.988 ;
			RECT	141.977 75.924 142.009 75.988 ;
			RECT	142.145 75.924 142.177 75.988 ;
			RECT	142.313 75.924 142.345 75.988 ;
			RECT	142.481 75.924 142.513 75.988 ;
			RECT	142.649 75.924 142.681 75.988 ;
			RECT	142.817 75.924 142.849 75.988 ;
			RECT	142.985 75.924 143.017 75.988 ;
			RECT	143.153 75.924 143.185 75.988 ;
			RECT	143.321 75.924 143.353 75.988 ;
			RECT	143.489 75.924 143.521 75.988 ;
			RECT	143.657 75.924 143.689 75.988 ;
			RECT	143.825 75.924 143.857 75.988 ;
			RECT	143.993 75.924 144.025 75.988 ;
			RECT	144.161 75.924 144.193 75.988 ;
			RECT	144.329 75.924 144.361 75.988 ;
			RECT	144.497 75.924 144.529 75.988 ;
			RECT	144.665 75.924 144.697 75.988 ;
			RECT	144.833 75.924 144.865 75.988 ;
			RECT	145.001 75.924 145.033 75.988 ;
			RECT	145.169 75.924 145.201 75.988 ;
			RECT	145.337 75.924 145.369 75.988 ;
			RECT	145.505 75.924 145.537 75.988 ;
			RECT	145.673 75.924 145.705 75.988 ;
			RECT	145.841 75.924 145.873 75.988 ;
			RECT	146.009 75.924 146.041 75.988 ;
			RECT	146.177 75.924 146.209 75.988 ;
			RECT	146.345 75.924 146.377 75.988 ;
			RECT	146.513 75.924 146.545 75.988 ;
			RECT	146.681 75.924 146.713 75.988 ;
			RECT	146.849 75.924 146.881 75.988 ;
			RECT	147.017 75.924 147.049 75.988 ;
			RECT	147.185 75.924 147.217 75.988 ;
			RECT	147.316 75.94 147.348 75.972 ;
			RECT	147.437 75.94 147.469 75.972 ;
			RECT	147.567 75.924 147.599 75.988 ;
			RECT	149.879 75.924 149.911 75.988 ;
			RECT	151.13 75.924 151.194 75.988 ;
			RECT	151.81 75.924 151.842 75.988 ;
			RECT	152.249 75.924 152.281 75.988 ;
			RECT	153.56 75.924 153.624 75.988 ;
			RECT	156.601 75.924 156.633 75.988 ;
			RECT	156.731 75.94 156.763 75.972 ;
			RECT	156.852 75.94 156.884 75.972 ;
			RECT	156.983 75.924 157.015 75.988 ;
			RECT	157.151 75.924 157.183 75.988 ;
			RECT	157.319 75.924 157.351 75.988 ;
			RECT	157.487 75.924 157.519 75.988 ;
			RECT	157.655 75.924 157.687 75.988 ;
			RECT	157.823 75.924 157.855 75.988 ;
			RECT	157.991 75.924 158.023 75.988 ;
			RECT	158.159 75.924 158.191 75.988 ;
			RECT	158.327 75.924 158.359 75.988 ;
			RECT	158.495 75.924 158.527 75.988 ;
			RECT	158.663 75.924 158.695 75.988 ;
			RECT	158.831 75.924 158.863 75.988 ;
			RECT	158.999 75.924 159.031 75.988 ;
			RECT	159.167 75.924 159.199 75.988 ;
			RECT	159.335 75.924 159.367 75.988 ;
			RECT	159.503 75.924 159.535 75.988 ;
			RECT	159.671 75.924 159.703 75.988 ;
			RECT	159.839 75.924 159.871 75.988 ;
			RECT	160.007 75.924 160.039 75.988 ;
			RECT	160.175 75.924 160.207 75.988 ;
			RECT	160.343 75.924 160.375 75.988 ;
			RECT	160.511 75.924 160.543 75.988 ;
			RECT	160.679 75.924 160.711 75.988 ;
			RECT	160.847 75.924 160.879 75.988 ;
			RECT	161.015 75.924 161.047 75.988 ;
			RECT	161.183 75.924 161.215 75.988 ;
			RECT	161.351 75.924 161.383 75.988 ;
			RECT	161.519 75.924 161.551 75.988 ;
			RECT	161.687 75.924 161.719 75.988 ;
			RECT	161.855 75.924 161.887 75.988 ;
			RECT	162.023 75.924 162.055 75.988 ;
			RECT	162.191 75.924 162.223 75.988 ;
			RECT	162.359 75.924 162.391 75.988 ;
			RECT	162.527 75.924 162.559 75.988 ;
			RECT	162.695 75.924 162.727 75.988 ;
			RECT	162.863 75.924 162.895 75.988 ;
			RECT	163.031 75.924 163.063 75.988 ;
			RECT	163.199 75.924 163.231 75.988 ;
			RECT	163.367 75.924 163.399 75.988 ;
			RECT	163.535 75.924 163.567 75.988 ;
			RECT	163.703 75.924 163.735 75.988 ;
			RECT	163.871 75.924 163.903 75.988 ;
			RECT	164.039 75.924 164.071 75.988 ;
			RECT	164.207 75.924 164.239 75.988 ;
			RECT	164.375 75.924 164.407 75.988 ;
			RECT	164.543 75.924 164.575 75.988 ;
			RECT	164.711 75.924 164.743 75.988 ;
			RECT	164.879 75.924 164.911 75.988 ;
			RECT	165.047 75.924 165.079 75.988 ;
			RECT	165.215 75.924 165.247 75.988 ;
			RECT	165.383 75.924 165.415 75.988 ;
			RECT	165.551 75.924 165.583 75.988 ;
			RECT	165.719 75.924 165.751 75.988 ;
			RECT	165.887 75.924 165.919 75.988 ;
			RECT	166.055 75.924 166.087 75.988 ;
			RECT	166.223 75.924 166.255 75.988 ;
			RECT	166.391 75.924 166.423 75.988 ;
			RECT	166.559 75.924 166.591 75.988 ;
			RECT	166.727 75.924 166.759 75.988 ;
			RECT	166.895 75.924 166.927 75.988 ;
			RECT	167.063 75.924 167.095 75.988 ;
			RECT	167.231 75.924 167.263 75.988 ;
			RECT	167.399 75.924 167.431 75.988 ;
			RECT	167.567 75.924 167.599 75.988 ;
			RECT	167.735 75.924 167.767 75.988 ;
			RECT	167.903 75.924 167.935 75.988 ;
			RECT	168.071 75.924 168.103 75.988 ;
			RECT	168.239 75.924 168.271 75.988 ;
			RECT	168.407 75.924 168.439 75.988 ;
			RECT	168.575 75.924 168.607 75.988 ;
			RECT	168.743 75.924 168.775 75.988 ;
			RECT	168.911 75.924 168.943 75.988 ;
			RECT	169.079 75.924 169.111 75.988 ;
			RECT	169.247 75.924 169.279 75.988 ;
			RECT	169.415 75.924 169.447 75.988 ;
			RECT	169.583 75.924 169.615 75.988 ;
			RECT	169.751 75.924 169.783 75.988 ;
			RECT	169.919 75.924 169.951 75.988 ;
			RECT	170.087 75.924 170.119 75.988 ;
			RECT	170.255 75.924 170.287 75.988 ;
			RECT	170.423 75.924 170.455 75.988 ;
			RECT	170.591 75.924 170.623 75.988 ;
			RECT	170.759 75.924 170.791 75.988 ;
			RECT	170.927 75.924 170.959 75.988 ;
			RECT	171.095 75.924 171.127 75.988 ;
			RECT	171.263 75.924 171.295 75.988 ;
			RECT	171.431 75.924 171.463 75.988 ;
			RECT	171.599 75.924 171.631 75.988 ;
			RECT	171.767 75.924 171.799 75.988 ;
			RECT	171.935 75.924 171.967 75.988 ;
			RECT	172.103 75.924 172.135 75.988 ;
			RECT	172.271 75.924 172.303 75.988 ;
			RECT	172.439 75.924 172.471 75.988 ;
			RECT	172.607 75.924 172.639 75.988 ;
			RECT	172.775 75.924 172.807 75.988 ;
			RECT	172.943 75.924 172.975 75.988 ;
			RECT	173.111 75.924 173.143 75.988 ;
			RECT	173.279 75.924 173.311 75.988 ;
			RECT	173.447 75.924 173.479 75.988 ;
			RECT	173.615 75.924 173.647 75.988 ;
			RECT	173.783 75.924 173.815 75.988 ;
			RECT	173.951 75.924 173.983 75.988 ;
			RECT	174.119 75.924 174.151 75.988 ;
			RECT	174.287 75.924 174.319 75.988 ;
			RECT	174.455 75.924 174.487 75.988 ;
			RECT	174.623 75.924 174.655 75.988 ;
			RECT	174.791 75.924 174.823 75.988 ;
			RECT	174.959 75.924 174.991 75.988 ;
			RECT	175.127 75.924 175.159 75.988 ;
			RECT	175.295 75.924 175.327 75.988 ;
			RECT	175.463 75.924 175.495 75.988 ;
			RECT	175.631 75.924 175.663 75.988 ;
			RECT	175.799 75.924 175.831 75.988 ;
			RECT	175.967 75.924 175.999 75.988 ;
			RECT	176.135 75.924 176.167 75.988 ;
			RECT	176.303 75.924 176.335 75.988 ;
			RECT	176.471 75.924 176.503 75.988 ;
			RECT	176.639 75.924 176.671 75.988 ;
			RECT	176.807 75.924 176.839 75.988 ;
			RECT	176.975 75.924 177.007 75.988 ;
			RECT	177.143 75.924 177.175 75.988 ;
			RECT	177.311 75.924 177.343 75.988 ;
			RECT	177.479 75.924 177.511 75.988 ;
			RECT	177.647 75.924 177.679 75.988 ;
			RECT	177.815 75.924 177.847 75.988 ;
			RECT	177.983 75.924 178.015 75.988 ;
			RECT	178.151 75.924 178.183 75.988 ;
			RECT	178.319 75.924 178.351 75.988 ;
			RECT	178.487 75.924 178.519 75.988 ;
			RECT	178.655 75.924 178.687 75.988 ;
			RECT	178.823 75.924 178.855 75.988 ;
			RECT	178.991 75.924 179.023 75.988 ;
			RECT	179.159 75.924 179.191 75.988 ;
			RECT	179.327 75.924 179.359 75.988 ;
			RECT	179.495 75.924 179.527 75.988 ;
			RECT	179.663 75.924 179.695 75.988 ;
			RECT	179.831 75.924 179.863 75.988 ;
			RECT	179.999 75.924 180.031 75.988 ;
			RECT	180.167 75.924 180.199 75.988 ;
			RECT	180.335 75.924 180.367 75.988 ;
			RECT	180.503 75.924 180.535 75.988 ;
			RECT	180.671 75.924 180.703 75.988 ;
			RECT	180.839 75.924 180.871 75.988 ;
			RECT	181.007 75.924 181.039 75.988 ;
			RECT	181.175 75.924 181.207 75.988 ;
			RECT	181.343 75.924 181.375 75.988 ;
			RECT	181.511 75.924 181.543 75.988 ;
			RECT	181.679 75.924 181.711 75.988 ;
			RECT	181.847 75.924 181.879 75.988 ;
			RECT	182.015 75.924 182.047 75.988 ;
			RECT	182.183 75.924 182.215 75.988 ;
			RECT	182.351 75.924 182.383 75.988 ;
			RECT	182.519 75.924 182.551 75.988 ;
			RECT	182.687 75.924 182.719 75.988 ;
			RECT	182.855 75.924 182.887 75.988 ;
			RECT	183.023 75.924 183.055 75.988 ;
			RECT	183.191 75.924 183.223 75.988 ;
			RECT	183.359 75.924 183.391 75.988 ;
			RECT	183.527 75.924 183.559 75.988 ;
			RECT	183.695 75.924 183.727 75.988 ;
			RECT	183.863 75.924 183.895 75.988 ;
			RECT	184.031 75.924 184.063 75.988 ;
			RECT	184.199 75.924 184.231 75.988 ;
			RECT	184.367 75.924 184.399 75.988 ;
			RECT	184.535 75.924 184.567 75.988 ;
			RECT	184.703 75.924 184.735 75.988 ;
			RECT	184.871 75.924 184.903 75.988 ;
			RECT	185.039 75.924 185.071 75.988 ;
			RECT	185.207 75.924 185.239 75.988 ;
			RECT	185.375 75.924 185.407 75.988 ;
			RECT	185.543 75.924 185.575 75.988 ;
			RECT	185.711 75.924 185.743 75.988 ;
			RECT	185.879 75.924 185.911 75.988 ;
			RECT	186.047 75.924 186.079 75.988 ;
			RECT	186.215 75.924 186.247 75.988 ;
			RECT	186.383 75.924 186.415 75.988 ;
			RECT	186.551 75.924 186.583 75.988 ;
			RECT	186.719 75.924 186.751 75.988 ;
			RECT	186.887 75.924 186.919 75.988 ;
			RECT	187.055 75.924 187.087 75.988 ;
			RECT	187.223 75.924 187.255 75.988 ;
			RECT	187.391 75.924 187.423 75.988 ;
			RECT	187.559 75.924 187.591 75.988 ;
			RECT	187.727 75.924 187.759 75.988 ;
			RECT	187.895 75.924 187.927 75.988 ;
			RECT	188.063 75.924 188.095 75.988 ;
			RECT	188.231 75.924 188.263 75.988 ;
			RECT	188.399 75.924 188.431 75.988 ;
			RECT	188.567 75.924 188.599 75.988 ;
			RECT	188.735 75.924 188.767 75.988 ;
			RECT	188.903 75.924 188.935 75.988 ;
			RECT	189.071 75.924 189.103 75.988 ;
			RECT	189.239 75.924 189.271 75.988 ;
			RECT	189.407 75.924 189.439 75.988 ;
			RECT	189.575 75.924 189.607 75.988 ;
			RECT	189.743 75.924 189.775 75.988 ;
			RECT	189.911 75.924 189.943 75.988 ;
			RECT	190.079 75.924 190.111 75.988 ;
			RECT	190.247 75.924 190.279 75.988 ;
			RECT	190.415 75.924 190.447 75.988 ;
			RECT	190.583 75.924 190.615 75.988 ;
			RECT	190.751 75.924 190.783 75.988 ;
			RECT	190.919 75.924 190.951 75.988 ;
			RECT	191.087 75.924 191.119 75.988 ;
			RECT	191.255 75.924 191.287 75.988 ;
			RECT	191.423 75.924 191.455 75.988 ;
			RECT	191.591 75.924 191.623 75.988 ;
			RECT	191.759 75.924 191.791 75.988 ;
			RECT	191.927 75.924 191.959 75.988 ;
			RECT	192.095 75.924 192.127 75.988 ;
			RECT	192.263 75.924 192.295 75.988 ;
			RECT	192.431 75.924 192.463 75.988 ;
			RECT	192.599 75.924 192.631 75.988 ;
			RECT	192.767 75.924 192.799 75.988 ;
			RECT	192.935 75.924 192.967 75.988 ;
			RECT	193.103 75.924 193.135 75.988 ;
			RECT	193.271 75.924 193.303 75.988 ;
			RECT	193.439 75.924 193.471 75.988 ;
			RECT	193.607 75.924 193.639 75.988 ;
			RECT	193.775 75.924 193.807 75.988 ;
			RECT	193.943 75.924 193.975 75.988 ;
			RECT	194.111 75.924 194.143 75.988 ;
			RECT	194.279 75.924 194.311 75.988 ;
			RECT	194.447 75.924 194.479 75.988 ;
			RECT	194.615 75.924 194.647 75.988 ;
			RECT	194.783 75.924 194.815 75.988 ;
			RECT	194.951 75.924 194.983 75.988 ;
			RECT	195.119 75.924 195.151 75.988 ;
			RECT	195.287 75.924 195.319 75.988 ;
			RECT	195.455 75.924 195.487 75.988 ;
			RECT	195.623 75.924 195.655 75.988 ;
			RECT	195.791 75.924 195.823 75.988 ;
			RECT	195.959 75.924 195.991 75.988 ;
			RECT	196.127 75.924 196.159 75.988 ;
			RECT	196.295 75.924 196.327 75.988 ;
			RECT	196.463 75.924 196.495 75.988 ;
			RECT	196.631 75.924 196.663 75.988 ;
			RECT	196.799 75.924 196.831 75.988 ;
			RECT	196.967 75.924 196.999 75.988 ;
			RECT	197.135 75.924 197.167 75.988 ;
			RECT	197.303 75.924 197.335 75.988 ;
			RECT	197.471 75.924 197.503 75.988 ;
			RECT	197.639 75.924 197.671 75.988 ;
			RECT	197.807 75.924 197.839 75.988 ;
			RECT	197.975 75.924 198.007 75.988 ;
			RECT	198.143 75.924 198.175 75.988 ;
			RECT	198.311 75.924 198.343 75.988 ;
			RECT	198.479 75.924 198.511 75.988 ;
			RECT	198.647 75.924 198.679 75.988 ;
			RECT	198.815 75.924 198.847 75.988 ;
			RECT	198.983 75.924 199.015 75.988 ;
			RECT	199.151 75.924 199.183 75.988 ;
			RECT	199.319 75.924 199.351 75.988 ;
			RECT	199.487 75.924 199.519 75.988 ;
			RECT	199.655 75.924 199.687 75.988 ;
			RECT	199.823 75.924 199.855 75.988 ;
			RECT	199.991 75.924 200.023 75.988 ;
			RECT	200.121 75.94 200.153 75.972 ;
			RECT	200.243 75.935 200.275 75.967 ;
			RECT	200.373 75.924 200.405 75.988 ;
			RECT	200.9 75.924 200.932 75.988 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 27.28 201.665 27.4 ;
			LAYER	J3 ;
			RECT	0.755 27.308 0.787 27.372 ;
			RECT	1.645 27.308 1.709 27.372 ;
			RECT	2.323 27.308 2.387 27.372 ;
			RECT	3.438 27.308 3.47 27.372 ;
			RECT	3.585 27.308 3.617 27.372 ;
			RECT	4.195 27.308 4.227 27.372 ;
			RECT	4.72 27.308 4.752 27.372 ;
			RECT	4.944 27.308 5.008 27.372 ;
			RECT	5.267 27.308 5.299 27.372 ;
			RECT	5.797 27.308 5.829 27.372 ;
			RECT	5.927 27.329 5.959 27.361 ;
			RECT	6.049 27.324 6.081 27.356 ;
			RECT	6.179 27.308 6.211 27.372 ;
			RECT	6.347 27.308 6.379 27.372 ;
			RECT	6.515 27.308 6.547 27.372 ;
			RECT	6.683 27.308 6.715 27.372 ;
			RECT	6.851 27.308 6.883 27.372 ;
			RECT	7.019 27.308 7.051 27.372 ;
			RECT	7.187 27.308 7.219 27.372 ;
			RECT	7.355 27.308 7.387 27.372 ;
			RECT	7.523 27.308 7.555 27.372 ;
			RECT	7.691 27.308 7.723 27.372 ;
			RECT	7.859 27.308 7.891 27.372 ;
			RECT	8.027 27.308 8.059 27.372 ;
			RECT	8.195 27.308 8.227 27.372 ;
			RECT	8.363 27.308 8.395 27.372 ;
			RECT	8.531 27.308 8.563 27.372 ;
			RECT	8.699 27.308 8.731 27.372 ;
			RECT	8.867 27.308 8.899 27.372 ;
			RECT	9.035 27.308 9.067 27.372 ;
			RECT	9.203 27.308 9.235 27.372 ;
			RECT	9.371 27.308 9.403 27.372 ;
			RECT	9.539 27.308 9.571 27.372 ;
			RECT	9.707 27.308 9.739 27.372 ;
			RECT	9.875 27.308 9.907 27.372 ;
			RECT	10.043 27.308 10.075 27.372 ;
			RECT	10.211 27.308 10.243 27.372 ;
			RECT	10.379 27.308 10.411 27.372 ;
			RECT	10.547 27.308 10.579 27.372 ;
			RECT	10.715 27.308 10.747 27.372 ;
			RECT	10.883 27.308 10.915 27.372 ;
			RECT	11.051 27.308 11.083 27.372 ;
			RECT	11.219 27.308 11.251 27.372 ;
			RECT	11.387 27.308 11.419 27.372 ;
			RECT	11.555 27.308 11.587 27.372 ;
			RECT	11.723 27.308 11.755 27.372 ;
			RECT	11.891 27.308 11.923 27.372 ;
			RECT	12.059 27.308 12.091 27.372 ;
			RECT	12.227 27.308 12.259 27.372 ;
			RECT	12.395 27.308 12.427 27.372 ;
			RECT	12.563 27.308 12.595 27.372 ;
			RECT	12.731 27.308 12.763 27.372 ;
			RECT	12.899 27.308 12.931 27.372 ;
			RECT	13.067 27.308 13.099 27.372 ;
			RECT	13.235 27.308 13.267 27.372 ;
			RECT	13.403 27.308 13.435 27.372 ;
			RECT	13.571 27.308 13.603 27.372 ;
			RECT	13.739 27.308 13.771 27.372 ;
			RECT	13.907 27.308 13.939 27.372 ;
			RECT	14.075 27.308 14.107 27.372 ;
			RECT	14.243 27.308 14.275 27.372 ;
			RECT	14.411 27.308 14.443 27.372 ;
			RECT	14.579 27.308 14.611 27.372 ;
			RECT	14.747 27.308 14.779 27.372 ;
			RECT	14.915 27.308 14.947 27.372 ;
			RECT	15.083 27.308 15.115 27.372 ;
			RECT	15.251 27.308 15.283 27.372 ;
			RECT	15.419 27.308 15.451 27.372 ;
			RECT	15.587 27.308 15.619 27.372 ;
			RECT	15.755 27.308 15.787 27.372 ;
			RECT	15.923 27.308 15.955 27.372 ;
			RECT	16.091 27.308 16.123 27.372 ;
			RECT	16.259 27.308 16.291 27.372 ;
			RECT	16.427 27.308 16.459 27.372 ;
			RECT	16.595 27.308 16.627 27.372 ;
			RECT	16.763 27.308 16.795 27.372 ;
			RECT	16.931 27.308 16.963 27.372 ;
			RECT	17.099 27.308 17.131 27.372 ;
			RECT	17.267 27.308 17.299 27.372 ;
			RECT	17.435 27.308 17.467 27.372 ;
			RECT	17.603 27.308 17.635 27.372 ;
			RECT	17.771 27.308 17.803 27.372 ;
			RECT	17.939 27.308 17.971 27.372 ;
			RECT	18.107 27.308 18.139 27.372 ;
			RECT	18.275 27.308 18.307 27.372 ;
			RECT	18.443 27.308 18.475 27.372 ;
			RECT	18.611 27.308 18.643 27.372 ;
			RECT	18.779 27.308 18.811 27.372 ;
			RECT	18.947 27.308 18.979 27.372 ;
			RECT	19.115 27.308 19.147 27.372 ;
			RECT	19.283 27.308 19.315 27.372 ;
			RECT	19.451 27.308 19.483 27.372 ;
			RECT	19.619 27.308 19.651 27.372 ;
			RECT	19.787 27.308 19.819 27.372 ;
			RECT	19.955 27.308 19.987 27.372 ;
			RECT	20.123 27.308 20.155 27.372 ;
			RECT	20.291 27.308 20.323 27.372 ;
			RECT	20.459 27.308 20.491 27.372 ;
			RECT	20.627 27.308 20.659 27.372 ;
			RECT	20.795 27.308 20.827 27.372 ;
			RECT	20.963 27.308 20.995 27.372 ;
			RECT	21.131 27.308 21.163 27.372 ;
			RECT	21.299 27.308 21.331 27.372 ;
			RECT	21.467 27.308 21.499 27.372 ;
			RECT	21.635 27.308 21.667 27.372 ;
			RECT	21.803 27.308 21.835 27.372 ;
			RECT	21.971 27.308 22.003 27.372 ;
			RECT	22.139 27.308 22.171 27.372 ;
			RECT	22.307 27.308 22.339 27.372 ;
			RECT	22.475 27.308 22.507 27.372 ;
			RECT	22.643 27.308 22.675 27.372 ;
			RECT	22.811 27.308 22.843 27.372 ;
			RECT	22.979 27.308 23.011 27.372 ;
			RECT	23.147 27.308 23.179 27.372 ;
			RECT	23.315 27.308 23.347 27.372 ;
			RECT	23.483 27.308 23.515 27.372 ;
			RECT	23.651 27.308 23.683 27.372 ;
			RECT	23.819 27.308 23.851 27.372 ;
			RECT	23.987 27.308 24.019 27.372 ;
			RECT	24.155 27.308 24.187 27.372 ;
			RECT	24.323 27.308 24.355 27.372 ;
			RECT	24.491 27.308 24.523 27.372 ;
			RECT	24.659 27.308 24.691 27.372 ;
			RECT	24.827 27.308 24.859 27.372 ;
			RECT	24.995 27.308 25.027 27.372 ;
			RECT	25.163 27.308 25.195 27.372 ;
			RECT	25.331 27.308 25.363 27.372 ;
			RECT	25.499 27.308 25.531 27.372 ;
			RECT	25.667 27.308 25.699 27.372 ;
			RECT	25.835 27.308 25.867 27.372 ;
			RECT	26.003 27.308 26.035 27.372 ;
			RECT	26.171 27.308 26.203 27.372 ;
			RECT	26.339 27.308 26.371 27.372 ;
			RECT	26.507 27.308 26.539 27.372 ;
			RECT	26.675 27.308 26.707 27.372 ;
			RECT	26.843 27.308 26.875 27.372 ;
			RECT	27.011 27.308 27.043 27.372 ;
			RECT	27.179 27.308 27.211 27.372 ;
			RECT	27.347 27.308 27.379 27.372 ;
			RECT	27.515 27.308 27.547 27.372 ;
			RECT	27.683 27.308 27.715 27.372 ;
			RECT	27.851 27.308 27.883 27.372 ;
			RECT	28.019 27.308 28.051 27.372 ;
			RECT	28.187 27.308 28.219 27.372 ;
			RECT	28.355 27.308 28.387 27.372 ;
			RECT	28.523 27.308 28.555 27.372 ;
			RECT	28.691 27.308 28.723 27.372 ;
			RECT	28.859 27.308 28.891 27.372 ;
			RECT	29.027 27.308 29.059 27.372 ;
			RECT	29.195 27.308 29.227 27.372 ;
			RECT	29.363 27.308 29.395 27.372 ;
			RECT	29.531 27.308 29.563 27.372 ;
			RECT	29.699 27.308 29.731 27.372 ;
			RECT	29.867 27.308 29.899 27.372 ;
			RECT	30.035 27.308 30.067 27.372 ;
			RECT	30.203 27.308 30.235 27.372 ;
			RECT	30.371 27.308 30.403 27.372 ;
			RECT	30.539 27.308 30.571 27.372 ;
			RECT	30.707 27.308 30.739 27.372 ;
			RECT	30.875 27.308 30.907 27.372 ;
			RECT	31.043 27.308 31.075 27.372 ;
			RECT	31.211 27.308 31.243 27.372 ;
			RECT	31.379 27.308 31.411 27.372 ;
			RECT	31.547 27.308 31.579 27.372 ;
			RECT	31.715 27.308 31.747 27.372 ;
			RECT	31.883 27.308 31.915 27.372 ;
			RECT	32.051 27.308 32.083 27.372 ;
			RECT	32.219 27.308 32.251 27.372 ;
			RECT	32.387 27.308 32.419 27.372 ;
			RECT	32.555 27.308 32.587 27.372 ;
			RECT	32.723 27.308 32.755 27.372 ;
			RECT	32.891 27.308 32.923 27.372 ;
			RECT	33.059 27.308 33.091 27.372 ;
			RECT	33.227 27.308 33.259 27.372 ;
			RECT	33.395 27.308 33.427 27.372 ;
			RECT	33.563 27.308 33.595 27.372 ;
			RECT	33.731 27.308 33.763 27.372 ;
			RECT	33.899 27.308 33.931 27.372 ;
			RECT	34.067 27.308 34.099 27.372 ;
			RECT	34.235 27.308 34.267 27.372 ;
			RECT	34.403 27.308 34.435 27.372 ;
			RECT	34.571 27.308 34.603 27.372 ;
			RECT	34.739 27.308 34.771 27.372 ;
			RECT	34.907 27.308 34.939 27.372 ;
			RECT	35.075 27.308 35.107 27.372 ;
			RECT	35.243 27.308 35.275 27.372 ;
			RECT	35.411 27.308 35.443 27.372 ;
			RECT	35.579 27.308 35.611 27.372 ;
			RECT	35.747 27.308 35.779 27.372 ;
			RECT	35.915 27.308 35.947 27.372 ;
			RECT	36.083 27.308 36.115 27.372 ;
			RECT	36.251 27.308 36.283 27.372 ;
			RECT	36.419 27.308 36.451 27.372 ;
			RECT	36.587 27.308 36.619 27.372 ;
			RECT	36.755 27.308 36.787 27.372 ;
			RECT	36.923 27.308 36.955 27.372 ;
			RECT	37.091 27.308 37.123 27.372 ;
			RECT	37.259 27.308 37.291 27.372 ;
			RECT	37.427 27.308 37.459 27.372 ;
			RECT	37.595 27.308 37.627 27.372 ;
			RECT	37.763 27.308 37.795 27.372 ;
			RECT	37.931 27.308 37.963 27.372 ;
			RECT	38.099 27.308 38.131 27.372 ;
			RECT	38.267 27.308 38.299 27.372 ;
			RECT	38.435 27.308 38.467 27.372 ;
			RECT	38.603 27.308 38.635 27.372 ;
			RECT	38.771 27.308 38.803 27.372 ;
			RECT	38.939 27.308 38.971 27.372 ;
			RECT	39.107 27.308 39.139 27.372 ;
			RECT	39.275 27.308 39.307 27.372 ;
			RECT	39.443 27.308 39.475 27.372 ;
			RECT	39.611 27.308 39.643 27.372 ;
			RECT	39.779 27.308 39.811 27.372 ;
			RECT	39.947 27.308 39.979 27.372 ;
			RECT	40.115 27.308 40.147 27.372 ;
			RECT	40.283 27.308 40.315 27.372 ;
			RECT	40.451 27.308 40.483 27.372 ;
			RECT	40.619 27.308 40.651 27.372 ;
			RECT	40.787 27.308 40.819 27.372 ;
			RECT	40.955 27.308 40.987 27.372 ;
			RECT	41.123 27.308 41.155 27.372 ;
			RECT	41.291 27.308 41.323 27.372 ;
			RECT	41.459 27.308 41.491 27.372 ;
			RECT	41.627 27.308 41.659 27.372 ;
			RECT	41.795 27.308 41.827 27.372 ;
			RECT	41.963 27.308 41.995 27.372 ;
			RECT	42.131 27.308 42.163 27.372 ;
			RECT	42.299 27.308 42.331 27.372 ;
			RECT	42.467 27.308 42.499 27.372 ;
			RECT	42.635 27.308 42.667 27.372 ;
			RECT	42.803 27.308 42.835 27.372 ;
			RECT	42.971 27.308 43.003 27.372 ;
			RECT	43.139 27.308 43.171 27.372 ;
			RECT	43.307 27.308 43.339 27.372 ;
			RECT	43.475 27.308 43.507 27.372 ;
			RECT	43.643 27.308 43.675 27.372 ;
			RECT	43.811 27.308 43.843 27.372 ;
			RECT	43.979 27.308 44.011 27.372 ;
			RECT	44.147 27.308 44.179 27.372 ;
			RECT	44.315 27.308 44.347 27.372 ;
			RECT	44.483 27.308 44.515 27.372 ;
			RECT	44.651 27.308 44.683 27.372 ;
			RECT	44.819 27.308 44.851 27.372 ;
			RECT	44.987 27.308 45.019 27.372 ;
			RECT	45.155 27.308 45.187 27.372 ;
			RECT	45.323 27.308 45.355 27.372 ;
			RECT	45.491 27.308 45.523 27.372 ;
			RECT	45.659 27.308 45.691 27.372 ;
			RECT	45.827 27.308 45.859 27.372 ;
			RECT	45.995 27.308 46.027 27.372 ;
			RECT	46.163 27.308 46.195 27.372 ;
			RECT	46.331 27.308 46.363 27.372 ;
			RECT	46.499 27.308 46.531 27.372 ;
			RECT	46.667 27.308 46.699 27.372 ;
			RECT	46.835 27.308 46.867 27.372 ;
			RECT	47.003 27.308 47.035 27.372 ;
			RECT	47.171 27.308 47.203 27.372 ;
			RECT	47.339 27.308 47.371 27.372 ;
			RECT	47.507 27.308 47.539 27.372 ;
			RECT	47.675 27.308 47.707 27.372 ;
			RECT	47.843 27.308 47.875 27.372 ;
			RECT	48.011 27.308 48.043 27.372 ;
			RECT	48.179 27.308 48.211 27.372 ;
			RECT	48.347 27.308 48.379 27.372 ;
			RECT	48.515 27.308 48.547 27.372 ;
			RECT	48.683 27.308 48.715 27.372 ;
			RECT	48.851 27.308 48.883 27.372 ;
			RECT	49.019 27.308 49.051 27.372 ;
			RECT	49.187 27.308 49.219 27.372 ;
			RECT	49.318 27.324 49.35 27.356 ;
			RECT	49.439 27.324 49.471 27.356 ;
			RECT	49.569 27.308 49.601 27.372 ;
			RECT	51.881 27.308 51.913 27.372 ;
			RECT	53.132 27.308 53.196 27.372 ;
			RECT	53.812 27.308 53.844 27.372 ;
			RECT	54.251 27.308 54.283 27.372 ;
			RECT	55.562 27.308 55.626 27.372 ;
			RECT	58.603 27.308 58.635 27.372 ;
			RECT	58.733 27.324 58.765 27.356 ;
			RECT	58.854 27.324 58.886 27.356 ;
			RECT	58.985 27.308 59.017 27.372 ;
			RECT	59.153 27.308 59.185 27.372 ;
			RECT	59.321 27.308 59.353 27.372 ;
			RECT	59.489 27.308 59.521 27.372 ;
			RECT	59.657 27.308 59.689 27.372 ;
			RECT	59.825 27.308 59.857 27.372 ;
			RECT	59.993 27.308 60.025 27.372 ;
			RECT	60.161 27.308 60.193 27.372 ;
			RECT	60.329 27.308 60.361 27.372 ;
			RECT	60.497 27.308 60.529 27.372 ;
			RECT	60.665 27.308 60.697 27.372 ;
			RECT	60.833 27.308 60.865 27.372 ;
			RECT	61.001 27.308 61.033 27.372 ;
			RECT	61.169 27.308 61.201 27.372 ;
			RECT	61.337 27.308 61.369 27.372 ;
			RECT	61.505 27.308 61.537 27.372 ;
			RECT	61.673 27.308 61.705 27.372 ;
			RECT	61.841 27.308 61.873 27.372 ;
			RECT	62.009 27.308 62.041 27.372 ;
			RECT	62.177 27.308 62.209 27.372 ;
			RECT	62.345 27.308 62.377 27.372 ;
			RECT	62.513 27.308 62.545 27.372 ;
			RECT	62.681 27.308 62.713 27.372 ;
			RECT	62.849 27.308 62.881 27.372 ;
			RECT	63.017 27.308 63.049 27.372 ;
			RECT	63.185 27.308 63.217 27.372 ;
			RECT	63.353 27.308 63.385 27.372 ;
			RECT	63.521 27.308 63.553 27.372 ;
			RECT	63.689 27.308 63.721 27.372 ;
			RECT	63.857 27.308 63.889 27.372 ;
			RECT	64.025 27.308 64.057 27.372 ;
			RECT	64.193 27.308 64.225 27.372 ;
			RECT	64.361 27.308 64.393 27.372 ;
			RECT	64.529 27.308 64.561 27.372 ;
			RECT	64.697 27.308 64.729 27.372 ;
			RECT	64.865 27.308 64.897 27.372 ;
			RECT	65.033 27.308 65.065 27.372 ;
			RECT	65.201 27.308 65.233 27.372 ;
			RECT	65.369 27.308 65.401 27.372 ;
			RECT	65.537 27.308 65.569 27.372 ;
			RECT	65.705 27.308 65.737 27.372 ;
			RECT	65.873 27.308 65.905 27.372 ;
			RECT	66.041 27.308 66.073 27.372 ;
			RECT	66.209 27.308 66.241 27.372 ;
			RECT	66.377 27.308 66.409 27.372 ;
			RECT	66.545 27.308 66.577 27.372 ;
			RECT	66.713 27.308 66.745 27.372 ;
			RECT	66.881 27.308 66.913 27.372 ;
			RECT	67.049 27.308 67.081 27.372 ;
			RECT	67.217 27.308 67.249 27.372 ;
			RECT	67.385 27.308 67.417 27.372 ;
			RECT	67.553 27.308 67.585 27.372 ;
			RECT	67.721 27.308 67.753 27.372 ;
			RECT	67.889 27.308 67.921 27.372 ;
			RECT	68.057 27.308 68.089 27.372 ;
			RECT	68.225 27.308 68.257 27.372 ;
			RECT	68.393 27.308 68.425 27.372 ;
			RECT	68.561 27.308 68.593 27.372 ;
			RECT	68.729 27.308 68.761 27.372 ;
			RECT	68.897 27.308 68.929 27.372 ;
			RECT	69.065 27.308 69.097 27.372 ;
			RECT	69.233 27.308 69.265 27.372 ;
			RECT	69.401 27.308 69.433 27.372 ;
			RECT	69.569 27.308 69.601 27.372 ;
			RECT	69.737 27.308 69.769 27.372 ;
			RECT	69.905 27.308 69.937 27.372 ;
			RECT	70.073 27.308 70.105 27.372 ;
			RECT	70.241 27.308 70.273 27.372 ;
			RECT	70.409 27.308 70.441 27.372 ;
			RECT	70.577 27.308 70.609 27.372 ;
			RECT	70.745 27.308 70.777 27.372 ;
			RECT	70.913 27.308 70.945 27.372 ;
			RECT	71.081 27.308 71.113 27.372 ;
			RECT	71.249 27.308 71.281 27.372 ;
			RECT	71.417 27.308 71.449 27.372 ;
			RECT	71.585 27.308 71.617 27.372 ;
			RECT	71.753 27.308 71.785 27.372 ;
			RECT	71.921 27.308 71.953 27.372 ;
			RECT	72.089 27.308 72.121 27.372 ;
			RECT	72.257 27.308 72.289 27.372 ;
			RECT	72.425 27.308 72.457 27.372 ;
			RECT	72.593 27.308 72.625 27.372 ;
			RECT	72.761 27.308 72.793 27.372 ;
			RECT	72.929 27.308 72.961 27.372 ;
			RECT	73.097 27.308 73.129 27.372 ;
			RECT	73.265 27.308 73.297 27.372 ;
			RECT	73.433 27.308 73.465 27.372 ;
			RECT	73.601 27.308 73.633 27.372 ;
			RECT	73.769 27.308 73.801 27.372 ;
			RECT	73.937 27.308 73.969 27.372 ;
			RECT	74.105 27.308 74.137 27.372 ;
			RECT	74.273 27.308 74.305 27.372 ;
			RECT	74.441 27.308 74.473 27.372 ;
			RECT	74.609 27.308 74.641 27.372 ;
			RECT	74.777 27.308 74.809 27.372 ;
			RECT	74.945 27.308 74.977 27.372 ;
			RECT	75.113 27.308 75.145 27.372 ;
			RECT	75.281 27.308 75.313 27.372 ;
			RECT	75.449 27.308 75.481 27.372 ;
			RECT	75.617 27.308 75.649 27.372 ;
			RECT	75.785 27.308 75.817 27.372 ;
			RECT	75.953 27.308 75.985 27.372 ;
			RECT	76.121 27.308 76.153 27.372 ;
			RECT	76.289 27.308 76.321 27.372 ;
			RECT	76.457 27.308 76.489 27.372 ;
			RECT	76.625 27.308 76.657 27.372 ;
			RECT	76.793 27.308 76.825 27.372 ;
			RECT	76.961 27.308 76.993 27.372 ;
			RECT	77.129 27.308 77.161 27.372 ;
			RECT	77.297 27.308 77.329 27.372 ;
			RECT	77.465 27.308 77.497 27.372 ;
			RECT	77.633 27.308 77.665 27.372 ;
			RECT	77.801 27.308 77.833 27.372 ;
			RECT	77.969 27.308 78.001 27.372 ;
			RECT	78.137 27.308 78.169 27.372 ;
			RECT	78.305 27.308 78.337 27.372 ;
			RECT	78.473 27.308 78.505 27.372 ;
			RECT	78.641 27.308 78.673 27.372 ;
			RECT	78.809 27.308 78.841 27.372 ;
			RECT	78.977 27.308 79.009 27.372 ;
			RECT	79.145 27.308 79.177 27.372 ;
			RECT	79.313 27.308 79.345 27.372 ;
			RECT	79.481 27.308 79.513 27.372 ;
			RECT	79.649 27.308 79.681 27.372 ;
			RECT	79.817 27.308 79.849 27.372 ;
			RECT	79.985 27.308 80.017 27.372 ;
			RECT	80.153 27.308 80.185 27.372 ;
			RECT	80.321 27.308 80.353 27.372 ;
			RECT	80.489 27.308 80.521 27.372 ;
			RECT	80.657 27.308 80.689 27.372 ;
			RECT	80.825 27.308 80.857 27.372 ;
			RECT	80.993 27.308 81.025 27.372 ;
			RECT	81.161 27.308 81.193 27.372 ;
			RECT	81.329 27.308 81.361 27.372 ;
			RECT	81.497 27.308 81.529 27.372 ;
			RECT	81.665 27.308 81.697 27.372 ;
			RECT	81.833 27.308 81.865 27.372 ;
			RECT	82.001 27.308 82.033 27.372 ;
			RECT	82.169 27.308 82.201 27.372 ;
			RECT	82.337 27.308 82.369 27.372 ;
			RECT	82.505 27.308 82.537 27.372 ;
			RECT	82.673 27.308 82.705 27.372 ;
			RECT	82.841 27.308 82.873 27.372 ;
			RECT	83.009 27.308 83.041 27.372 ;
			RECT	83.177 27.308 83.209 27.372 ;
			RECT	83.345 27.308 83.377 27.372 ;
			RECT	83.513 27.308 83.545 27.372 ;
			RECT	83.681 27.308 83.713 27.372 ;
			RECT	83.849 27.308 83.881 27.372 ;
			RECT	84.017 27.308 84.049 27.372 ;
			RECT	84.185 27.308 84.217 27.372 ;
			RECT	84.353 27.308 84.385 27.372 ;
			RECT	84.521 27.308 84.553 27.372 ;
			RECT	84.689 27.308 84.721 27.372 ;
			RECT	84.857 27.308 84.889 27.372 ;
			RECT	85.025 27.308 85.057 27.372 ;
			RECT	85.193 27.308 85.225 27.372 ;
			RECT	85.361 27.308 85.393 27.372 ;
			RECT	85.529 27.308 85.561 27.372 ;
			RECT	85.697 27.308 85.729 27.372 ;
			RECT	85.865 27.308 85.897 27.372 ;
			RECT	86.033 27.308 86.065 27.372 ;
			RECT	86.201 27.308 86.233 27.372 ;
			RECT	86.369 27.308 86.401 27.372 ;
			RECT	86.537 27.308 86.569 27.372 ;
			RECT	86.705 27.308 86.737 27.372 ;
			RECT	86.873 27.308 86.905 27.372 ;
			RECT	87.041 27.308 87.073 27.372 ;
			RECT	87.209 27.308 87.241 27.372 ;
			RECT	87.377 27.308 87.409 27.372 ;
			RECT	87.545 27.308 87.577 27.372 ;
			RECT	87.713 27.308 87.745 27.372 ;
			RECT	87.881 27.308 87.913 27.372 ;
			RECT	88.049 27.308 88.081 27.372 ;
			RECT	88.217 27.308 88.249 27.372 ;
			RECT	88.385 27.308 88.417 27.372 ;
			RECT	88.553 27.308 88.585 27.372 ;
			RECT	88.721 27.308 88.753 27.372 ;
			RECT	88.889 27.308 88.921 27.372 ;
			RECT	89.057 27.308 89.089 27.372 ;
			RECT	89.225 27.308 89.257 27.372 ;
			RECT	89.393 27.308 89.425 27.372 ;
			RECT	89.561 27.308 89.593 27.372 ;
			RECT	89.729 27.308 89.761 27.372 ;
			RECT	89.897 27.308 89.929 27.372 ;
			RECT	90.065 27.308 90.097 27.372 ;
			RECT	90.233 27.308 90.265 27.372 ;
			RECT	90.401 27.308 90.433 27.372 ;
			RECT	90.569 27.308 90.601 27.372 ;
			RECT	90.737 27.308 90.769 27.372 ;
			RECT	90.905 27.308 90.937 27.372 ;
			RECT	91.073 27.308 91.105 27.372 ;
			RECT	91.241 27.308 91.273 27.372 ;
			RECT	91.409 27.308 91.441 27.372 ;
			RECT	91.577 27.308 91.609 27.372 ;
			RECT	91.745 27.308 91.777 27.372 ;
			RECT	91.913 27.308 91.945 27.372 ;
			RECT	92.081 27.308 92.113 27.372 ;
			RECT	92.249 27.308 92.281 27.372 ;
			RECT	92.417 27.308 92.449 27.372 ;
			RECT	92.585 27.308 92.617 27.372 ;
			RECT	92.753 27.308 92.785 27.372 ;
			RECT	92.921 27.308 92.953 27.372 ;
			RECT	93.089 27.308 93.121 27.372 ;
			RECT	93.257 27.308 93.289 27.372 ;
			RECT	93.425 27.308 93.457 27.372 ;
			RECT	93.593 27.308 93.625 27.372 ;
			RECT	93.761 27.308 93.793 27.372 ;
			RECT	93.929 27.308 93.961 27.372 ;
			RECT	94.097 27.308 94.129 27.372 ;
			RECT	94.265 27.308 94.297 27.372 ;
			RECT	94.433 27.308 94.465 27.372 ;
			RECT	94.601 27.308 94.633 27.372 ;
			RECT	94.769 27.308 94.801 27.372 ;
			RECT	94.937 27.308 94.969 27.372 ;
			RECT	95.105 27.308 95.137 27.372 ;
			RECT	95.273 27.308 95.305 27.372 ;
			RECT	95.441 27.308 95.473 27.372 ;
			RECT	95.609 27.308 95.641 27.372 ;
			RECT	95.777 27.308 95.809 27.372 ;
			RECT	95.945 27.308 95.977 27.372 ;
			RECT	96.113 27.308 96.145 27.372 ;
			RECT	96.281 27.308 96.313 27.372 ;
			RECT	96.449 27.308 96.481 27.372 ;
			RECT	96.617 27.308 96.649 27.372 ;
			RECT	96.785 27.308 96.817 27.372 ;
			RECT	96.953 27.308 96.985 27.372 ;
			RECT	97.121 27.308 97.153 27.372 ;
			RECT	97.289 27.308 97.321 27.372 ;
			RECT	97.457 27.308 97.489 27.372 ;
			RECT	97.625 27.308 97.657 27.372 ;
			RECT	97.793 27.308 97.825 27.372 ;
			RECT	97.961 27.308 97.993 27.372 ;
			RECT	98.129 27.308 98.161 27.372 ;
			RECT	98.297 27.308 98.329 27.372 ;
			RECT	98.465 27.308 98.497 27.372 ;
			RECT	98.633 27.308 98.665 27.372 ;
			RECT	98.801 27.308 98.833 27.372 ;
			RECT	98.969 27.308 99.001 27.372 ;
			RECT	99.137 27.308 99.169 27.372 ;
			RECT	99.305 27.308 99.337 27.372 ;
			RECT	99.473 27.308 99.505 27.372 ;
			RECT	99.641 27.308 99.673 27.372 ;
			RECT	99.809 27.308 99.841 27.372 ;
			RECT	99.977 27.308 100.009 27.372 ;
			RECT	100.145 27.308 100.177 27.372 ;
			RECT	100.313 27.308 100.345 27.372 ;
			RECT	100.481 27.308 100.513 27.372 ;
			RECT	100.649 27.308 100.681 27.372 ;
			RECT	100.817 27.308 100.849 27.372 ;
			RECT	100.985 27.308 101.017 27.372 ;
			RECT	101.153 27.308 101.185 27.372 ;
			RECT	101.321 27.308 101.353 27.372 ;
			RECT	101.489 27.308 101.521 27.372 ;
			RECT	101.657 27.308 101.689 27.372 ;
			RECT	101.825 27.308 101.857 27.372 ;
			RECT	101.993 27.308 102.025 27.372 ;
			RECT	102.123 27.324 102.155 27.356 ;
			RECT	102.245 27.329 102.277 27.361 ;
			RECT	102.375 27.308 102.407 27.372 ;
			RECT	103.795 27.308 103.827 27.372 ;
			RECT	103.925 27.329 103.957 27.361 ;
			RECT	104.047 27.324 104.079 27.356 ;
			RECT	104.177 27.308 104.209 27.372 ;
			RECT	104.345 27.308 104.377 27.372 ;
			RECT	104.513 27.308 104.545 27.372 ;
			RECT	104.681 27.308 104.713 27.372 ;
			RECT	104.849 27.308 104.881 27.372 ;
			RECT	105.017 27.308 105.049 27.372 ;
			RECT	105.185 27.308 105.217 27.372 ;
			RECT	105.353 27.308 105.385 27.372 ;
			RECT	105.521 27.308 105.553 27.372 ;
			RECT	105.689 27.308 105.721 27.372 ;
			RECT	105.857 27.308 105.889 27.372 ;
			RECT	106.025 27.308 106.057 27.372 ;
			RECT	106.193 27.308 106.225 27.372 ;
			RECT	106.361 27.308 106.393 27.372 ;
			RECT	106.529 27.308 106.561 27.372 ;
			RECT	106.697 27.308 106.729 27.372 ;
			RECT	106.865 27.308 106.897 27.372 ;
			RECT	107.033 27.308 107.065 27.372 ;
			RECT	107.201 27.308 107.233 27.372 ;
			RECT	107.369 27.308 107.401 27.372 ;
			RECT	107.537 27.308 107.569 27.372 ;
			RECT	107.705 27.308 107.737 27.372 ;
			RECT	107.873 27.308 107.905 27.372 ;
			RECT	108.041 27.308 108.073 27.372 ;
			RECT	108.209 27.308 108.241 27.372 ;
			RECT	108.377 27.308 108.409 27.372 ;
			RECT	108.545 27.308 108.577 27.372 ;
			RECT	108.713 27.308 108.745 27.372 ;
			RECT	108.881 27.308 108.913 27.372 ;
			RECT	109.049 27.308 109.081 27.372 ;
			RECT	109.217 27.308 109.249 27.372 ;
			RECT	109.385 27.308 109.417 27.372 ;
			RECT	109.553 27.308 109.585 27.372 ;
			RECT	109.721 27.308 109.753 27.372 ;
			RECT	109.889 27.308 109.921 27.372 ;
			RECT	110.057 27.308 110.089 27.372 ;
			RECT	110.225 27.308 110.257 27.372 ;
			RECT	110.393 27.308 110.425 27.372 ;
			RECT	110.561 27.308 110.593 27.372 ;
			RECT	110.729 27.308 110.761 27.372 ;
			RECT	110.897 27.308 110.929 27.372 ;
			RECT	111.065 27.308 111.097 27.372 ;
			RECT	111.233 27.308 111.265 27.372 ;
			RECT	111.401 27.308 111.433 27.372 ;
			RECT	111.569 27.308 111.601 27.372 ;
			RECT	111.737 27.308 111.769 27.372 ;
			RECT	111.905 27.308 111.937 27.372 ;
			RECT	112.073 27.308 112.105 27.372 ;
			RECT	112.241 27.308 112.273 27.372 ;
			RECT	112.409 27.308 112.441 27.372 ;
			RECT	112.577 27.308 112.609 27.372 ;
			RECT	112.745 27.308 112.777 27.372 ;
			RECT	112.913 27.308 112.945 27.372 ;
			RECT	113.081 27.308 113.113 27.372 ;
			RECT	113.249 27.308 113.281 27.372 ;
			RECT	113.417 27.308 113.449 27.372 ;
			RECT	113.585 27.308 113.617 27.372 ;
			RECT	113.753 27.308 113.785 27.372 ;
			RECT	113.921 27.308 113.953 27.372 ;
			RECT	114.089 27.308 114.121 27.372 ;
			RECT	114.257 27.308 114.289 27.372 ;
			RECT	114.425 27.308 114.457 27.372 ;
			RECT	114.593 27.308 114.625 27.372 ;
			RECT	114.761 27.308 114.793 27.372 ;
			RECT	114.929 27.308 114.961 27.372 ;
			RECT	115.097 27.308 115.129 27.372 ;
			RECT	115.265 27.308 115.297 27.372 ;
			RECT	115.433 27.308 115.465 27.372 ;
			RECT	115.601 27.308 115.633 27.372 ;
			RECT	115.769 27.308 115.801 27.372 ;
			RECT	115.937 27.308 115.969 27.372 ;
			RECT	116.105 27.308 116.137 27.372 ;
			RECT	116.273 27.308 116.305 27.372 ;
			RECT	116.441 27.308 116.473 27.372 ;
			RECT	116.609 27.308 116.641 27.372 ;
			RECT	116.777 27.308 116.809 27.372 ;
			RECT	116.945 27.308 116.977 27.372 ;
			RECT	117.113 27.308 117.145 27.372 ;
			RECT	117.281 27.308 117.313 27.372 ;
			RECT	117.449 27.308 117.481 27.372 ;
			RECT	117.617 27.308 117.649 27.372 ;
			RECT	117.785 27.308 117.817 27.372 ;
			RECT	117.953 27.308 117.985 27.372 ;
			RECT	118.121 27.308 118.153 27.372 ;
			RECT	118.289 27.308 118.321 27.372 ;
			RECT	118.457 27.308 118.489 27.372 ;
			RECT	118.625 27.308 118.657 27.372 ;
			RECT	118.793 27.308 118.825 27.372 ;
			RECT	118.961 27.308 118.993 27.372 ;
			RECT	119.129 27.308 119.161 27.372 ;
			RECT	119.297 27.308 119.329 27.372 ;
			RECT	119.465 27.308 119.497 27.372 ;
			RECT	119.633 27.308 119.665 27.372 ;
			RECT	119.801 27.308 119.833 27.372 ;
			RECT	119.969 27.308 120.001 27.372 ;
			RECT	120.137 27.308 120.169 27.372 ;
			RECT	120.305 27.308 120.337 27.372 ;
			RECT	120.473 27.308 120.505 27.372 ;
			RECT	120.641 27.308 120.673 27.372 ;
			RECT	120.809 27.308 120.841 27.372 ;
			RECT	120.977 27.308 121.009 27.372 ;
			RECT	121.145 27.308 121.177 27.372 ;
			RECT	121.313 27.308 121.345 27.372 ;
			RECT	121.481 27.308 121.513 27.372 ;
			RECT	121.649 27.308 121.681 27.372 ;
			RECT	121.817 27.308 121.849 27.372 ;
			RECT	121.985 27.308 122.017 27.372 ;
			RECT	122.153 27.308 122.185 27.372 ;
			RECT	122.321 27.308 122.353 27.372 ;
			RECT	122.489 27.308 122.521 27.372 ;
			RECT	122.657 27.308 122.689 27.372 ;
			RECT	122.825 27.308 122.857 27.372 ;
			RECT	122.993 27.308 123.025 27.372 ;
			RECT	123.161 27.308 123.193 27.372 ;
			RECT	123.329 27.308 123.361 27.372 ;
			RECT	123.497 27.308 123.529 27.372 ;
			RECT	123.665 27.308 123.697 27.372 ;
			RECT	123.833 27.308 123.865 27.372 ;
			RECT	124.001 27.308 124.033 27.372 ;
			RECT	124.169 27.308 124.201 27.372 ;
			RECT	124.337 27.308 124.369 27.372 ;
			RECT	124.505 27.308 124.537 27.372 ;
			RECT	124.673 27.308 124.705 27.372 ;
			RECT	124.841 27.308 124.873 27.372 ;
			RECT	125.009 27.308 125.041 27.372 ;
			RECT	125.177 27.308 125.209 27.372 ;
			RECT	125.345 27.308 125.377 27.372 ;
			RECT	125.513 27.308 125.545 27.372 ;
			RECT	125.681 27.308 125.713 27.372 ;
			RECT	125.849 27.308 125.881 27.372 ;
			RECT	126.017 27.308 126.049 27.372 ;
			RECT	126.185 27.308 126.217 27.372 ;
			RECT	126.353 27.308 126.385 27.372 ;
			RECT	126.521 27.308 126.553 27.372 ;
			RECT	126.689 27.308 126.721 27.372 ;
			RECT	126.857 27.308 126.889 27.372 ;
			RECT	127.025 27.308 127.057 27.372 ;
			RECT	127.193 27.308 127.225 27.372 ;
			RECT	127.361 27.308 127.393 27.372 ;
			RECT	127.529 27.308 127.561 27.372 ;
			RECT	127.697 27.308 127.729 27.372 ;
			RECT	127.865 27.308 127.897 27.372 ;
			RECT	128.033 27.308 128.065 27.372 ;
			RECT	128.201 27.308 128.233 27.372 ;
			RECT	128.369 27.308 128.401 27.372 ;
			RECT	128.537 27.308 128.569 27.372 ;
			RECT	128.705 27.308 128.737 27.372 ;
			RECT	128.873 27.308 128.905 27.372 ;
			RECT	129.041 27.308 129.073 27.372 ;
			RECT	129.209 27.308 129.241 27.372 ;
			RECT	129.377 27.308 129.409 27.372 ;
			RECT	129.545 27.308 129.577 27.372 ;
			RECT	129.713 27.308 129.745 27.372 ;
			RECT	129.881 27.308 129.913 27.372 ;
			RECT	130.049 27.308 130.081 27.372 ;
			RECT	130.217 27.308 130.249 27.372 ;
			RECT	130.385 27.308 130.417 27.372 ;
			RECT	130.553 27.308 130.585 27.372 ;
			RECT	130.721 27.308 130.753 27.372 ;
			RECT	130.889 27.308 130.921 27.372 ;
			RECT	131.057 27.308 131.089 27.372 ;
			RECT	131.225 27.308 131.257 27.372 ;
			RECT	131.393 27.308 131.425 27.372 ;
			RECT	131.561 27.308 131.593 27.372 ;
			RECT	131.729 27.308 131.761 27.372 ;
			RECT	131.897 27.308 131.929 27.372 ;
			RECT	132.065 27.308 132.097 27.372 ;
			RECT	132.233 27.308 132.265 27.372 ;
			RECT	132.401 27.308 132.433 27.372 ;
			RECT	132.569 27.308 132.601 27.372 ;
			RECT	132.737 27.308 132.769 27.372 ;
			RECT	132.905 27.308 132.937 27.372 ;
			RECT	133.073 27.308 133.105 27.372 ;
			RECT	133.241 27.308 133.273 27.372 ;
			RECT	133.409 27.308 133.441 27.372 ;
			RECT	133.577 27.308 133.609 27.372 ;
			RECT	133.745 27.308 133.777 27.372 ;
			RECT	133.913 27.308 133.945 27.372 ;
			RECT	134.081 27.308 134.113 27.372 ;
			RECT	134.249 27.308 134.281 27.372 ;
			RECT	134.417 27.308 134.449 27.372 ;
			RECT	134.585 27.308 134.617 27.372 ;
			RECT	134.753 27.308 134.785 27.372 ;
			RECT	134.921 27.308 134.953 27.372 ;
			RECT	135.089 27.308 135.121 27.372 ;
			RECT	135.257 27.308 135.289 27.372 ;
			RECT	135.425 27.308 135.457 27.372 ;
			RECT	135.593 27.308 135.625 27.372 ;
			RECT	135.761 27.308 135.793 27.372 ;
			RECT	135.929 27.308 135.961 27.372 ;
			RECT	136.097 27.308 136.129 27.372 ;
			RECT	136.265 27.308 136.297 27.372 ;
			RECT	136.433 27.308 136.465 27.372 ;
			RECT	136.601 27.308 136.633 27.372 ;
			RECT	136.769 27.308 136.801 27.372 ;
			RECT	136.937 27.308 136.969 27.372 ;
			RECT	137.105 27.308 137.137 27.372 ;
			RECT	137.273 27.308 137.305 27.372 ;
			RECT	137.441 27.308 137.473 27.372 ;
			RECT	137.609 27.308 137.641 27.372 ;
			RECT	137.777 27.308 137.809 27.372 ;
			RECT	137.945 27.308 137.977 27.372 ;
			RECT	138.113 27.308 138.145 27.372 ;
			RECT	138.281 27.308 138.313 27.372 ;
			RECT	138.449 27.308 138.481 27.372 ;
			RECT	138.617 27.308 138.649 27.372 ;
			RECT	138.785 27.308 138.817 27.372 ;
			RECT	138.953 27.308 138.985 27.372 ;
			RECT	139.121 27.308 139.153 27.372 ;
			RECT	139.289 27.308 139.321 27.372 ;
			RECT	139.457 27.308 139.489 27.372 ;
			RECT	139.625 27.308 139.657 27.372 ;
			RECT	139.793 27.308 139.825 27.372 ;
			RECT	139.961 27.308 139.993 27.372 ;
			RECT	140.129 27.308 140.161 27.372 ;
			RECT	140.297 27.308 140.329 27.372 ;
			RECT	140.465 27.308 140.497 27.372 ;
			RECT	140.633 27.308 140.665 27.372 ;
			RECT	140.801 27.308 140.833 27.372 ;
			RECT	140.969 27.308 141.001 27.372 ;
			RECT	141.137 27.308 141.169 27.372 ;
			RECT	141.305 27.308 141.337 27.372 ;
			RECT	141.473 27.308 141.505 27.372 ;
			RECT	141.641 27.308 141.673 27.372 ;
			RECT	141.809 27.308 141.841 27.372 ;
			RECT	141.977 27.308 142.009 27.372 ;
			RECT	142.145 27.308 142.177 27.372 ;
			RECT	142.313 27.308 142.345 27.372 ;
			RECT	142.481 27.308 142.513 27.372 ;
			RECT	142.649 27.308 142.681 27.372 ;
			RECT	142.817 27.308 142.849 27.372 ;
			RECT	142.985 27.308 143.017 27.372 ;
			RECT	143.153 27.308 143.185 27.372 ;
			RECT	143.321 27.308 143.353 27.372 ;
			RECT	143.489 27.308 143.521 27.372 ;
			RECT	143.657 27.308 143.689 27.372 ;
			RECT	143.825 27.308 143.857 27.372 ;
			RECT	143.993 27.308 144.025 27.372 ;
			RECT	144.161 27.308 144.193 27.372 ;
			RECT	144.329 27.308 144.361 27.372 ;
			RECT	144.497 27.308 144.529 27.372 ;
			RECT	144.665 27.308 144.697 27.372 ;
			RECT	144.833 27.308 144.865 27.372 ;
			RECT	145.001 27.308 145.033 27.372 ;
			RECT	145.169 27.308 145.201 27.372 ;
			RECT	145.337 27.308 145.369 27.372 ;
			RECT	145.505 27.308 145.537 27.372 ;
			RECT	145.673 27.308 145.705 27.372 ;
			RECT	145.841 27.308 145.873 27.372 ;
			RECT	146.009 27.308 146.041 27.372 ;
			RECT	146.177 27.308 146.209 27.372 ;
			RECT	146.345 27.308 146.377 27.372 ;
			RECT	146.513 27.308 146.545 27.372 ;
			RECT	146.681 27.308 146.713 27.372 ;
			RECT	146.849 27.308 146.881 27.372 ;
			RECT	147.017 27.308 147.049 27.372 ;
			RECT	147.185 27.308 147.217 27.372 ;
			RECT	147.316 27.324 147.348 27.356 ;
			RECT	147.437 27.324 147.469 27.356 ;
			RECT	147.567 27.308 147.599 27.372 ;
			RECT	149.879 27.308 149.911 27.372 ;
			RECT	151.13 27.308 151.194 27.372 ;
			RECT	151.81 27.308 151.842 27.372 ;
			RECT	152.249 27.308 152.281 27.372 ;
			RECT	153.56 27.308 153.624 27.372 ;
			RECT	156.601 27.308 156.633 27.372 ;
			RECT	156.731 27.324 156.763 27.356 ;
			RECT	156.852 27.324 156.884 27.356 ;
			RECT	156.983 27.308 157.015 27.372 ;
			RECT	157.151 27.308 157.183 27.372 ;
			RECT	157.319 27.308 157.351 27.372 ;
			RECT	157.487 27.308 157.519 27.372 ;
			RECT	157.655 27.308 157.687 27.372 ;
			RECT	157.823 27.308 157.855 27.372 ;
			RECT	157.991 27.308 158.023 27.372 ;
			RECT	158.159 27.308 158.191 27.372 ;
			RECT	158.327 27.308 158.359 27.372 ;
			RECT	158.495 27.308 158.527 27.372 ;
			RECT	158.663 27.308 158.695 27.372 ;
			RECT	158.831 27.308 158.863 27.372 ;
			RECT	158.999 27.308 159.031 27.372 ;
			RECT	159.167 27.308 159.199 27.372 ;
			RECT	159.335 27.308 159.367 27.372 ;
			RECT	159.503 27.308 159.535 27.372 ;
			RECT	159.671 27.308 159.703 27.372 ;
			RECT	159.839 27.308 159.871 27.372 ;
			RECT	160.007 27.308 160.039 27.372 ;
			RECT	160.175 27.308 160.207 27.372 ;
			RECT	160.343 27.308 160.375 27.372 ;
			RECT	160.511 27.308 160.543 27.372 ;
			RECT	160.679 27.308 160.711 27.372 ;
			RECT	160.847 27.308 160.879 27.372 ;
			RECT	161.015 27.308 161.047 27.372 ;
			RECT	161.183 27.308 161.215 27.372 ;
			RECT	161.351 27.308 161.383 27.372 ;
			RECT	161.519 27.308 161.551 27.372 ;
			RECT	161.687 27.308 161.719 27.372 ;
			RECT	161.855 27.308 161.887 27.372 ;
			RECT	162.023 27.308 162.055 27.372 ;
			RECT	162.191 27.308 162.223 27.372 ;
			RECT	162.359 27.308 162.391 27.372 ;
			RECT	162.527 27.308 162.559 27.372 ;
			RECT	162.695 27.308 162.727 27.372 ;
			RECT	162.863 27.308 162.895 27.372 ;
			RECT	163.031 27.308 163.063 27.372 ;
			RECT	163.199 27.308 163.231 27.372 ;
			RECT	163.367 27.308 163.399 27.372 ;
			RECT	163.535 27.308 163.567 27.372 ;
			RECT	163.703 27.308 163.735 27.372 ;
			RECT	163.871 27.308 163.903 27.372 ;
			RECT	164.039 27.308 164.071 27.372 ;
			RECT	164.207 27.308 164.239 27.372 ;
			RECT	164.375 27.308 164.407 27.372 ;
			RECT	164.543 27.308 164.575 27.372 ;
			RECT	164.711 27.308 164.743 27.372 ;
			RECT	164.879 27.308 164.911 27.372 ;
			RECT	165.047 27.308 165.079 27.372 ;
			RECT	165.215 27.308 165.247 27.372 ;
			RECT	165.383 27.308 165.415 27.372 ;
			RECT	165.551 27.308 165.583 27.372 ;
			RECT	165.719 27.308 165.751 27.372 ;
			RECT	165.887 27.308 165.919 27.372 ;
			RECT	166.055 27.308 166.087 27.372 ;
			RECT	166.223 27.308 166.255 27.372 ;
			RECT	166.391 27.308 166.423 27.372 ;
			RECT	166.559 27.308 166.591 27.372 ;
			RECT	166.727 27.308 166.759 27.372 ;
			RECT	166.895 27.308 166.927 27.372 ;
			RECT	167.063 27.308 167.095 27.372 ;
			RECT	167.231 27.308 167.263 27.372 ;
			RECT	167.399 27.308 167.431 27.372 ;
			RECT	167.567 27.308 167.599 27.372 ;
			RECT	167.735 27.308 167.767 27.372 ;
			RECT	167.903 27.308 167.935 27.372 ;
			RECT	168.071 27.308 168.103 27.372 ;
			RECT	168.239 27.308 168.271 27.372 ;
			RECT	168.407 27.308 168.439 27.372 ;
			RECT	168.575 27.308 168.607 27.372 ;
			RECT	168.743 27.308 168.775 27.372 ;
			RECT	168.911 27.308 168.943 27.372 ;
			RECT	169.079 27.308 169.111 27.372 ;
			RECT	169.247 27.308 169.279 27.372 ;
			RECT	169.415 27.308 169.447 27.372 ;
			RECT	169.583 27.308 169.615 27.372 ;
			RECT	169.751 27.308 169.783 27.372 ;
			RECT	169.919 27.308 169.951 27.372 ;
			RECT	170.087 27.308 170.119 27.372 ;
			RECT	170.255 27.308 170.287 27.372 ;
			RECT	170.423 27.308 170.455 27.372 ;
			RECT	170.591 27.308 170.623 27.372 ;
			RECT	170.759 27.308 170.791 27.372 ;
			RECT	170.927 27.308 170.959 27.372 ;
			RECT	171.095 27.308 171.127 27.372 ;
			RECT	171.263 27.308 171.295 27.372 ;
			RECT	171.431 27.308 171.463 27.372 ;
			RECT	171.599 27.308 171.631 27.372 ;
			RECT	171.767 27.308 171.799 27.372 ;
			RECT	171.935 27.308 171.967 27.372 ;
			RECT	172.103 27.308 172.135 27.372 ;
			RECT	172.271 27.308 172.303 27.372 ;
			RECT	172.439 27.308 172.471 27.372 ;
			RECT	172.607 27.308 172.639 27.372 ;
			RECT	172.775 27.308 172.807 27.372 ;
			RECT	172.943 27.308 172.975 27.372 ;
			RECT	173.111 27.308 173.143 27.372 ;
			RECT	173.279 27.308 173.311 27.372 ;
			RECT	173.447 27.308 173.479 27.372 ;
			RECT	173.615 27.308 173.647 27.372 ;
			RECT	173.783 27.308 173.815 27.372 ;
			RECT	173.951 27.308 173.983 27.372 ;
			RECT	174.119 27.308 174.151 27.372 ;
			RECT	174.287 27.308 174.319 27.372 ;
			RECT	174.455 27.308 174.487 27.372 ;
			RECT	174.623 27.308 174.655 27.372 ;
			RECT	174.791 27.308 174.823 27.372 ;
			RECT	174.959 27.308 174.991 27.372 ;
			RECT	175.127 27.308 175.159 27.372 ;
			RECT	175.295 27.308 175.327 27.372 ;
			RECT	175.463 27.308 175.495 27.372 ;
			RECT	175.631 27.308 175.663 27.372 ;
			RECT	175.799 27.308 175.831 27.372 ;
			RECT	175.967 27.308 175.999 27.372 ;
			RECT	176.135 27.308 176.167 27.372 ;
			RECT	176.303 27.308 176.335 27.372 ;
			RECT	176.471 27.308 176.503 27.372 ;
			RECT	176.639 27.308 176.671 27.372 ;
			RECT	176.807 27.308 176.839 27.372 ;
			RECT	176.975 27.308 177.007 27.372 ;
			RECT	177.143 27.308 177.175 27.372 ;
			RECT	177.311 27.308 177.343 27.372 ;
			RECT	177.479 27.308 177.511 27.372 ;
			RECT	177.647 27.308 177.679 27.372 ;
			RECT	177.815 27.308 177.847 27.372 ;
			RECT	177.983 27.308 178.015 27.372 ;
			RECT	178.151 27.308 178.183 27.372 ;
			RECT	178.319 27.308 178.351 27.372 ;
			RECT	178.487 27.308 178.519 27.372 ;
			RECT	178.655 27.308 178.687 27.372 ;
			RECT	178.823 27.308 178.855 27.372 ;
			RECT	178.991 27.308 179.023 27.372 ;
			RECT	179.159 27.308 179.191 27.372 ;
			RECT	179.327 27.308 179.359 27.372 ;
			RECT	179.495 27.308 179.527 27.372 ;
			RECT	179.663 27.308 179.695 27.372 ;
			RECT	179.831 27.308 179.863 27.372 ;
			RECT	179.999 27.308 180.031 27.372 ;
			RECT	180.167 27.308 180.199 27.372 ;
			RECT	180.335 27.308 180.367 27.372 ;
			RECT	180.503 27.308 180.535 27.372 ;
			RECT	180.671 27.308 180.703 27.372 ;
			RECT	180.839 27.308 180.871 27.372 ;
			RECT	181.007 27.308 181.039 27.372 ;
			RECT	181.175 27.308 181.207 27.372 ;
			RECT	181.343 27.308 181.375 27.372 ;
			RECT	181.511 27.308 181.543 27.372 ;
			RECT	181.679 27.308 181.711 27.372 ;
			RECT	181.847 27.308 181.879 27.372 ;
			RECT	182.015 27.308 182.047 27.372 ;
			RECT	182.183 27.308 182.215 27.372 ;
			RECT	182.351 27.308 182.383 27.372 ;
			RECT	182.519 27.308 182.551 27.372 ;
			RECT	182.687 27.308 182.719 27.372 ;
			RECT	182.855 27.308 182.887 27.372 ;
			RECT	183.023 27.308 183.055 27.372 ;
			RECT	183.191 27.308 183.223 27.372 ;
			RECT	183.359 27.308 183.391 27.372 ;
			RECT	183.527 27.308 183.559 27.372 ;
			RECT	183.695 27.308 183.727 27.372 ;
			RECT	183.863 27.308 183.895 27.372 ;
			RECT	184.031 27.308 184.063 27.372 ;
			RECT	184.199 27.308 184.231 27.372 ;
			RECT	184.367 27.308 184.399 27.372 ;
			RECT	184.535 27.308 184.567 27.372 ;
			RECT	184.703 27.308 184.735 27.372 ;
			RECT	184.871 27.308 184.903 27.372 ;
			RECT	185.039 27.308 185.071 27.372 ;
			RECT	185.207 27.308 185.239 27.372 ;
			RECT	185.375 27.308 185.407 27.372 ;
			RECT	185.543 27.308 185.575 27.372 ;
			RECT	185.711 27.308 185.743 27.372 ;
			RECT	185.879 27.308 185.911 27.372 ;
			RECT	186.047 27.308 186.079 27.372 ;
			RECT	186.215 27.308 186.247 27.372 ;
			RECT	186.383 27.308 186.415 27.372 ;
			RECT	186.551 27.308 186.583 27.372 ;
			RECT	186.719 27.308 186.751 27.372 ;
			RECT	186.887 27.308 186.919 27.372 ;
			RECT	187.055 27.308 187.087 27.372 ;
			RECT	187.223 27.308 187.255 27.372 ;
			RECT	187.391 27.308 187.423 27.372 ;
			RECT	187.559 27.308 187.591 27.372 ;
			RECT	187.727 27.308 187.759 27.372 ;
			RECT	187.895 27.308 187.927 27.372 ;
			RECT	188.063 27.308 188.095 27.372 ;
			RECT	188.231 27.308 188.263 27.372 ;
			RECT	188.399 27.308 188.431 27.372 ;
			RECT	188.567 27.308 188.599 27.372 ;
			RECT	188.735 27.308 188.767 27.372 ;
			RECT	188.903 27.308 188.935 27.372 ;
			RECT	189.071 27.308 189.103 27.372 ;
			RECT	189.239 27.308 189.271 27.372 ;
			RECT	189.407 27.308 189.439 27.372 ;
			RECT	189.575 27.308 189.607 27.372 ;
			RECT	189.743 27.308 189.775 27.372 ;
			RECT	189.911 27.308 189.943 27.372 ;
			RECT	190.079 27.308 190.111 27.372 ;
			RECT	190.247 27.308 190.279 27.372 ;
			RECT	190.415 27.308 190.447 27.372 ;
			RECT	190.583 27.308 190.615 27.372 ;
			RECT	190.751 27.308 190.783 27.372 ;
			RECT	190.919 27.308 190.951 27.372 ;
			RECT	191.087 27.308 191.119 27.372 ;
			RECT	191.255 27.308 191.287 27.372 ;
			RECT	191.423 27.308 191.455 27.372 ;
			RECT	191.591 27.308 191.623 27.372 ;
			RECT	191.759 27.308 191.791 27.372 ;
			RECT	191.927 27.308 191.959 27.372 ;
			RECT	192.095 27.308 192.127 27.372 ;
			RECT	192.263 27.308 192.295 27.372 ;
			RECT	192.431 27.308 192.463 27.372 ;
			RECT	192.599 27.308 192.631 27.372 ;
			RECT	192.767 27.308 192.799 27.372 ;
			RECT	192.935 27.308 192.967 27.372 ;
			RECT	193.103 27.308 193.135 27.372 ;
			RECT	193.271 27.308 193.303 27.372 ;
			RECT	193.439 27.308 193.471 27.372 ;
			RECT	193.607 27.308 193.639 27.372 ;
			RECT	193.775 27.308 193.807 27.372 ;
			RECT	193.943 27.308 193.975 27.372 ;
			RECT	194.111 27.308 194.143 27.372 ;
			RECT	194.279 27.308 194.311 27.372 ;
			RECT	194.447 27.308 194.479 27.372 ;
			RECT	194.615 27.308 194.647 27.372 ;
			RECT	194.783 27.308 194.815 27.372 ;
			RECT	194.951 27.308 194.983 27.372 ;
			RECT	195.119 27.308 195.151 27.372 ;
			RECT	195.287 27.308 195.319 27.372 ;
			RECT	195.455 27.308 195.487 27.372 ;
			RECT	195.623 27.308 195.655 27.372 ;
			RECT	195.791 27.308 195.823 27.372 ;
			RECT	195.959 27.308 195.991 27.372 ;
			RECT	196.127 27.308 196.159 27.372 ;
			RECT	196.295 27.308 196.327 27.372 ;
			RECT	196.463 27.308 196.495 27.372 ;
			RECT	196.631 27.308 196.663 27.372 ;
			RECT	196.799 27.308 196.831 27.372 ;
			RECT	196.967 27.308 196.999 27.372 ;
			RECT	197.135 27.308 197.167 27.372 ;
			RECT	197.303 27.308 197.335 27.372 ;
			RECT	197.471 27.308 197.503 27.372 ;
			RECT	197.639 27.308 197.671 27.372 ;
			RECT	197.807 27.308 197.839 27.372 ;
			RECT	197.975 27.308 198.007 27.372 ;
			RECT	198.143 27.308 198.175 27.372 ;
			RECT	198.311 27.308 198.343 27.372 ;
			RECT	198.479 27.308 198.511 27.372 ;
			RECT	198.647 27.308 198.679 27.372 ;
			RECT	198.815 27.308 198.847 27.372 ;
			RECT	198.983 27.308 199.015 27.372 ;
			RECT	199.151 27.308 199.183 27.372 ;
			RECT	199.319 27.308 199.351 27.372 ;
			RECT	199.487 27.308 199.519 27.372 ;
			RECT	199.655 27.308 199.687 27.372 ;
			RECT	199.823 27.308 199.855 27.372 ;
			RECT	199.991 27.308 200.023 27.372 ;
			RECT	200.121 27.324 200.153 27.356 ;
			RECT	200.243 27.329 200.275 27.361 ;
			RECT	200.373 27.308 200.405 27.372 ;
			RECT	200.9 27.308 200.932 27.372 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 25.36 201.665 25.48 ;
			LAYER	J3 ;
			RECT	0.755 25.388 0.787 25.452 ;
			RECT	1.645 25.388 1.709 25.452 ;
			RECT	2.323 25.388 2.387 25.452 ;
			RECT	3.438 25.388 3.47 25.452 ;
			RECT	3.585 25.388 3.617 25.452 ;
			RECT	4.195 25.388 4.227 25.452 ;
			RECT	4.72 25.388 4.752 25.452 ;
			RECT	4.944 25.388 5.008 25.452 ;
			RECT	5.267 25.388 5.299 25.452 ;
			RECT	5.797 25.388 5.829 25.452 ;
			RECT	5.927 25.409 5.959 25.441 ;
			RECT	6.049 25.404 6.081 25.436 ;
			RECT	6.179 25.388 6.211 25.452 ;
			RECT	6.347 25.388 6.379 25.452 ;
			RECT	6.515 25.388 6.547 25.452 ;
			RECT	6.683 25.388 6.715 25.452 ;
			RECT	6.851 25.388 6.883 25.452 ;
			RECT	7.019 25.388 7.051 25.452 ;
			RECT	7.187 25.388 7.219 25.452 ;
			RECT	7.355 25.388 7.387 25.452 ;
			RECT	7.523 25.388 7.555 25.452 ;
			RECT	7.691 25.388 7.723 25.452 ;
			RECT	7.859 25.388 7.891 25.452 ;
			RECT	8.027 25.388 8.059 25.452 ;
			RECT	8.195 25.388 8.227 25.452 ;
			RECT	8.363 25.388 8.395 25.452 ;
			RECT	8.531 25.388 8.563 25.452 ;
			RECT	8.699 25.388 8.731 25.452 ;
			RECT	8.867 25.388 8.899 25.452 ;
			RECT	9.035 25.388 9.067 25.452 ;
			RECT	9.203 25.388 9.235 25.452 ;
			RECT	9.371 25.388 9.403 25.452 ;
			RECT	9.539 25.388 9.571 25.452 ;
			RECT	9.707 25.388 9.739 25.452 ;
			RECT	9.875 25.388 9.907 25.452 ;
			RECT	10.043 25.388 10.075 25.452 ;
			RECT	10.211 25.388 10.243 25.452 ;
			RECT	10.379 25.388 10.411 25.452 ;
			RECT	10.547 25.388 10.579 25.452 ;
			RECT	10.715 25.388 10.747 25.452 ;
			RECT	10.883 25.388 10.915 25.452 ;
			RECT	11.051 25.388 11.083 25.452 ;
			RECT	11.219 25.388 11.251 25.452 ;
			RECT	11.387 25.388 11.419 25.452 ;
			RECT	11.555 25.388 11.587 25.452 ;
			RECT	11.723 25.388 11.755 25.452 ;
			RECT	11.891 25.388 11.923 25.452 ;
			RECT	12.059 25.388 12.091 25.452 ;
			RECT	12.227 25.388 12.259 25.452 ;
			RECT	12.395 25.388 12.427 25.452 ;
			RECT	12.563 25.388 12.595 25.452 ;
			RECT	12.731 25.388 12.763 25.452 ;
			RECT	12.899 25.388 12.931 25.452 ;
			RECT	13.067 25.388 13.099 25.452 ;
			RECT	13.235 25.388 13.267 25.452 ;
			RECT	13.403 25.388 13.435 25.452 ;
			RECT	13.571 25.388 13.603 25.452 ;
			RECT	13.739 25.388 13.771 25.452 ;
			RECT	13.907 25.388 13.939 25.452 ;
			RECT	14.075 25.388 14.107 25.452 ;
			RECT	14.243 25.388 14.275 25.452 ;
			RECT	14.411 25.388 14.443 25.452 ;
			RECT	14.579 25.388 14.611 25.452 ;
			RECT	14.747 25.388 14.779 25.452 ;
			RECT	14.915 25.388 14.947 25.452 ;
			RECT	15.083 25.388 15.115 25.452 ;
			RECT	15.251 25.388 15.283 25.452 ;
			RECT	15.419 25.388 15.451 25.452 ;
			RECT	15.587 25.388 15.619 25.452 ;
			RECT	15.755 25.388 15.787 25.452 ;
			RECT	15.923 25.388 15.955 25.452 ;
			RECT	16.091 25.388 16.123 25.452 ;
			RECT	16.259 25.388 16.291 25.452 ;
			RECT	16.427 25.388 16.459 25.452 ;
			RECT	16.595 25.388 16.627 25.452 ;
			RECT	16.763 25.388 16.795 25.452 ;
			RECT	16.931 25.388 16.963 25.452 ;
			RECT	17.099 25.388 17.131 25.452 ;
			RECT	17.267 25.388 17.299 25.452 ;
			RECT	17.435 25.388 17.467 25.452 ;
			RECT	17.603 25.388 17.635 25.452 ;
			RECT	17.771 25.388 17.803 25.452 ;
			RECT	17.939 25.388 17.971 25.452 ;
			RECT	18.107 25.388 18.139 25.452 ;
			RECT	18.275 25.388 18.307 25.452 ;
			RECT	18.443 25.388 18.475 25.452 ;
			RECT	18.611 25.388 18.643 25.452 ;
			RECT	18.779 25.388 18.811 25.452 ;
			RECT	18.947 25.388 18.979 25.452 ;
			RECT	19.115 25.388 19.147 25.452 ;
			RECT	19.283 25.388 19.315 25.452 ;
			RECT	19.451 25.388 19.483 25.452 ;
			RECT	19.619 25.388 19.651 25.452 ;
			RECT	19.787 25.388 19.819 25.452 ;
			RECT	19.955 25.388 19.987 25.452 ;
			RECT	20.123 25.388 20.155 25.452 ;
			RECT	20.291 25.388 20.323 25.452 ;
			RECT	20.459 25.388 20.491 25.452 ;
			RECT	20.627 25.388 20.659 25.452 ;
			RECT	20.795 25.388 20.827 25.452 ;
			RECT	20.963 25.388 20.995 25.452 ;
			RECT	21.131 25.388 21.163 25.452 ;
			RECT	21.299 25.388 21.331 25.452 ;
			RECT	21.467 25.388 21.499 25.452 ;
			RECT	21.635 25.388 21.667 25.452 ;
			RECT	21.803 25.388 21.835 25.452 ;
			RECT	21.971 25.388 22.003 25.452 ;
			RECT	22.139 25.388 22.171 25.452 ;
			RECT	22.307 25.388 22.339 25.452 ;
			RECT	22.475 25.388 22.507 25.452 ;
			RECT	22.643 25.388 22.675 25.452 ;
			RECT	22.811 25.388 22.843 25.452 ;
			RECT	22.979 25.388 23.011 25.452 ;
			RECT	23.147 25.388 23.179 25.452 ;
			RECT	23.315 25.388 23.347 25.452 ;
			RECT	23.483 25.388 23.515 25.452 ;
			RECT	23.651 25.388 23.683 25.452 ;
			RECT	23.819 25.388 23.851 25.452 ;
			RECT	23.987 25.388 24.019 25.452 ;
			RECT	24.155 25.388 24.187 25.452 ;
			RECT	24.323 25.388 24.355 25.452 ;
			RECT	24.491 25.388 24.523 25.452 ;
			RECT	24.659 25.388 24.691 25.452 ;
			RECT	24.827 25.388 24.859 25.452 ;
			RECT	24.995 25.388 25.027 25.452 ;
			RECT	25.163 25.388 25.195 25.452 ;
			RECT	25.331 25.388 25.363 25.452 ;
			RECT	25.499 25.388 25.531 25.452 ;
			RECT	25.667 25.388 25.699 25.452 ;
			RECT	25.835 25.388 25.867 25.452 ;
			RECT	26.003 25.388 26.035 25.452 ;
			RECT	26.171 25.388 26.203 25.452 ;
			RECT	26.339 25.388 26.371 25.452 ;
			RECT	26.507 25.388 26.539 25.452 ;
			RECT	26.675 25.388 26.707 25.452 ;
			RECT	26.843 25.388 26.875 25.452 ;
			RECT	27.011 25.388 27.043 25.452 ;
			RECT	27.179 25.388 27.211 25.452 ;
			RECT	27.347 25.388 27.379 25.452 ;
			RECT	27.515 25.388 27.547 25.452 ;
			RECT	27.683 25.388 27.715 25.452 ;
			RECT	27.851 25.388 27.883 25.452 ;
			RECT	28.019 25.388 28.051 25.452 ;
			RECT	28.187 25.388 28.219 25.452 ;
			RECT	28.355 25.388 28.387 25.452 ;
			RECT	28.523 25.388 28.555 25.452 ;
			RECT	28.691 25.388 28.723 25.452 ;
			RECT	28.859 25.388 28.891 25.452 ;
			RECT	29.027 25.388 29.059 25.452 ;
			RECT	29.195 25.388 29.227 25.452 ;
			RECT	29.363 25.388 29.395 25.452 ;
			RECT	29.531 25.388 29.563 25.452 ;
			RECT	29.699 25.388 29.731 25.452 ;
			RECT	29.867 25.388 29.899 25.452 ;
			RECT	30.035 25.388 30.067 25.452 ;
			RECT	30.203 25.388 30.235 25.452 ;
			RECT	30.371 25.388 30.403 25.452 ;
			RECT	30.539 25.388 30.571 25.452 ;
			RECT	30.707 25.388 30.739 25.452 ;
			RECT	30.875 25.388 30.907 25.452 ;
			RECT	31.043 25.388 31.075 25.452 ;
			RECT	31.211 25.388 31.243 25.452 ;
			RECT	31.379 25.388 31.411 25.452 ;
			RECT	31.547 25.388 31.579 25.452 ;
			RECT	31.715 25.388 31.747 25.452 ;
			RECT	31.883 25.388 31.915 25.452 ;
			RECT	32.051 25.388 32.083 25.452 ;
			RECT	32.219 25.388 32.251 25.452 ;
			RECT	32.387 25.388 32.419 25.452 ;
			RECT	32.555 25.388 32.587 25.452 ;
			RECT	32.723 25.388 32.755 25.452 ;
			RECT	32.891 25.388 32.923 25.452 ;
			RECT	33.059 25.388 33.091 25.452 ;
			RECT	33.227 25.388 33.259 25.452 ;
			RECT	33.395 25.388 33.427 25.452 ;
			RECT	33.563 25.388 33.595 25.452 ;
			RECT	33.731 25.388 33.763 25.452 ;
			RECT	33.899 25.388 33.931 25.452 ;
			RECT	34.067 25.388 34.099 25.452 ;
			RECT	34.235 25.388 34.267 25.452 ;
			RECT	34.403 25.388 34.435 25.452 ;
			RECT	34.571 25.388 34.603 25.452 ;
			RECT	34.739 25.388 34.771 25.452 ;
			RECT	34.907 25.388 34.939 25.452 ;
			RECT	35.075 25.388 35.107 25.452 ;
			RECT	35.243 25.388 35.275 25.452 ;
			RECT	35.411 25.388 35.443 25.452 ;
			RECT	35.579 25.388 35.611 25.452 ;
			RECT	35.747 25.388 35.779 25.452 ;
			RECT	35.915 25.388 35.947 25.452 ;
			RECT	36.083 25.388 36.115 25.452 ;
			RECT	36.251 25.388 36.283 25.452 ;
			RECT	36.419 25.388 36.451 25.452 ;
			RECT	36.587 25.388 36.619 25.452 ;
			RECT	36.755 25.388 36.787 25.452 ;
			RECT	36.923 25.388 36.955 25.452 ;
			RECT	37.091 25.388 37.123 25.452 ;
			RECT	37.259 25.388 37.291 25.452 ;
			RECT	37.427 25.388 37.459 25.452 ;
			RECT	37.595 25.388 37.627 25.452 ;
			RECT	37.763 25.388 37.795 25.452 ;
			RECT	37.931 25.388 37.963 25.452 ;
			RECT	38.099 25.388 38.131 25.452 ;
			RECT	38.267 25.388 38.299 25.452 ;
			RECT	38.435 25.388 38.467 25.452 ;
			RECT	38.603 25.388 38.635 25.452 ;
			RECT	38.771 25.388 38.803 25.452 ;
			RECT	38.939 25.388 38.971 25.452 ;
			RECT	39.107 25.388 39.139 25.452 ;
			RECT	39.275 25.388 39.307 25.452 ;
			RECT	39.443 25.388 39.475 25.452 ;
			RECT	39.611 25.388 39.643 25.452 ;
			RECT	39.779 25.388 39.811 25.452 ;
			RECT	39.947 25.388 39.979 25.452 ;
			RECT	40.115 25.388 40.147 25.452 ;
			RECT	40.283 25.388 40.315 25.452 ;
			RECT	40.451 25.388 40.483 25.452 ;
			RECT	40.619 25.388 40.651 25.452 ;
			RECT	40.787 25.388 40.819 25.452 ;
			RECT	40.955 25.388 40.987 25.452 ;
			RECT	41.123 25.388 41.155 25.452 ;
			RECT	41.291 25.388 41.323 25.452 ;
			RECT	41.459 25.388 41.491 25.452 ;
			RECT	41.627 25.388 41.659 25.452 ;
			RECT	41.795 25.388 41.827 25.452 ;
			RECT	41.963 25.388 41.995 25.452 ;
			RECT	42.131 25.388 42.163 25.452 ;
			RECT	42.299 25.388 42.331 25.452 ;
			RECT	42.467 25.388 42.499 25.452 ;
			RECT	42.635 25.388 42.667 25.452 ;
			RECT	42.803 25.388 42.835 25.452 ;
			RECT	42.971 25.388 43.003 25.452 ;
			RECT	43.139 25.388 43.171 25.452 ;
			RECT	43.307 25.388 43.339 25.452 ;
			RECT	43.475 25.388 43.507 25.452 ;
			RECT	43.643 25.388 43.675 25.452 ;
			RECT	43.811 25.388 43.843 25.452 ;
			RECT	43.979 25.388 44.011 25.452 ;
			RECT	44.147 25.388 44.179 25.452 ;
			RECT	44.315 25.388 44.347 25.452 ;
			RECT	44.483 25.388 44.515 25.452 ;
			RECT	44.651 25.388 44.683 25.452 ;
			RECT	44.819 25.388 44.851 25.452 ;
			RECT	44.987 25.388 45.019 25.452 ;
			RECT	45.155 25.388 45.187 25.452 ;
			RECT	45.323 25.388 45.355 25.452 ;
			RECT	45.491 25.388 45.523 25.452 ;
			RECT	45.659 25.388 45.691 25.452 ;
			RECT	45.827 25.388 45.859 25.452 ;
			RECT	45.995 25.388 46.027 25.452 ;
			RECT	46.163 25.388 46.195 25.452 ;
			RECT	46.331 25.388 46.363 25.452 ;
			RECT	46.499 25.388 46.531 25.452 ;
			RECT	46.667 25.388 46.699 25.452 ;
			RECT	46.835 25.388 46.867 25.452 ;
			RECT	47.003 25.388 47.035 25.452 ;
			RECT	47.171 25.388 47.203 25.452 ;
			RECT	47.339 25.388 47.371 25.452 ;
			RECT	47.507 25.388 47.539 25.452 ;
			RECT	47.675 25.388 47.707 25.452 ;
			RECT	47.843 25.388 47.875 25.452 ;
			RECT	48.011 25.388 48.043 25.452 ;
			RECT	48.179 25.388 48.211 25.452 ;
			RECT	48.347 25.388 48.379 25.452 ;
			RECT	48.515 25.388 48.547 25.452 ;
			RECT	48.683 25.388 48.715 25.452 ;
			RECT	48.851 25.388 48.883 25.452 ;
			RECT	49.019 25.388 49.051 25.452 ;
			RECT	49.187 25.388 49.219 25.452 ;
			RECT	49.318 25.404 49.35 25.436 ;
			RECT	49.439 25.404 49.471 25.436 ;
			RECT	49.569 25.388 49.601 25.452 ;
			RECT	51.881 25.388 51.913 25.452 ;
			RECT	53.132 25.388 53.196 25.452 ;
			RECT	53.812 25.388 53.844 25.452 ;
			RECT	54.251 25.388 54.283 25.452 ;
			RECT	55.562 25.388 55.626 25.452 ;
			RECT	58.603 25.388 58.635 25.452 ;
			RECT	58.733 25.404 58.765 25.436 ;
			RECT	58.854 25.404 58.886 25.436 ;
			RECT	58.985 25.388 59.017 25.452 ;
			RECT	59.153 25.388 59.185 25.452 ;
			RECT	59.321 25.388 59.353 25.452 ;
			RECT	59.489 25.388 59.521 25.452 ;
			RECT	59.657 25.388 59.689 25.452 ;
			RECT	59.825 25.388 59.857 25.452 ;
			RECT	59.993 25.388 60.025 25.452 ;
			RECT	60.161 25.388 60.193 25.452 ;
			RECT	60.329 25.388 60.361 25.452 ;
			RECT	60.497 25.388 60.529 25.452 ;
			RECT	60.665 25.388 60.697 25.452 ;
			RECT	60.833 25.388 60.865 25.452 ;
			RECT	61.001 25.388 61.033 25.452 ;
			RECT	61.169 25.388 61.201 25.452 ;
			RECT	61.337 25.388 61.369 25.452 ;
			RECT	61.505 25.388 61.537 25.452 ;
			RECT	61.673 25.388 61.705 25.452 ;
			RECT	61.841 25.388 61.873 25.452 ;
			RECT	62.009 25.388 62.041 25.452 ;
			RECT	62.177 25.388 62.209 25.452 ;
			RECT	62.345 25.388 62.377 25.452 ;
			RECT	62.513 25.388 62.545 25.452 ;
			RECT	62.681 25.388 62.713 25.452 ;
			RECT	62.849 25.388 62.881 25.452 ;
			RECT	63.017 25.388 63.049 25.452 ;
			RECT	63.185 25.388 63.217 25.452 ;
			RECT	63.353 25.388 63.385 25.452 ;
			RECT	63.521 25.388 63.553 25.452 ;
			RECT	63.689 25.388 63.721 25.452 ;
			RECT	63.857 25.388 63.889 25.452 ;
			RECT	64.025 25.388 64.057 25.452 ;
			RECT	64.193 25.388 64.225 25.452 ;
			RECT	64.361 25.388 64.393 25.452 ;
			RECT	64.529 25.388 64.561 25.452 ;
			RECT	64.697 25.388 64.729 25.452 ;
			RECT	64.865 25.388 64.897 25.452 ;
			RECT	65.033 25.388 65.065 25.452 ;
			RECT	65.201 25.388 65.233 25.452 ;
			RECT	65.369 25.388 65.401 25.452 ;
			RECT	65.537 25.388 65.569 25.452 ;
			RECT	65.705 25.388 65.737 25.452 ;
			RECT	65.873 25.388 65.905 25.452 ;
			RECT	66.041 25.388 66.073 25.452 ;
			RECT	66.209 25.388 66.241 25.452 ;
			RECT	66.377 25.388 66.409 25.452 ;
			RECT	66.545 25.388 66.577 25.452 ;
			RECT	66.713 25.388 66.745 25.452 ;
			RECT	66.881 25.388 66.913 25.452 ;
			RECT	67.049 25.388 67.081 25.452 ;
			RECT	67.217 25.388 67.249 25.452 ;
			RECT	67.385 25.388 67.417 25.452 ;
			RECT	67.553 25.388 67.585 25.452 ;
			RECT	67.721 25.388 67.753 25.452 ;
			RECT	67.889 25.388 67.921 25.452 ;
			RECT	68.057 25.388 68.089 25.452 ;
			RECT	68.225 25.388 68.257 25.452 ;
			RECT	68.393 25.388 68.425 25.452 ;
			RECT	68.561 25.388 68.593 25.452 ;
			RECT	68.729 25.388 68.761 25.452 ;
			RECT	68.897 25.388 68.929 25.452 ;
			RECT	69.065 25.388 69.097 25.452 ;
			RECT	69.233 25.388 69.265 25.452 ;
			RECT	69.401 25.388 69.433 25.452 ;
			RECT	69.569 25.388 69.601 25.452 ;
			RECT	69.737 25.388 69.769 25.452 ;
			RECT	69.905 25.388 69.937 25.452 ;
			RECT	70.073 25.388 70.105 25.452 ;
			RECT	70.241 25.388 70.273 25.452 ;
			RECT	70.409 25.388 70.441 25.452 ;
			RECT	70.577 25.388 70.609 25.452 ;
			RECT	70.745 25.388 70.777 25.452 ;
			RECT	70.913 25.388 70.945 25.452 ;
			RECT	71.081 25.388 71.113 25.452 ;
			RECT	71.249 25.388 71.281 25.452 ;
			RECT	71.417 25.388 71.449 25.452 ;
			RECT	71.585 25.388 71.617 25.452 ;
			RECT	71.753 25.388 71.785 25.452 ;
			RECT	71.921 25.388 71.953 25.452 ;
			RECT	72.089 25.388 72.121 25.452 ;
			RECT	72.257 25.388 72.289 25.452 ;
			RECT	72.425 25.388 72.457 25.452 ;
			RECT	72.593 25.388 72.625 25.452 ;
			RECT	72.761 25.388 72.793 25.452 ;
			RECT	72.929 25.388 72.961 25.452 ;
			RECT	73.097 25.388 73.129 25.452 ;
			RECT	73.265 25.388 73.297 25.452 ;
			RECT	73.433 25.388 73.465 25.452 ;
			RECT	73.601 25.388 73.633 25.452 ;
			RECT	73.769 25.388 73.801 25.452 ;
			RECT	73.937 25.388 73.969 25.452 ;
			RECT	74.105 25.388 74.137 25.452 ;
			RECT	74.273 25.388 74.305 25.452 ;
			RECT	74.441 25.388 74.473 25.452 ;
			RECT	74.609 25.388 74.641 25.452 ;
			RECT	74.777 25.388 74.809 25.452 ;
			RECT	74.945 25.388 74.977 25.452 ;
			RECT	75.113 25.388 75.145 25.452 ;
			RECT	75.281 25.388 75.313 25.452 ;
			RECT	75.449 25.388 75.481 25.452 ;
			RECT	75.617 25.388 75.649 25.452 ;
			RECT	75.785 25.388 75.817 25.452 ;
			RECT	75.953 25.388 75.985 25.452 ;
			RECT	76.121 25.388 76.153 25.452 ;
			RECT	76.289 25.388 76.321 25.452 ;
			RECT	76.457 25.388 76.489 25.452 ;
			RECT	76.625 25.388 76.657 25.452 ;
			RECT	76.793 25.388 76.825 25.452 ;
			RECT	76.961 25.388 76.993 25.452 ;
			RECT	77.129 25.388 77.161 25.452 ;
			RECT	77.297 25.388 77.329 25.452 ;
			RECT	77.465 25.388 77.497 25.452 ;
			RECT	77.633 25.388 77.665 25.452 ;
			RECT	77.801 25.388 77.833 25.452 ;
			RECT	77.969 25.388 78.001 25.452 ;
			RECT	78.137 25.388 78.169 25.452 ;
			RECT	78.305 25.388 78.337 25.452 ;
			RECT	78.473 25.388 78.505 25.452 ;
			RECT	78.641 25.388 78.673 25.452 ;
			RECT	78.809 25.388 78.841 25.452 ;
			RECT	78.977 25.388 79.009 25.452 ;
			RECT	79.145 25.388 79.177 25.452 ;
			RECT	79.313 25.388 79.345 25.452 ;
			RECT	79.481 25.388 79.513 25.452 ;
			RECT	79.649 25.388 79.681 25.452 ;
			RECT	79.817 25.388 79.849 25.452 ;
			RECT	79.985 25.388 80.017 25.452 ;
			RECT	80.153 25.388 80.185 25.452 ;
			RECT	80.321 25.388 80.353 25.452 ;
			RECT	80.489 25.388 80.521 25.452 ;
			RECT	80.657 25.388 80.689 25.452 ;
			RECT	80.825 25.388 80.857 25.452 ;
			RECT	80.993 25.388 81.025 25.452 ;
			RECT	81.161 25.388 81.193 25.452 ;
			RECT	81.329 25.388 81.361 25.452 ;
			RECT	81.497 25.388 81.529 25.452 ;
			RECT	81.665 25.388 81.697 25.452 ;
			RECT	81.833 25.388 81.865 25.452 ;
			RECT	82.001 25.388 82.033 25.452 ;
			RECT	82.169 25.388 82.201 25.452 ;
			RECT	82.337 25.388 82.369 25.452 ;
			RECT	82.505 25.388 82.537 25.452 ;
			RECT	82.673 25.388 82.705 25.452 ;
			RECT	82.841 25.388 82.873 25.452 ;
			RECT	83.009 25.388 83.041 25.452 ;
			RECT	83.177 25.388 83.209 25.452 ;
			RECT	83.345 25.388 83.377 25.452 ;
			RECT	83.513 25.388 83.545 25.452 ;
			RECT	83.681 25.388 83.713 25.452 ;
			RECT	83.849 25.388 83.881 25.452 ;
			RECT	84.017 25.388 84.049 25.452 ;
			RECT	84.185 25.388 84.217 25.452 ;
			RECT	84.353 25.388 84.385 25.452 ;
			RECT	84.521 25.388 84.553 25.452 ;
			RECT	84.689 25.388 84.721 25.452 ;
			RECT	84.857 25.388 84.889 25.452 ;
			RECT	85.025 25.388 85.057 25.452 ;
			RECT	85.193 25.388 85.225 25.452 ;
			RECT	85.361 25.388 85.393 25.452 ;
			RECT	85.529 25.388 85.561 25.452 ;
			RECT	85.697 25.388 85.729 25.452 ;
			RECT	85.865 25.388 85.897 25.452 ;
			RECT	86.033 25.388 86.065 25.452 ;
			RECT	86.201 25.388 86.233 25.452 ;
			RECT	86.369 25.388 86.401 25.452 ;
			RECT	86.537 25.388 86.569 25.452 ;
			RECT	86.705 25.388 86.737 25.452 ;
			RECT	86.873 25.388 86.905 25.452 ;
			RECT	87.041 25.388 87.073 25.452 ;
			RECT	87.209 25.388 87.241 25.452 ;
			RECT	87.377 25.388 87.409 25.452 ;
			RECT	87.545 25.388 87.577 25.452 ;
			RECT	87.713 25.388 87.745 25.452 ;
			RECT	87.881 25.388 87.913 25.452 ;
			RECT	88.049 25.388 88.081 25.452 ;
			RECT	88.217 25.388 88.249 25.452 ;
			RECT	88.385 25.388 88.417 25.452 ;
			RECT	88.553 25.388 88.585 25.452 ;
			RECT	88.721 25.388 88.753 25.452 ;
			RECT	88.889 25.388 88.921 25.452 ;
			RECT	89.057 25.388 89.089 25.452 ;
			RECT	89.225 25.388 89.257 25.452 ;
			RECT	89.393 25.388 89.425 25.452 ;
			RECT	89.561 25.388 89.593 25.452 ;
			RECT	89.729 25.388 89.761 25.452 ;
			RECT	89.897 25.388 89.929 25.452 ;
			RECT	90.065 25.388 90.097 25.452 ;
			RECT	90.233 25.388 90.265 25.452 ;
			RECT	90.401 25.388 90.433 25.452 ;
			RECT	90.569 25.388 90.601 25.452 ;
			RECT	90.737 25.388 90.769 25.452 ;
			RECT	90.905 25.388 90.937 25.452 ;
			RECT	91.073 25.388 91.105 25.452 ;
			RECT	91.241 25.388 91.273 25.452 ;
			RECT	91.409 25.388 91.441 25.452 ;
			RECT	91.577 25.388 91.609 25.452 ;
			RECT	91.745 25.388 91.777 25.452 ;
			RECT	91.913 25.388 91.945 25.452 ;
			RECT	92.081 25.388 92.113 25.452 ;
			RECT	92.249 25.388 92.281 25.452 ;
			RECT	92.417 25.388 92.449 25.452 ;
			RECT	92.585 25.388 92.617 25.452 ;
			RECT	92.753 25.388 92.785 25.452 ;
			RECT	92.921 25.388 92.953 25.452 ;
			RECT	93.089 25.388 93.121 25.452 ;
			RECT	93.257 25.388 93.289 25.452 ;
			RECT	93.425 25.388 93.457 25.452 ;
			RECT	93.593 25.388 93.625 25.452 ;
			RECT	93.761 25.388 93.793 25.452 ;
			RECT	93.929 25.388 93.961 25.452 ;
			RECT	94.097 25.388 94.129 25.452 ;
			RECT	94.265 25.388 94.297 25.452 ;
			RECT	94.433 25.388 94.465 25.452 ;
			RECT	94.601 25.388 94.633 25.452 ;
			RECT	94.769 25.388 94.801 25.452 ;
			RECT	94.937 25.388 94.969 25.452 ;
			RECT	95.105 25.388 95.137 25.452 ;
			RECT	95.273 25.388 95.305 25.452 ;
			RECT	95.441 25.388 95.473 25.452 ;
			RECT	95.609 25.388 95.641 25.452 ;
			RECT	95.777 25.388 95.809 25.452 ;
			RECT	95.945 25.388 95.977 25.452 ;
			RECT	96.113 25.388 96.145 25.452 ;
			RECT	96.281 25.388 96.313 25.452 ;
			RECT	96.449 25.388 96.481 25.452 ;
			RECT	96.617 25.388 96.649 25.452 ;
			RECT	96.785 25.388 96.817 25.452 ;
			RECT	96.953 25.388 96.985 25.452 ;
			RECT	97.121 25.388 97.153 25.452 ;
			RECT	97.289 25.388 97.321 25.452 ;
			RECT	97.457 25.388 97.489 25.452 ;
			RECT	97.625 25.388 97.657 25.452 ;
			RECT	97.793 25.388 97.825 25.452 ;
			RECT	97.961 25.388 97.993 25.452 ;
			RECT	98.129 25.388 98.161 25.452 ;
			RECT	98.297 25.388 98.329 25.452 ;
			RECT	98.465 25.388 98.497 25.452 ;
			RECT	98.633 25.388 98.665 25.452 ;
			RECT	98.801 25.388 98.833 25.452 ;
			RECT	98.969 25.388 99.001 25.452 ;
			RECT	99.137 25.388 99.169 25.452 ;
			RECT	99.305 25.388 99.337 25.452 ;
			RECT	99.473 25.388 99.505 25.452 ;
			RECT	99.641 25.388 99.673 25.452 ;
			RECT	99.809 25.388 99.841 25.452 ;
			RECT	99.977 25.388 100.009 25.452 ;
			RECT	100.145 25.388 100.177 25.452 ;
			RECT	100.313 25.388 100.345 25.452 ;
			RECT	100.481 25.388 100.513 25.452 ;
			RECT	100.649 25.388 100.681 25.452 ;
			RECT	100.817 25.388 100.849 25.452 ;
			RECT	100.985 25.388 101.017 25.452 ;
			RECT	101.153 25.388 101.185 25.452 ;
			RECT	101.321 25.388 101.353 25.452 ;
			RECT	101.489 25.388 101.521 25.452 ;
			RECT	101.657 25.388 101.689 25.452 ;
			RECT	101.825 25.388 101.857 25.452 ;
			RECT	101.993 25.388 102.025 25.452 ;
			RECT	102.123 25.404 102.155 25.436 ;
			RECT	102.245 25.409 102.277 25.441 ;
			RECT	102.375 25.388 102.407 25.452 ;
			RECT	103.795 25.388 103.827 25.452 ;
			RECT	103.925 25.409 103.957 25.441 ;
			RECT	104.047 25.404 104.079 25.436 ;
			RECT	104.177 25.388 104.209 25.452 ;
			RECT	104.345 25.388 104.377 25.452 ;
			RECT	104.513 25.388 104.545 25.452 ;
			RECT	104.681 25.388 104.713 25.452 ;
			RECT	104.849 25.388 104.881 25.452 ;
			RECT	105.017 25.388 105.049 25.452 ;
			RECT	105.185 25.388 105.217 25.452 ;
			RECT	105.353 25.388 105.385 25.452 ;
			RECT	105.521 25.388 105.553 25.452 ;
			RECT	105.689 25.388 105.721 25.452 ;
			RECT	105.857 25.388 105.889 25.452 ;
			RECT	106.025 25.388 106.057 25.452 ;
			RECT	106.193 25.388 106.225 25.452 ;
			RECT	106.361 25.388 106.393 25.452 ;
			RECT	106.529 25.388 106.561 25.452 ;
			RECT	106.697 25.388 106.729 25.452 ;
			RECT	106.865 25.388 106.897 25.452 ;
			RECT	107.033 25.388 107.065 25.452 ;
			RECT	107.201 25.388 107.233 25.452 ;
			RECT	107.369 25.388 107.401 25.452 ;
			RECT	107.537 25.388 107.569 25.452 ;
			RECT	107.705 25.388 107.737 25.452 ;
			RECT	107.873 25.388 107.905 25.452 ;
			RECT	108.041 25.388 108.073 25.452 ;
			RECT	108.209 25.388 108.241 25.452 ;
			RECT	108.377 25.388 108.409 25.452 ;
			RECT	108.545 25.388 108.577 25.452 ;
			RECT	108.713 25.388 108.745 25.452 ;
			RECT	108.881 25.388 108.913 25.452 ;
			RECT	109.049 25.388 109.081 25.452 ;
			RECT	109.217 25.388 109.249 25.452 ;
			RECT	109.385 25.388 109.417 25.452 ;
			RECT	109.553 25.388 109.585 25.452 ;
			RECT	109.721 25.388 109.753 25.452 ;
			RECT	109.889 25.388 109.921 25.452 ;
			RECT	110.057 25.388 110.089 25.452 ;
			RECT	110.225 25.388 110.257 25.452 ;
			RECT	110.393 25.388 110.425 25.452 ;
			RECT	110.561 25.388 110.593 25.452 ;
			RECT	110.729 25.388 110.761 25.452 ;
			RECT	110.897 25.388 110.929 25.452 ;
			RECT	111.065 25.388 111.097 25.452 ;
			RECT	111.233 25.388 111.265 25.452 ;
			RECT	111.401 25.388 111.433 25.452 ;
			RECT	111.569 25.388 111.601 25.452 ;
			RECT	111.737 25.388 111.769 25.452 ;
			RECT	111.905 25.388 111.937 25.452 ;
			RECT	112.073 25.388 112.105 25.452 ;
			RECT	112.241 25.388 112.273 25.452 ;
			RECT	112.409 25.388 112.441 25.452 ;
			RECT	112.577 25.388 112.609 25.452 ;
			RECT	112.745 25.388 112.777 25.452 ;
			RECT	112.913 25.388 112.945 25.452 ;
			RECT	113.081 25.388 113.113 25.452 ;
			RECT	113.249 25.388 113.281 25.452 ;
			RECT	113.417 25.388 113.449 25.452 ;
			RECT	113.585 25.388 113.617 25.452 ;
			RECT	113.753 25.388 113.785 25.452 ;
			RECT	113.921 25.388 113.953 25.452 ;
			RECT	114.089 25.388 114.121 25.452 ;
			RECT	114.257 25.388 114.289 25.452 ;
			RECT	114.425 25.388 114.457 25.452 ;
			RECT	114.593 25.388 114.625 25.452 ;
			RECT	114.761 25.388 114.793 25.452 ;
			RECT	114.929 25.388 114.961 25.452 ;
			RECT	115.097 25.388 115.129 25.452 ;
			RECT	115.265 25.388 115.297 25.452 ;
			RECT	115.433 25.388 115.465 25.452 ;
			RECT	115.601 25.388 115.633 25.452 ;
			RECT	115.769 25.388 115.801 25.452 ;
			RECT	115.937 25.388 115.969 25.452 ;
			RECT	116.105 25.388 116.137 25.452 ;
			RECT	116.273 25.388 116.305 25.452 ;
			RECT	116.441 25.388 116.473 25.452 ;
			RECT	116.609 25.388 116.641 25.452 ;
			RECT	116.777 25.388 116.809 25.452 ;
			RECT	116.945 25.388 116.977 25.452 ;
			RECT	117.113 25.388 117.145 25.452 ;
			RECT	117.281 25.388 117.313 25.452 ;
			RECT	117.449 25.388 117.481 25.452 ;
			RECT	117.617 25.388 117.649 25.452 ;
			RECT	117.785 25.388 117.817 25.452 ;
			RECT	117.953 25.388 117.985 25.452 ;
			RECT	118.121 25.388 118.153 25.452 ;
			RECT	118.289 25.388 118.321 25.452 ;
			RECT	118.457 25.388 118.489 25.452 ;
			RECT	118.625 25.388 118.657 25.452 ;
			RECT	118.793 25.388 118.825 25.452 ;
			RECT	118.961 25.388 118.993 25.452 ;
			RECT	119.129 25.388 119.161 25.452 ;
			RECT	119.297 25.388 119.329 25.452 ;
			RECT	119.465 25.388 119.497 25.452 ;
			RECT	119.633 25.388 119.665 25.452 ;
			RECT	119.801 25.388 119.833 25.452 ;
			RECT	119.969 25.388 120.001 25.452 ;
			RECT	120.137 25.388 120.169 25.452 ;
			RECT	120.305 25.388 120.337 25.452 ;
			RECT	120.473 25.388 120.505 25.452 ;
			RECT	120.641 25.388 120.673 25.452 ;
			RECT	120.809 25.388 120.841 25.452 ;
			RECT	120.977 25.388 121.009 25.452 ;
			RECT	121.145 25.388 121.177 25.452 ;
			RECT	121.313 25.388 121.345 25.452 ;
			RECT	121.481 25.388 121.513 25.452 ;
			RECT	121.649 25.388 121.681 25.452 ;
			RECT	121.817 25.388 121.849 25.452 ;
			RECT	121.985 25.388 122.017 25.452 ;
			RECT	122.153 25.388 122.185 25.452 ;
			RECT	122.321 25.388 122.353 25.452 ;
			RECT	122.489 25.388 122.521 25.452 ;
			RECT	122.657 25.388 122.689 25.452 ;
			RECT	122.825 25.388 122.857 25.452 ;
			RECT	122.993 25.388 123.025 25.452 ;
			RECT	123.161 25.388 123.193 25.452 ;
			RECT	123.329 25.388 123.361 25.452 ;
			RECT	123.497 25.388 123.529 25.452 ;
			RECT	123.665 25.388 123.697 25.452 ;
			RECT	123.833 25.388 123.865 25.452 ;
			RECT	124.001 25.388 124.033 25.452 ;
			RECT	124.169 25.388 124.201 25.452 ;
			RECT	124.337 25.388 124.369 25.452 ;
			RECT	124.505 25.388 124.537 25.452 ;
			RECT	124.673 25.388 124.705 25.452 ;
			RECT	124.841 25.388 124.873 25.452 ;
			RECT	125.009 25.388 125.041 25.452 ;
			RECT	125.177 25.388 125.209 25.452 ;
			RECT	125.345 25.388 125.377 25.452 ;
			RECT	125.513 25.388 125.545 25.452 ;
			RECT	125.681 25.388 125.713 25.452 ;
			RECT	125.849 25.388 125.881 25.452 ;
			RECT	126.017 25.388 126.049 25.452 ;
			RECT	126.185 25.388 126.217 25.452 ;
			RECT	126.353 25.388 126.385 25.452 ;
			RECT	126.521 25.388 126.553 25.452 ;
			RECT	126.689 25.388 126.721 25.452 ;
			RECT	126.857 25.388 126.889 25.452 ;
			RECT	127.025 25.388 127.057 25.452 ;
			RECT	127.193 25.388 127.225 25.452 ;
			RECT	127.361 25.388 127.393 25.452 ;
			RECT	127.529 25.388 127.561 25.452 ;
			RECT	127.697 25.388 127.729 25.452 ;
			RECT	127.865 25.388 127.897 25.452 ;
			RECT	128.033 25.388 128.065 25.452 ;
			RECT	128.201 25.388 128.233 25.452 ;
			RECT	128.369 25.388 128.401 25.452 ;
			RECT	128.537 25.388 128.569 25.452 ;
			RECT	128.705 25.388 128.737 25.452 ;
			RECT	128.873 25.388 128.905 25.452 ;
			RECT	129.041 25.388 129.073 25.452 ;
			RECT	129.209 25.388 129.241 25.452 ;
			RECT	129.377 25.388 129.409 25.452 ;
			RECT	129.545 25.388 129.577 25.452 ;
			RECT	129.713 25.388 129.745 25.452 ;
			RECT	129.881 25.388 129.913 25.452 ;
			RECT	130.049 25.388 130.081 25.452 ;
			RECT	130.217 25.388 130.249 25.452 ;
			RECT	130.385 25.388 130.417 25.452 ;
			RECT	130.553 25.388 130.585 25.452 ;
			RECT	130.721 25.388 130.753 25.452 ;
			RECT	130.889 25.388 130.921 25.452 ;
			RECT	131.057 25.388 131.089 25.452 ;
			RECT	131.225 25.388 131.257 25.452 ;
			RECT	131.393 25.388 131.425 25.452 ;
			RECT	131.561 25.388 131.593 25.452 ;
			RECT	131.729 25.388 131.761 25.452 ;
			RECT	131.897 25.388 131.929 25.452 ;
			RECT	132.065 25.388 132.097 25.452 ;
			RECT	132.233 25.388 132.265 25.452 ;
			RECT	132.401 25.388 132.433 25.452 ;
			RECT	132.569 25.388 132.601 25.452 ;
			RECT	132.737 25.388 132.769 25.452 ;
			RECT	132.905 25.388 132.937 25.452 ;
			RECT	133.073 25.388 133.105 25.452 ;
			RECT	133.241 25.388 133.273 25.452 ;
			RECT	133.409 25.388 133.441 25.452 ;
			RECT	133.577 25.388 133.609 25.452 ;
			RECT	133.745 25.388 133.777 25.452 ;
			RECT	133.913 25.388 133.945 25.452 ;
			RECT	134.081 25.388 134.113 25.452 ;
			RECT	134.249 25.388 134.281 25.452 ;
			RECT	134.417 25.388 134.449 25.452 ;
			RECT	134.585 25.388 134.617 25.452 ;
			RECT	134.753 25.388 134.785 25.452 ;
			RECT	134.921 25.388 134.953 25.452 ;
			RECT	135.089 25.388 135.121 25.452 ;
			RECT	135.257 25.388 135.289 25.452 ;
			RECT	135.425 25.388 135.457 25.452 ;
			RECT	135.593 25.388 135.625 25.452 ;
			RECT	135.761 25.388 135.793 25.452 ;
			RECT	135.929 25.388 135.961 25.452 ;
			RECT	136.097 25.388 136.129 25.452 ;
			RECT	136.265 25.388 136.297 25.452 ;
			RECT	136.433 25.388 136.465 25.452 ;
			RECT	136.601 25.388 136.633 25.452 ;
			RECT	136.769 25.388 136.801 25.452 ;
			RECT	136.937 25.388 136.969 25.452 ;
			RECT	137.105 25.388 137.137 25.452 ;
			RECT	137.273 25.388 137.305 25.452 ;
			RECT	137.441 25.388 137.473 25.452 ;
			RECT	137.609 25.388 137.641 25.452 ;
			RECT	137.777 25.388 137.809 25.452 ;
			RECT	137.945 25.388 137.977 25.452 ;
			RECT	138.113 25.388 138.145 25.452 ;
			RECT	138.281 25.388 138.313 25.452 ;
			RECT	138.449 25.388 138.481 25.452 ;
			RECT	138.617 25.388 138.649 25.452 ;
			RECT	138.785 25.388 138.817 25.452 ;
			RECT	138.953 25.388 138.985 25.452 ;
			RECT	139.121 25.388 139.153 25.452 ;
			RECT	139.289 25.388 139.321 25.452 ;
			RECT	139.457 25.388 139.489 25.452 ;
			RECT	139.625 25.388 139.657 25.452 ;
			RECT	139.793 25.388 139.825 25.452 ;
			RECT	139.961 25.388 139.993 25.452 ;
			RECT	140.129 25.388 140.161 25.452 ;
			RECT	140.297 25.388 140.329 25.452 ;
			RECT	140.465 25.388 140.497 25.452 ;
			RECT	140.633 25.388 140.665 25.452 ;
			RECT	140.801 25.388 140.833 25.452 ;
			RECT	140.969 25.388 141.001 25.452 ;
			RECT	141.137 25.388 141.169 25.452 ;
			RECT	141.305 25.388 141.337 25.452 ;
			RECT	141.473 25.388 141.505 25.452 ;
			RECT	141.641 25.388 141.673 25.452 ;
			RECT	141.809 25.388 141.841 25.452 ;
			RECT	141.977 25.388 142.009 25.452 ;
			RECT	142.145 25.388 142.177 25.452 ;
			RECT	142.313 25.388 142.345 25.452 ;
			RECT	142.481 25.388 142.513 25.452 ;
			RECT	142.649 25.388 142.681 25.452 ;
			RECT	142.817 25.388 142.849 25.452 ;
			RECT	142.985 25.388 143.017 25.452 ;
			RECT	143.153 25.388 143.185 25.452 ;
			RECT	143.321 25.388 143.353 25.452 ;
			RECT	143.489 25.388 143.521 25.452 ;
			RECT	143.657 25.388 143.689 25.452 ;
			RECT	143.825 25.388 143.857 25.452 ;
			RECT	143.993 25.388 144.025 25.452 ;
			RECT	144.161 25.388 144.193 25.452 ;
			RECT	144.329 25.388 144.361 25.452 ;
			RECT	144.497 25.388 144.529 25.452 ;
			RECT	144.665 25.388 144.697 25.452 ;
			RECT	144.833 25.388 144.865 25.452 ;
			RECT	145.001 25.388 145.033 25.452 ;
			RECT	145.169 25.388 145.201 25.452 ;
			RECT	145.337 25.388 145.369 25.452 ;
			RECT	145.505 25.388 145.537 25.452 ;
			RECT	145.673 25.388 145.705 25.452 ;
			RECT	145.841 25.388 145.873 25.452 ;
			RECT	146.009 25.388 146.041 25.452 ;
			RECT	146.177 25.388 146.209 25.452 ;
			RECT	146.345 25.388 146.377 25.452 ;
			RECT	146.513 25.388 146.545 25.452 ;
			RECT	146.681 25.388 146.713 25.452 ;
			RECT	146.849 25.388 146.881 25.452 ;
			RECT	147.017 25.388 147.049 25.452 ;
			RECT	147.185 25.388 147.217 25.452 ;
			RECT	147.316 25.404 147.348 25.436 ;
			RECT	147.437 25.404 147.469 25.436 ;
			RECT	147.567 25.388 147.599 25.452 ;
			RECT	149.879 25.388 149.911 25.452 ;
			RECT	151.13 25.388 151.194 25.452 ;
			RECT	151.81 25.388 151.842 25.452 ;
			RECT	152.249 25.388 152.281 25.452 ;
			RECT	153.56 25.388 153.624 25.452 ;
			RECT	156.601 25.388 156.633 25.452 ;
			RECT	156.731 25.404 156.763 25.436 ;
			RECT	156.852 25.404 156.884 25.436 ;
			RECT	156.983 25.388 157.015 25.452 ;
			RECT	157.151 25.388 157.183 25.452 ;
			RECT	157.319 25.388 157.351 25.452 ;
			RECT	157.487 25.388 157.519 25.452 ;
			RECT	157.655 25.388 157.687 25.452 ;
			RECT	157.823 25.388 157.855 25.452 ;
			RECT	157.991 25.388 158.023 25.452 ;
			RECT	158.159 25.388 158.191 25.452 ;
			RECT	158.327 25.388 158.359 25.452 ;
			RECT	158.495 25.388 158.527 25.452 ;
			RECT	158.663 25.388 158.695 25.452 ;
			RECT	158.831 25.388 158.863 25.452 ;
			RECT	158.999 25.388 159.031 25.452 ;
			RECT	159.167 25.388 159.199 25.452 ;
			RECT	159.335 25.388 159.367 25.452 ;
			RECT	159.503 25.388 159.535 25.452 ;
			RECT	159.671 25.388 159.703 25.452 ;
			RECT	159.839 25.388 159.871 25.452 ;
			RECT	160.007 25.388 160.039 25.452 ;
			RECT	160.175 25.388 160.207 25.452 ;
			RECT	160.343 25.388 160.375 25.452 ;
			RECT	160.511 25.388 160.543 25.452 ;
			RECT	160.679 25.388 160.711 25.452 ;
			RECT	160.847 25.388 160.879 25.452 ;
			RECT	161.015 25.388 161.047 25.452 ;
			RECT	161.183 25.388 161.215 25.452 ;
			RECT	161.351 25.388 161.383 25.452 ;
			RECT	161.519 25.388 161.551 25.452 ;
			RECT	161.687 25.388 161.719 25.452 ;
			RECT	161.855 25.388 161.887 25.452 ;
			RECT	162.023 25.388 162.055 25.452 ;
			RECT	162.191 25.388 162.223 25.452 ;
			RECT	162.359 25.388 162.391 25.452 ;
			RECT	162.527 25.388 162.559 25.452 ;
			RECT	162.695 25.388 162.727 25.452 ;
			RECT	162.863 25.388 162.895 25.452 ;
			RECT	163.031 25.388 163.063 25.452 ;
			RECT	163.199 25.388 163.231 25.452 ;
			RECT	163.367 25.388 163.399 25.452 ;
			RECT	163.535 25.388 163.567 25.452 ;
			RECT	163.703 25.388 163.735 25.452 ;
			RECT	163.871 25.388 163.903 25.452 ;
			RECT	164.039 25.388 164.071 25.452 ;
			RECT	164.207 25.388 164.239 25.452 ;
			RECT	164.375 25.388 164.407 25.452 ;
			RECT	164.543 25.388 164.575 25.452 ;
			RECT	164.711 25.388 164.743 25.452 ;
			RECT	164.879 25.388 164.911 25.452 ;
			RECT	165.047 25.388 165.079 25.452 ;
			RECT	165.215 25.388 165.247 25.452 ;
			RECT	165.383 25.388 165.415 25.452 ;
			RECT	165.551 25.388 165.583 25.452 ;
			RECT	165.719 25.388 165.751 25.452 ;
			RECT	165.887 25.388 165.919 25.452 ;
			RECT	166.055 25.388 166.087 25.452 ;
			RECT	166.223 25.388 166.255 25.452 ;
			RECT	166.391 25.388 166.423 25.452 ;
			RECT	166.559 25.388 166.591 25.452 ;
			RECT	166.727 25.388 166.759 25.452 ;
			RECT	166.895 25.388 166.927 25.452 ;
			RECT	167.063 25.388 167.095 25.452 ;
			RECT	167.231 25.388 167.263 25.452 ;
			RECT	167.399 25.388 167.431 25.452 ;
			RECT	167.567 25.388 167.599 25.452 ;
			RECT	167.735 25.388 167.767 25.452 ;
			RECT	167.903 25.388 167.935 25.452 ;
			RECT	168.071 25.388 168.103 25.452 ;
			RECT	168.239 25.388 168.271 25.452 ;
			RECT	168.407 25.388 168.439 25.452 ;
			RECT	168.575 25.388 168.607 25.452 ;
			RECT	168.743 25.388 168.775 25.452 ;
			RECT	168.911 25.388 168.943 25.452 ;
			RECT	169.079 25.388 169.111 25.452 ;
			RECT	169.247 25.388 169.279 25.452 ;
			RECT	169.415 25.388 169.447 25.452 ;
			RECT	169.583 25.388 169.615 25.452 ;
			RECT	169.751 25.388 169.783 25.452 ;
			RECT	169.919 25.388 169.951 25.452 ;
			RECT	170.087 25.388 170.119 25.452 ;
			RECT	170.255 25.388 170.287 25.452 ;
			RECT	170.423 25.388 170.455 25.452 ;
			RECT	170.591 25.388 170.623 25.452 ;
			RECT	170.759 25.388 170.791 25.452 ;
			RECT	170.927 25.388 170.959 25.452 ;
			RECT	171.095 25.388 171.127 25.452 ;
			RECT	171.263 25.388 171.295 25.452 ;
			RECT	171.431 25.388 171.463 25.452 ;
			RECT	171.599 25.388 171.631 25.452 ;
			RECT	171.767 25.388 171.799 25.452 ;
			RECT	171.935 25.388 171.967 25.452 ;
			RECT	172.103 25.388 172.135 25.452 ;
			RECT	172.271 25.388 172.303 25.452 ;
			RECT	172.439 25.388 172.471 25.452 ;
			RECT	172.607 25.388 172.639 25.452 ;
			RECT	172.775 25.388 172.807 25.452 ;
			RECT	172.943 25.388 172.975 25.452 ;
			RECT	173.111 25.388 173.143 25.452 ;
			RECT	173.279 25.388 173.311 25.452 ;
			RECT	173.447 25.388 173.479 25.452 ;
			RECT	173.615 25.388 173.647 25.452 ;
			RECT	173.783 25.388 173.815 25.452 ;
			RECT	173.951 25.388 173.983 25.452 ;
			RECT	174.119 25.388 174.151 25.452 ;
			RECT	174.287 25.388 174.319 25.452 ;
			RECT	174.455 25.388 174.487 25.452 ;
			RECT	174.623 25.388 174.655 25.452 ;
			RECT	174.791 25.388 174.823 25.452 ;
			RECT	174.959 25.388 174.991 25.452 ;
			RECT	175.127 25.388 175.159 25.452 ;
			RECT	175.295 25.388 175.327 25.452 ;
			RECT	175.463 25.388 175.495 25.452 ;
			RECT	175.631 25.388 175.663 25.452 ;
			RECT	175.799 25.388 175.831 25.452 ;
			RECT	175.967 25.388 175.999 25.452 ;
			RECT	176.135 25.388 176.167 25.452 ;
			RECT	176.303 25.388 176.335 25.452 ;
			RECT	176.471 25.388 176.503 25.452 ;
			RECT	176.639 25.388 176.671 25.452 ;
			RECT	176.807 25.388 176.839 25.452 ;
			RECT	176.975 25.388 177.007 25.452 ;
			RECT	177.143 25.388 177.175 25.452 ;
			RECT	177.311 25.388 177.343 25.452 ;
			RECT	177.479 25.388 177.511 25.452 ;
			RECT	177.647 25.388 177.679 25.452 ;
			RECT	177.815 25.388 177.847 25.452 ;
			RECT	177.983 25.388 178.015 25.452 ;
			RECT	178.151 25.388 178.183 25.452 ;
			RECT	178.319 25.388 178.351 25.452 ;
			RECT	178.487 25.388 178.519 25.452 ;
			RECT	178.655 25.388 178.687 25.452 ;
			RECT	178.823 25.388 178.855 25.452 ;
			RECT	178.991 25.388 179.023 25.452 ;
			RECT	179.159 25.388 179.191 25.452 ;
			RECT	179.327 25.388 179.359 25.452 ;
			RECT	179.495 25.388 179.527 25.452 ;
			RECT	179.663 25.388 179.695 25.452 ;
			RECT	179.831 25.388 179.863 25.452 ;
			RECT	179.999 25.388 180.031 25.452 ;
			RECT	180.167 25.388 180.199 25.452 ;
			RECT	180.335 25.388 180.367 25.452 ;
			RECT	180.503 25.388 180.535 25.452 ;
			RECT	180.671 25.388 180.703 25.452 ;
			RECT	180.839 25.388 180.871 25.452 ;
			RECT	181.007 25.388 181.039 25.452 ;
			RECT	181.175 25.388 181.207 25.452 ;
			RECT	181.343 25.388 181.375 25.452 ;
			RECT	181.511 25.388 181.543 25.452 ;
			RECT	181.679 25.388 181.711 25.452 ;
			RECT	181.847 25.388 181.879 25.452 ;
			RECT	182.015 25.388 182.047 25.452 ;
			RECT	182.183 25.388 182.215 25.452 ;
			RECT	182.351 25.388 182.383 25.452 ;
			RECT	182.519 25.388 182.551 25.452 ;
			RECT	182.687 25.388 182.719 25.452 ;
			RECT	182.855 25.388 182.887 25.452 ;
			RECT	183.023 25.388 183.055 25.452 ;
			RECT	183.191 25.388 183.223 25.452 ;
			RECT	183.359 25.388 183.391 25.452 ;
			RECT	183.527 25.388 183.559 25.452 ;
			RECT	183.695 25.388 183.727 25.452 ;
			RECT	183.863 25.388 183.895 25.452 ;
			RECT	184.031 25.388 184.063 25.452 ;
			RECT	184.199 25.388 184.231 25.452 ;
			RECT	184.367 25.388 184.399 25.452 ;
			RECT	184.535 25.388 184.567 25.452 ;
			RECT	184.703 25.388 184.735 25.452 ;
			RECT	184.871 25.388 184.903 25.452 ;
			RECT	185.039 25.388 185.071 25.452 ;
			RECT	185.207 25.388 185.239 25.452 ;
			RECT	185.375 25.388 185.407 25.452 ;
			RECT	185.543 25.388 185.575 25.452 ;
			RECT	185.711 25.388 185.743 25.452 ;
			RECT	185.879 25.388 185.911 25.452 ;
			RECT	186.047 25.388 186.079 25.452 ;
			RECT	186.215 25.388 186.247 25.452 ;
			RECT	186.383 25.388 186.415 25.452 ;
			RECT	186.551 25.388 186.583 25.452 ;
			RECT	186.719 25.388 186.751 25.452 ;
			RECT	186.887 25.388 186.919 25.452 ;
			RECT	187.055 25.388 187.087 25.452 ;
			RECT	187.223 25.388 187.255 25.452 ;
			RECT	187.391 25.388 187.423 25.452 ;
			RECT	187.559 25.388 187.591 25.452 ;
			RECT	187.727 25.388 187.759 25.452 ;
			RECT	187.895 25.388 187.927 25.452 ;
			RECT	188.063 25.388 188.095 25.452 ;
			RECT	188.231 25.388 188.263 25.452 ;
			RECT	188.399 25.388 188.431 25.452 ;
			RECT	188.567 25.388 188.599 25.452 ;
			RECT	188.735 25.388 188.767 25.452 ;
			RECT	188.903 25.388 188.935 25.452 ;
			RECT	189.071 25.388 189.103 25.452 ;
			RECT	189.239 25.388 189.271 25.452 ;
			RECT	189.407 25.388 189.439 25.452 ;
			RECT	189.575 25.388 189.607 25.452 ;
			RECT	189.743 25.388 189.775 25.452 ;
			RECT	189.911 25.388 189.943 25.452 ;
			RECT	190.079 25.388 190.111 25.452 ;
			RECT	190.247 25.388 190.279 25.452 ;
			RECT	190.415 25.388 190.447 25.452 ;
			RECT	190.583 25.388 190.615 25.452 ;
			RECT	190.751 25.388 190.783 25.452 ;
			RECT	190.919 25.388 190.951 25.452 ;
			RECT	191.087 25.388 191.119 25.452 ;
			RECT	191.255 25.388 191.287 25.452 ;
			RECT	191.423 25.388 191.455 25.452 ;
			RECT	191.591 25.388 191.623 25.452 ;
			RECT	191.759 25.388 191.791 25.452 ;
			RECT	191.927 25.388 191.959 25.452 ;
			RECT	192.095 25.388 192.127 25.452 ;
			RECT	192.263 25.388 192.295 25.452 ;
			RECT	192.431 25.388 192.463 25.452 ;
			RECT	192.599 25.388 192.631 25.452 ;
			RECT	192.767 25.388 192.799 25.452 ;
			RECT	192.935 25.388 192.967 25.452 ;
			RECT	193.103 25.388 193.135 25.452 ;
			RECT	193.271 25.388 193.303 25.452 ;
			RECT	193.439 25.388 193.471 25.452 ;
			RECT	193.607 25.388 193.639 25.452 ;
			RECT	193.775 25.388 193.807 25.452 ;
			RECT	193.943 25.388 193.975 25.452 ;
			RECT	194.111 25.388 194.143 25.452 ;
			RECT	194.279 25.388 194.311 25.452 ;
			RECT	194.447 25.388 194.479 25.452 ;
			RECT	194.615 25.388 194.647 25.452 ;
			RECT	194.783 25.388 194.815 25.452 ;
			RECT	194.951 25.388 194.983 25.452 ;
			RECT	195.119 25.388 195.151 25.452 ;
			RECT	195.287 25.388 195.319 25.452 ;
			RECT	195.455 25.388 195.487 25.452 ;
			RECT	195.623 25.388 195.655 25.452 ;
			RECT	195.791 25.388 195.823 25.452 ;
			RECT	195.959 25.388 195.991 25.452 ;
			RECT	196.127 25.388 196.159 25.452 ;
			RECT	196.295 25.388 196.327 25.452 ;
			RECT	196.463 25.388 196.495 25.452 ;
			RECT	196.631 25.388 196.663 25.452 ;
			RECT	196.799 25.388 196.831 25.452 ;
			RECT	196.967 25.388 196.999 25.452 ;
			RECT	197.135 25.388 197.167 25.452 ;
			RECT	197.303 25.388 197.335 25.452 ;
			RECT	197.471 25.388 197.503 25.452 ;
			RECT	197.639 25.388 197.671 25.452 ;
			RECT	197.807 25.388 197.839 25.452 ;
			RECT	197.975 25.388 198.007 25.452 ;
			RECT	198.143 25.388 198.175 25.452 ;
			RECT	198.311 25.388 198.343 25.452 ;
			RECT	198.479 25.388 198.511 25.452 ;
			RECT	198.647 25.388 198.679 25.452 ;
			RECT	198.815 25.388 198.847 25.452 ;
			RECT	198.983 25.388 199.015 25.452 ;
			RECT	199.151 25.388 199.183 25.452 ;
			RECT	199.319 25.388 199.351 25.452 ;
			RECT	199.487 25.388 199.519 25.452 ;
			RECT	199.655 25.388 199.687 25.452 ;
			RECT	199.823 25.388 199.855 25.452 ;
			RECT	199.991 25.388 200.023 25.452 ;
			RECT	200.121 25.404 200.153 25.436 ;
			RECT	200.243 25.409 200.275 25.441 ;
			RECT	200.373 25.388 200.405 25.452 ;
			RECT	200.9 25.388 200.932 25.452 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 23.44 201.665 23.56 ;
			LAYER	J3 ;
			RECT	0.755 23.468 0.787 23.532 ;
			RECT	1.645 23.468 1.709 23.532 ;
			RECT	2.323 23.468 2.387 23.532 ;
			RECT	3.438 23.468 3.47 23.532 ;
			RECT	3.585 23.468 3.617 23.532 ;
			RECT	4.195 23.468 4.227 23.532 ;
			RECT	4.72 23.468 4.752 23.532 ;
			RECT	4.944 23.468 5.008 23.532 ;
			RECT	5.267 23.468 5.299 23.532 ;
			RECT	5.797 23.468 5.829 23.532 ;
			RECT	5.927 23.489 5.959 23.521 ;
			RECT	6.049 23.484 6.081 23.516 ;
			RECT	6.179 23.468 6.211 23.532 ;
			RECT	6.347 23.468 6.379 23.532 ;
			RECT	6.515 23.468 6.547 23.532 ;
			RECT	6.683 23.468 6.715 23.532 ;
			RECT	6.851 23.468 6.883 23.532 ;
			RECT	7.019 23.468 7.051 23.532 ;
			RECT	7.187 23.468 7.219 23.532 ;
			RECT	7.355 23.468 7.387 23.532 ;
			RECT	7.523 23.468 7.555 23.532 ;
			RECT	7.691 23.468 7.723 23.532 ;
			RECT	7.859 23.468 7.891 23.532 ;
			RECT	8.027 23.468 8.059 23.532 ;
			RECT	8.195 23.468 8.227 23.532 ;
			RECT	8.363 23.468 8.395 23.532 ;
			RECT	8.531 23.468 8.563 23.532 ;
			RECT	8.699 23.468 8.731 23.532 ;
			RECT	8.867 23.468 8.899 23.532 ;
			RECT	9.035 23.468 9.067 23.532 ;
			RECT	9.203 23.468 9.235 23.532 ;
			RECT	9.371 23.468 9.403 23.532 ;
			RECT	9.539 23.468 9.571 23.532 ;
			RECT	9.707 23.468 9.739 23.532 ;
			RECT	9.875 23.468 9.907 23.532 ;
			RECT	10.043 23.468 10.075 23.532 ;
			RECT	10.211 23.468 10.243 23.532 ;
			RECT	10.379 23.468 10.411 23.532 ;
			RECT	10.547 23.468 10.579 23.532 ;
			RECT	10.715 23.468 10.747 23.532 ;
			RECT	10.883 23.468 10.915 23.532 ;
			RECT	11.051 23.468 11.083 23.532 ;
			RECT	11.219 23.468 11.251 23.532 ;
			RECT	11.387 23.468 11.419 23.532 ;
			RECT	11.555 23.468 11.587 23.532 ;
			RECT	11.723 23.468 11.755 23.532 ;
			RECT	11.891 23.468 11.923 23.532 ;
			RECT	12.059 23.468 12.091 23.532 ;
			RECT	12.227 23.468 12.259 23.532 ;
			RECT	12.395 23.468 12.427 23.532 ;
			RECT	12.563 23.468 12.595 23.532 ;
			RECT	12.731 23.468 12.763 23.532 ;
			RECT	12.899 23.468 12.931 23.532 ;
			RECT	13.067 23.468 13.099 23.532 ;
			RECT	13.235 23.468 13.267 23.532 ;
			RECT	13.403 23.468 13.435 23.532 ;
			RECT	13.571 23.468 13.603 23.532 ;
			RECT	13.739 23.468 13.771 23.532 ;
			RECT	13.907 23.468 13.939 23.532 ;
			RECT	14.075 23.468 14.107 23.532 ;
			RECT	14.243 23.468 14.275 23.532 ;
			RECT	14.411 23.468 14.443 23.532 ;
			RECT	14.579 23.468 14.611 23.532 ;
			RECT	14.747 23.468 14.779 23.532 ;
			RECT	14.915 23.468 14.947 23.532 ;
			RECT	15.083 23.468 15.115 23.532 ;
			RECT	15.251 23.468 15.283 23.532 ;
			RECT	15.419 23.468 15.451 23.532 ;
			RECT	15.587 23.468 15.619 23.532 ;
			RECT	15.755 23.468 15.787 23.532 ;
			RECT	15.923 23.468 15.955 23.532 ;
			RECT	16.091 23.468 16.123 23.532 ;
			RECT	16.259 23.468 16.291 23.532 ;
			RECT	16.427 23.468 16.459 23.532 ;
			RECT	16.595 23.468 16.627 23.532 ;
			RECT	16.763 23.468 16.795 23.532 ;
			RECT	16.931 23.468 16.963 23.532 ;
			RECT	17.099 23.468 17.131 23.532 ;
			RECT	17.267 23.468 17.299 23.532 ;
			RECT	17.435 23.468 17.467 23.532 ;
			RECT	17.603 23.468 17.635 23.532 ;
			RECT	17.771 23.468 17.803 23.532 ;
			RECT	17.939 23.468 17.971 23.532 ;
			RECT	18.107 23.468 18.139 23.532 ;
			RECT	18.275 23.468 18.307 23.532 ;
			RECT	18.443 23.468 18.475 23.532 ;
			RECT	18.611 23.468 18.643 23.532 ;
			RECT	18.779 23.468 18.811 23.532 ;
			RECT	18.947 23.468 18.979 23.532 ;
			RECT	19.115 23.468 19.147 23.532 ;
			RECT	19.283 23.468 19.315 23.532 ;
			RECT	19.451 23.468 19.483 23.532 ;
			RECT	19.619 23.468 19.651 23.532 ;
			RECT	19.787 23.468 19.819 23.532 ;
			RECT	19.955 23.468 19.987 23.532 ;
			RECT	20.123 23.468 20.155 23.532 ;
			RECT	20.291 23.468 20.323 23.532 ;
			RECT	20.459 23.468 20.491 23.532 ;
			RECT	20.627 23.468 20.659 23.532 ;
			RECT	20.795 23.468 20.827 23.532 ;
			RECT	20.963 23.468 20.995 23.532 ;
			RECT	21.131 23.468 21.163 23.532 ;
			RECT	21.299 23.468 21.331 23.532 ;
			RECT	21.467 23.468 21.499 23.532 ;
			RECT	21.635 23.468 21.667 23.532 ;
			RECT	21.803 23.468 21.835 23.532 ;
			RECT	21.971 23.468 22.003 23.532 ;
			RECT	22.139 23.468 22.171 23.532 ;
			RECT	22.307 23.468 22.339 23.532 ;
			RECT	22.475 23.468 22.507 23.532 ;
			RECT	22.643 23.468 22.675 23.532 ;
			RECT	22.811 23.468 22.843 23.532 ;
			RECT	22.979 23.468 23.011 23.532 ;
			RECT	23.147 23.468 23.179 23.532 ;
			RECT	23.315 23.468 23.347 23.532 ;
			RECT	23.483 23.468 23.515 23.532 ;
			RECT	23.651 23.468 23.683 23.532 ;
			RECT	23.819 23.468 23.851 23.532 ;
			RECT	23.987 23.468 24.019 23.532 ;
			RECT	24.155 23.468 24.187 23.532 ;
			RECT	24.323 23.468 24.355 23.532 ;
			RECT	24.491 23.468 24.523 23.532 ;
			RECT	24.659 23.468 24.691 23.532 ;
			RECT	24.827 23.468 24.859 23.532 ;
			RECT	24.995 23.468 25.027 23.532 ;
			RECT	25.163 23.468 25.195 23.532 ;
			RECT	25.331 23.468 25.363 23.532 ;
			RECT	25.499 23.468 25.531 23.532 ;
			RECT	25.667 23.468 25.699 23.532 ;
			RECT	25.835 23.468 25.867 23.532 ;
			RECT	26.003 23.468 26.035 23.532 ;
			RECT	26.171 23.468 26.203 23.532 ;
			RECT	26.339 23.468 26.371 23.532 ;
			RECT	26.507 23.468 26.539 23.532 ;
			RECT	26.675 23.468 26.707 23.532 ;
			RECT	26.843 23.468 26.875 23.532 ;
			RECT	27.011 23.468 27.043 23.532 ;
			RECT	27.179 23.468 27.211 23.532 ;
			RECT	27.347 23.468 27.379 23.532 ;
			RECT	27.515 23.468 27.547 23.532 ;
			RECT	27.683 23.468 27.715 23.532 ;
			RECT	27.851 23.468 27.883 23.532 ;
			RECT	28.019 23.468 28.051 23.532 ;
			RECT	28.187 23.468 28.219 23.532 ;
			RECT	28.355 23.468 28.387 23.532 ;
			RECT	28.523 23.468 28.555 23.532 ;
			RECT	28.691 23.468 28.723 23.532 ;
			RECT	28.859 23.468 28.891 23.532 ;
			RECT	29.027 23.468 29.059 23.532 ;
			RECT	29.195 23.468 29.227 23.532 ;
			RECT	29.363 23.468 29.395 23.532 ;
			RECT	29.531 23.468 29.563 23.532 ;
			RECT	29.699 23.468 29.731 23.532 ;
			RECT	29.867 23.468 29.899 23.532 ;
			RECT	30.035 23.468 30.067 23.532 ;
			RECT	30.203 23.468 30.235 23.532 ;
			RECT	30.371 23.468 30.403 23.532 ;
			RECT	30.539 23.468 30.571 23.532 ;
			RECT	30.707 23.468 30.739 23.532 ;
			RECT	30.875 23.468 30.907 23.532 ;
			RECT	31.043 23.468 31.075 23.532 ;
			RECT	31.211 23.468 31.243 23.532 ;
			RECT	31.379 23.468 31.411 23.532 ;
			RECT	31.547 23.468 31.579 23.532 ;
			RECT	31.715 23.468 31.747 23.532 ;
			RECT	31.883 23.468 31.915 23.532 ;
			RECT	32.051 23.468 32.083 23.532 ;
			RECT	32.219 23.468 32.251 23.532 ;
			RECT	32.387 23.468 32.419 23.532 ;
			RECT	32.555 23.468 32.587 23.532 ;
			RECT	32.723 23.468 32.755 23.532 ;
			RECT	32.891 23.468 32.923 23.532 ;
			RECT	33.059 23.468 33.091 23.532 ;
			RECT	33.227 23.468 33.259 23.532 ;
			RECT	33.395 23.468 33.427 23.532 ;
			RECT	33.563 23.468 33.595 23.532 ;
			RECT	33.731 23.468 33.763 23.532 ;
			RECT	33.899 23.468 33.931 23.532 ;
			RECT	34.067 23.468 34.099 23.532 ;
			RECT	34.235 23.468 34.267 23.532 ;
			RECT	34.403 23.468 34.435 23.532 ;
			RECT	34.571 23.468 34.603 23.532 ;
			RECT	34.739 23.468 34.771 23.532 ;
			RECT	34.907 23.468 34.939 23.532 ;
			RECT	35.075 23.468 35.107 23.532 ;
			RECT	35.243 23.468 35.275 23.532 ;
			RECT	35.411 23.468 35.443 23.532 ;
			RECT	35.579 23.468 35.611 23.532 ;
			RECT	35.747 23.468 35.779 23.532 ;
			RECT	35.915 23.468 35.947 23.532 ;
			RECT	36.083 23.468 36.115 23.532 ;
			RECT	36.251 23.468 36.283 23.532 ;
			RECT	36.419 23.468 36.451 23.532 ;
			RECT	36.587 23.468 36.619 23.532 ;
			RECT	36.755 23.468 36.787 23.532 ;
			RECT	36.923 23.468 36.955 23.532 ;
			RECT	37.091 23.468 37.123 23.532 ;
			RECT	37.259 23.468 37.291 23.532 ;
			RECT	37.427 23.468 37.459 23.532 ;
			RECT	37.595 23.468 37.627 23.532 ;
			RECT	37.763 23.468 37.795 23.532 ;
			RECT	37.931 23.468 37.963 23.532 ;
			RECT	38.099 23.468 38.131 23.532 ;
			RECT	38.267 23.468 38.299 23.532 ;
			RECT	38.435 23.468 38.467 23.532 ;
			RECT	38.603 23.468 38.635 23.532 ;
			RECT	38.771 23.468 38.803 23.532 ;
			RECT	38.939 23.468 38.971 23.532 ;
			RECT	39.107 23.468 39.139 23.532 ;
			RECT	39.275 23.468 39.307 23.532 ;
			RECT	39.443 23.468 39.475 23.532 ;
			RECT	39.611 23.468 39.643 23.532 ;
			RECT	39.779 23.468 39.811 23.532 ;
			RECT	39.947 23.468 39.979 23.532 ;
			RECT	40.115 23.468 40.147 23.532 ;
			RECT	40.283 23.468 40.315 23.532 ;
			RECT	40.451 23.468 40.483 23.532 ;
			RECT	40.619 23.468 40.651 23.532 ;
			RECT	40.787 23.468 40.819 23.532 ;
			RECT	40.955 23.468 40.987 23.532 ;
			RECT	41.123 23.468 41.155 23.532 ;
			RECT	41.291 23.468 41.323 23.532 ;
			RECT	41.459 23.468 41.491 23.532 ;
			RECT	41.627 23.468 41.659 23.532 ;
			RECT	41.795 23.468 41.827 23.532 ;
			RECT	41.963 23.468 41.995 23.532 ;
			RECT	42.131 23.468 42.163 23.532 ;
			RECT	42.299 23.468 42.331 23.532 ;
			RECT	42.467 23.468 42.499 23.532 ;
			RECT	42.635 23.468 42.667 23.532 ;
			RECT	42.803 23.468 42.835 23.532 ;
			RECT	42.971 23.468 43.003 23.532 ;
			RECT	43.139 23.468 43.171 23.532 ;
			RECT	43.307 23.468 43.339 23.532 ;
			RECT	43.475 23.468 43.507 23.532 ;
			RECT	43.643 23.468 43.675 23.532 ;
			RECT	43.811 23.468 43.843 23.532 ;
			RECT	43.979 23.468 44.011 23.532 ;
			RECT	44.147 23.468 44.179 23.532 ;
			RECT	44.315 23.468 44.347 23.532 ;
			RECT	44.483 23.468 44.515 23.532 ;
			RECT	44.651 23.468 44.683 23.532 ;
			RECT	44.819 23.468 44.851 23.532 ;
			RECT	44.987 23.468 45.019 23.532 ;
			RECT	45.155 23.468 45.187 23.532 ;
			RECT	45.323 23.468 45.355 23.532 ;
			RECT	45.491 23.468 45.523 23.532 ;
			RECT	45.659 23.468 45.691 23.532 ;
			RECT	45.827 23.468 45.859 23.532 ;
			RECT	45.995 23.468 46.027 23.532 ;
			RECT	46.163 23.468 46.195 23.532 ;
			RECT	46.331 23.468 46.363 23.532 ;
			RECT	46.499 23.468 46.531 23.532 ;
			RECT	46.667 23.468 46.699 23.532 ;
			RECT	46.835 23.468 46.867 23.532 ;
			RECT	47.003 23.468 47.035 23.532 ;
			RECT	47.171 23.468 47.203 23.532 ;
			RECT	47.339 23.468 47.371 23.532 ;
			RECT	47.507 23.468 47.539 23.532 ;
			RECT	47.675 23.468 47.707 23.532 ;
			RECT	47.843 23.468 47.875 23.532 ;
			RECT	48.011 23.468 48.043 23.532 ;
			RECT	48.179 23.468 48.211 23.532 ;
			RECT	48.347 23.468 48.379 23.532 ;
			RECT	48.515 23.468 48.547 23.532 ;
			RECT	48.683 23.468 48.715 23.532 ;
			RECT	48.851 23.468 48.883 23.532 ;
			RECT	49.019 23.468 49.051 23.532 ;
			RECT	49.187 23.468 49.219 23.532 ;
			RECT	49.318 23.484 49.35 23.516 ;
			RECT	49.439 23.484 49.471 23.516 ;
			RECT	49.569 23.468 49.601 23.532 ;
			RECT	51.881 23.468 51.913 23.532 ;
			RECT	53.132 23.468 53.196 23.532 ;
			RECT	53.812 23.468 53.844 23.532 ;
			RECT	54.251 23.468 54.283 23.532 ;
			RECT	55.562 23.468 55.626 23.532 ;
			RECT	58.603 23.468 58.635 23.532 ;
			RECT	58.733 23.484 58.765 23.516 ;
			RECT	58.854 23.484 58.886 23.516 ;
			RECT	58.985 23.468 59.017 23.532 ;
			RECT	59.153 23.468 59.185 23.532 ;
			RECT	59.321 23.468 59.353 23.532 ;
			RECT	59.489 23.468 59.521 23.532 ;
			RECT	59.657 23.468 59.689 23.532 ;
			RECT	59.825 23.468 59.857 23.532 ;
			RECT	59.993 23.468 60.025 23.532 ;
			RECT	60.161 23.468 60.193 23.532 ;
			RECT	60.329 23.468 60.361 23.532 ;
			RECT	60.497 23.468 60.529 23.532 ;
			RECT	60.665 23.468 60.697 23.532 ;
			RECT	60.833 23.468 60.865 23.532 ;
			RECT	61.001 23.468 61.033 23.532 ;
			RECT	61.169 23.468 61.201 23.532 ;
			RECT	61.337 23.468 61.369 23.532 ;
			RECT	61.505 23.468 61.537 23.532 ;
			RECT	61.673 23.468 61.705 23.532 ;
			RECT	61.841 23.468 61.873 23.532 ;
			RECT	62.009 23.468 62.041 23.532 ;
			RECT	62.177 23.468 62.209 23.532 ;
			RECT	62.345 23.468 62.377 23.532 ;
			RECT	62.513 23.468 62.545 23.532 ;
			RECT	62.681 23.468 62.713 23.532 ;
			RECT	62.849 23.468 62.881 23.532 ;
			RECT	63.017 23.468 63.049 23.532 ;
			RECT	63.185 23.468 63.217 23.532 ;
			RECT	63.353 23.468 63.385 23.532 ;
			RECT	63.521 23.468 63.553 23.532 ;
			RECT	63.689 23.468 63.721 23.532 ;
			RECT	63.857 23.468 63.889 23.532 ;
			RECT	64.025 23.468 64.057 23.532 ;
			RECT	64.193 23.468 64.225 23.532 ;
			RECT	64.361 23.468 64.393 23.532 ;
			RECT	64.529 23.468 64.561 23.532 ;
			RECT	64.697 23.468 64.729 23.532 ;
			RECT	64.865 23.468 64.897 23.532 ;
			RECT	65.033 23.468 65.065 23.532 ;
			RECT	65.201 23.468 65.233 23.532 ;
			RECT	65.369 23.468 65.401 23.532 ;
			RECT	65.537 23.468 65.569 23.532 ;
			RECT	65.705 23.468 65.737 23.532 ;
			RECT	65.873 23.468 65.905 23.532 ;
			RECT	66.041 23.468 66.073 23.532 ;
			RECT	66.209 23.468 66.241 23.532 ;
			RECT	66.377 23.468 66.409 23.532 ;
			RECT	66.545 23.468 66.577 23.532 ;
			RECT	66.713 23.468 66.745 23.532 ;
			RECT	66.881 23.468 66.913 23.532 ;
			RECT	67.049 23.468 67.081 23.532 ;
			RECT	67.217 23.468 67.249 23.532 ;
			RECT	67.385 23.468 67.417 23.532 ;
			RECT	67.553 23.468 67.585 23.532 ;
			RECT	67.721 23.468 67.753 23.532 ;
			RECT	67.889 23.468 67.921 23.532 ;
			RECT	68.057 23.468 68.089 23.532 ;
			RECT	68.225 23.468 68.257 23.532 ;
			RECT	68.393 23.468 68.425 23.532 ;
			RECT	68.561 23.468 68.593 23.532 ;
			RECT	68.729 23.468 68.761 23.532 ;
			RECT	68.897 23.468 68.929 23.532 ;
			RECT	69.065 23.468 69.097 23.532 ;
			RECT	69.233 23.468 69.265 23.532 ;
			RECT	69.401 23.468 69.433 23.532 ;
			RECT	69.569 23.468 69.601 23.532 ;
			RECT	69.737 23.468 69.769 23.532 ;
			RECT	69.905 23.468 69.937 23.532 ;
			RECT	70.073 23.468 70.105 23.532 ;
			RECT	70.241 23.468 70.273 23.532 ;
			RECT	70.409 23.468 70.441 23.532 ;
			RECT	70.577 23.468 70.609 23.532 ;
			RECT	70.745 23.468 70.777 23.532 ;
			RECT	70.913 23.468 70.945 23.532 ;
			RECT	71.081 23.468 71.113 23.532 ;
			RECT	71.249 23.468 71.281 23.532 ;
			RECT	71.417 23.468 71.449 23.532 ;
			RECT	71.585 23.468 71.617 23.532 ;
			RECT	71.753 23.468 71.785 23.532 ;
			RECT	71.921 23.468 71.953 23.532 ;
			RECT	72.089 23.468 72.121 23.532 ;
			RECT	72.257 23.468 72.289 23.532 ;
			RECT	72.425 23.468 72.457 23.532 ;
			RECT	72.593 23.468 72.625 23.532 ;
			RECT	72.761 23.468 72.793 23.532 ;
			RECT	72.929 23.468 72.961 23.532 ;
			RECT	73.097 23.468 73.129 23.532 ;
			RECT	73.265 23.468 73.297 23.532 ;
			RECT	73.433 23.468 73.465 23.532 ;
			RECT	73.601 23.468 73.633 23.532 ;
			RECT	73.769 23.468 73.801 23.532 ;
			RECT	73.937 23.468 73.969 23.532 ;
			RECT	74.105 23.468 74.137 23.532 ;
			RECT	74.273 23.468 74.305 23.532 ;
			RECT	74.441 23.468 74.473 23.532 ;
			RECT	74.609 23.468 74.641 23.532 ;
			RECT	74.777 23.468 74.809 23.532 ;
			RECT	74.945 23.468 74.977 23.532 ;
			RECT	75.113 23.468 75.145 23.532 ;
			RECT	75.281 23.468 75.313 23.532 ;
			RECT	75.449 23.468 75.481 23.532 ;
			RECT	75.617 23.468 75.649 23.532 ;
			RECT	75.785 23.468 75.817 23.532 ;
			RECT	75.953 23.468 75.985 23.532 ;
			RECT	76.121 23.468 76.153 23.532 ;
			RECT	76.289 23.468 76.321 23.532 ;
			RECT	76.457 23.468 76.489 23.532 ;
			RECT	76.625 23.468 76.657 23.532 ;
			RECT	76.793 23.468 76.825 23.532 ;
			RECT	76.961 23.468 76.993 23.532 ;
			RECT	77.129 23.468 77.161 23.532 ;
			RECT	77.297 23.468 77.329 23.532 ;
			RECT	77.465 23.468 77.497 23.532 ;
			RECT	77.633 23.468 77.665 23.532 ;
			RECT	77.801 23.468 77.833 23.532 ;
			RECT	77.969 23.468 78.001 23.532 ;
			RECT	78.137 23.468 78.169 23.532 ;
			RECT	78.305 23.468 78.337 23.532 ;
			RECT	78.473 23.468 78.505 23.532 ;
			RECT	78.641 23.468 78.673 23.532 ;
			RECT	78.809 23.468 78.841 23.532 ;
			RECT	78.977 23.468 79.009 23.532 ;
			RECT	79.145 23.468 79.177 23.532 ;
			RECT	79.313 23.468 79.345 23.532 ;
			RECT	79.481 23.468 79.513 23.532 ;
			RECT	79.649 23.468 79.681 23.532 ;
			RECT	79.817 23.468 79.849 23.532 ;
			RECT	79.985 23.468 80.017 23.532 ;
			RECT	80.153 23.468 80.185 23.532 ;
			RECT	80.321 23.468 80.353 23.532 ;
			RECT	80.489 23.468 80.521 23.532 ;
			RECT	80.657 23.468 80.689 23.532 ;
			RECT	80.825 23.468 80.857 23.532 ;
			RECT	80.993 23.468 81.025 23.532 ;
			RECT	81.161 23.468 81.193 23.532 ;
			RECT	81.329 23.468 81.361 23.532 ;
			RECT	81.497 23.468 81.529 23.532 ;
			RECT	81.665 23.468 81.697 23.532 ;
			RECT	81.833 23.468 81.865 23.532 ;
			RECT	82.001 23.468 82.033 23.532 ;
			RECT	82.169 23.468 82.201 23.532 ;
			RECT	82.337 23.468 82.369 23.532 ;
			RECT	82.505 23.468 82.537 23.532 ;
			RECT	82.673 23.468 82.705 23.532 ;
			RECT	82.841 23.468 82.873 23.532 ;
			RECT	83.009 23.468 83.041 23.532 ;
			RECT	83.177 23.468 83.209 23.532 ;
			RECT	83.345 23.468 83.377 23.532 ;
			RECT	83.513 23.468 83.545 23.532 ;
			RECT	83.681 23.468 83.713 23.532 ;
			RECT	83.849 23.468 83.881 23.532 ;
			RECT	84.017 23.468 84.049 23.532 ;
			RECT	84.185 23.468 84.217 23.532 ;
			RECT	84.353 23.468 84.385 23.532 ;
			RECT	84.521 23.468 84.553 23.532 ;
			RECT	84.689 23.468 84.721 23.532 ;
			RECT	84.857 23.468 84.889 23.532 ;
			RECT	85.025 23.468 85.057 23.532 ;
			RECT	85.193 23.468 85.225 23.532 ;
			RECT	85.361 23.468 85.393 23.532 ;
			RECT	85.529 23.468 85.561 23.532 ;
			RECT	85.697 23.468 85.729 23.532 ;
			RECT	85.865 23.468 85.897 23.532 ;
			RECT	86.033 23.468 86.065 23.532 ;
			RECT	86.201 23.468 86.233 23.532 ;
			RECT	86.369 23.468 86.401 23.532 ;
			RECT	86.537 23.468 86.569 23.532 ;
			RECT	86.705 23.468 86.737 23.532 ;
			RECT	86.873 23.468 86.905 23.532 ;
			RECT	87.041 23.468 87.073 23.532 ;
			RECT	87.209 23.468 87.241 23.532 ;
			RECT	87.377 23.468 87.409 23.532 ;
			RECT	87.545 23.468 87.577 23.532 ;
			RECT	87.713 23.468 87.745 23.532 ;
			RECT	87.881 23.468 87.913 23.532 ;
			RECT	88.049 23.468 88.081 23.532 ;
			RECT	88.217 23.468 88.249 23.532 ;
			RECT	88.385 23.468 88.417 23.532 ;
			RECT	88.553 23.468 88.585 23.532 ;
			RECT	88.721 23.468 88.753 23.532 ;
			RECT	88.889 23.468 88.921 23.532 ;
			RECT	89.057 23.468 89.089 23.532 ;
			RECT	89.225 23.468 89.257 23.532 ;
			RECT	89.393 23.468 89.425 23.532 ;
			RECT	89.561 23.468 89.593 23.532 ;
			RECT	89.729 23.468 89.761 23.532 ;
			RECT	89.897 23.468 89.929 23.532 ;
			RECT	90.065 23.468 90.097 23.532 ;
			RECT	90.233 23.468 90.265 23.532 ;
			RECT	90.401 23.468 90.433 23.532 ;
			RECT	90.569 23.468 90.601 23.532 ;
			RECT	90.737 23.468 90.769 23.532 ;
			RECT	90.905 23.468 90.937 23.532 ;
			RECT	91.073 23.468 91.105 23.532 ;
			RECT	91.241 23.468 91.273 23.532 ;
			RECT	91.409 23.468 91.441 23.532 ;
			RECT	91.577 23.468 91.609 23.532 ;
			RECT	91.745 23.468 91.777 23.532 ;
			RECT	91.913 23.468 91.945 23.532 ;
			RECT	92.081 23.468 92.113 23.532 ;
			RECT	92.249 23.468 92.281 23.532 ;
			RECT	92.417 23.468 92.449 23.532 ;
			RECT	92.585 23.468 92.617 23.532 ;
			RECT	92.753 23.468 92.785 23.532 ;
			RECT	92.921 23.468 92.953 23.532 ;
			RECT	93.089 23.468 93.121 23.532 ;
			RECT	93.257 23.468 93.289 23.532 ;
			RECT	93.425 23.468 93.457 23.532 ;
			RECT	93.593 23.468 93.625 23.532 ;
			RECT	93.761 23.468 93.793 23.532 ;
			RECT	93.929 23.468 93.961 23.532 ;
			RECT	94.097 23.468 94.129 23.532 ;
			RECT	94.265 23.468 94.297 23.532 ;
			RECT	94.433 23.468 94.465 23.532 ;
			RECT	94.601 23.468 94.633 23.532 ;
			RECT	94.769 23.468 94.801 23.532 ;
			RECT	94.937 23.468 94.969 23.532 ;
			RECT	95.105 23.468 95.137 23.532 ;
			RECT	95.273 23.468 95.305 23.532 ;
			RECT	95.441 23.468 95.473 23.532 ;
			RECT	95.609 23.468 95.641 23.532 ;
			RECT	95.777 23.468 95.809 23.532 ;
			RECT	95.945 23.468 95.977 23.532 ;
			RECT	96.113 23.468 96.145 23.532 ;
			RECT	96.281 23.468 96.313 23.532 ;
			RECT	96.449 23.468 96.481 23.532 ;
			RECT	96.617 23.468 96.649 23.532 ;
			RECT	96.785 23.468 96.817 23.532 ;
			RECT	96.953 23.468 96.985 23.532 ;
			RECT	97.121 23.468 97.153 23.532 ;
			RECT	97.289 23.468 97.321 23.532 ;
			RECT	97.457 23.468 97.489 23.532 ;
			RECT	97.625 23.468 97.657 23.532 ;
			RECT	97.793 23.468 97.825 23.532 ;
			RECT	97.961 23.468 97.993 23.532 ;
			RECT	98.129 23.468 98.161 23.532 ;
			RECT	98.297 23.468 98.329 23.532 ;
			RECT	98.465 23.468 98.497 23.532 ;
			RECT	98.633 23.468 98.665 23.532 ;
			RECT	98.801 23.468 98.833 23.532 ;
			RECT	98.969 23.468 99.001 23.532 ;
			RECT	99.137 23.468 99.169 23.532 ;
			RECT	99.305 23.468 99.337 23.532 ;
			RECT	99.473 23.468 99.505 23.532 ;
			RECT	99.641 23.468 99.673 23.532 ;
			RECT	99.809 23.468 99.841 23.532 ;
			RECT	99.977 23.468 100.009 23.532 ;
			RECT	100.145 23.468 100.177 23.532 ;
			RECT	100.313 23.468 100.345 23.532 ;
			RECT	100.481 23.468 100.513 23.532 ;
			RECT	100.649 23.468 100.681 23.532 ;
			RECT	100.817 23.468 100.849 23.532 ;
			RECT	100.985 23.468 101.017 23.532 ;
			RECT	101.153 23.468 101.185 23.532 ;
			RECT	101.321 23.468 101.353 23.532 ;
			RECT	101.489 23.468 101.521 23.532 ;
			RECT	101.657 23.468 101.689 23.532 ;
			RECT	101.825 23.468 101.857 23.532 ;
			RECT	101.993 23.468 102.025 23.532 ;
			RECT	102.123 23.484 102.155 23.516 ;
			RECT	102.245 23.489 102.277 23.521 ;
			RECT	102.375 23.468 102.407 23.532 ;
			RECT	103.795 23.468 103.827 23.532 ;
			RECT	103.925 23.489 103.957 23.521 ;
			RECT	104.047 23.484 104.079 23.516 ;
			RECT	104.177 23.468 104.209 23.532 ;
			RECT	104.345 23.468 104.377 23.532 ;
			RECT	104.513 23.468 104.545 23.532 ;
			RECT	104.681 23.468 104.713 23.532 ;
			RECT	104.849 23.468 104.881 23.532 ;
			RECT	105.017 23.468 105.049 23.532 ;
			RECT	105.185 23.468 105.217 23.532 ;
			RECT	105.353 23.468 105.385 23.532 ;
			RECT	105.521 23.468 105.553 23.532 ;
			RECT	105.689 23.468 105.721 23.532 ;
			RECT	105.857 23.468 105.889 23.532 ;
			RECT	106.025 23.468 106.057 23.532 ;
			RECT	106.193 23.468 106.225 23.532 ;
			RECT	106.361 23.468 106.393 23.532 ;
			RECT	106.529 23.468 106.561 23.532 ;
			RECT	106.697 23.468 106.729 23.532 ;
			RECT	106.865 23.468 106.897 23.532 ;
			RECT	107.033 23.468 107.065 23.532 ;
			RECT	107.201 23.468 107.233 23.532 ;
			RECT	107.369 23.468 107.401 23.532 ;
			RECT	107.537 23.468 107.569 23.532 ;
			RECT	107.705 23.468 107.737 23.532 ;
			RECT	107.873 23.468 107.905 23.532 ;
			RECT	108.041 23.468 108.073 23.532 ;
			RECT	108.209 23.468 108.241 23.532 ;
			RECT	108.377 23.468 108.409 23.532 ;
			RECT	108.545 23.468 108.577 23.532 ;
			RECT	108.713 23.468 108.745 23.532 ;
			RECT	108.881 23.468 108.913 23.532 ;
			RECT	109.049 23.468 109.081 23.532 ;
			RECT	109.217 23.468 109.249 23.532 ;
			RECT	109.385 23.468 109.417 23.532 ;
			RECT	109.553 23.468 109.585 23.532 ;
			RECT	109.721 23.468 109.753 23.532 ;
			RECT	109.889 23.468 109.921 23.532 ;
			RECT	110.057 23.468 110.089 23.532 ;
			RECT	110.225 23.468 110.257 23.532 ;
			RECT	110.393 23.468 110.425 23.532 ;
			RECT	110.561 23.468 110.593 23.532 ;
			RECT	110.729 23.468 110.761 23.532 ;
			RECT	110.897 23.468 110.929 23.532 ;
			RECT	111.065 23.468 111.097 23.532 ;
			RECT	111.233 23.468 111.265 23.532 ;
			RECT	111.401 23.468 111.433 23.532 ;
			RECT	111.569 23.468 111.601 23.532 ;
			RECT	111.737 23.468 111.769 23.532 ;
			RECT	111.905 23.468 111.937 23.532 ;
			RECT	112.073 23.468 112.105 23.532 ;
			RECT	112.241 23.468 112.273 23.532 ;
			RECT	112.409 23.468 112.441 23.532 ;
			RECT	112.577 23.468 112.609 23.532 ;
			RECT	112.745 23.468 112.777 23.532 ;
			RECT	112.913 23.468 112.945 23.532 ;
			RECT	113.081 23.468 113.113 23.532 ;
			RECT	113.249 23.468 113.281 23.532 ;
			RECT	113.417 23.468 113.449 23.532 ;
			RECT	113.585 23.468 113.617 23.532 ;
			RECT	113.753 23.468 113.785 23.532 ;
			RECT	113.921 23.468 113.953 23.532 ;
			RECT	114.089 23.468 114.121 23.532 ;
			RECT	114.257 23.468 114.289 23.532 ;
			RECT	114.425 23.468 114.457 23.532 ;
			RECT	114.593 23.468 114.625 23.532 ;
			RECT	114.761 23.468 114.793 23.532 ;
			RECT	114.929 23.468 114.961 23.532 ;
			RECT	115.097 23.468 115.129 23.532 ;
			RECT	115.265 23.468 115.297 23.532 ;
			RECT	115.433 23.468 115.465 23.532 ;
			RECT	115.601 23.468 115.633 23.532 ;
			RECT	115.769 23.468 115.801 23.532 ;
			RECT	115.937 23.468 115.969 23.532 ;
			RECT	116.105 23.468 116.137 23.532 ;
			RECT	116.273 23.468 116.305 23.532 ;
			RECT	116.441 23.468 116.473 23.532 ;
			RECT	116.609 23.468 116.641 23.532 ;
			RECT	116.777 23.468 116.809 23.532 ;
			RECT	116.945 23.468 116.977 23.532 ;
			RECT	117.113 23.468 117.145 23.532 ;
			RECT	117.281 23.468 117.313 23.532 ;
			RECT	117.449 23.468 117.481 23.532 ;
			RECT	117.617 23.468 117.649 23.532 ;
			RECT	117.785 23.468 117.817 23.532 ;
			RECT	117.953 23.468 117.985 23.532 ;
			RECT	118.121 23.468 118.153 23.532 ;
			RECT	118.289 23.468 118.321 23.532 ;
			RECT	118.457 23.468 118.489 23.532 ;
			RECT	118.625 23.468 118.657 23.532 ;
			RECT	118.793 23.468 118.825 23.532 ;
			RECT	118.961 23.468 118.993 23.532 ;
			RECT	119.129 23.468 119.161 23.532 ;
			RECT	119.297 23.468 119.329 23.532 ;
			RECT	119.465 23.468 119.497 23.532 ;
			RECT	119.633 23.468 119.665 23.532 ;
			RECT	119.801 23.468 119.833 23.532 ;
			RECT	119.969 23.468 120.001 23.532 ;
			RECT	120.137 23.468 120.169 23.532 ;
			RECT	120.305 23.468 120.337 23.532 ;
			RECT	120.473 23.468 120.505 23.532 ;
			RECT	120.641 23.468 120.673 23.532 ;
			RECT	120.809 23.468 120.841 23.532 ;
			RECT	120.977 23.468 121.009 23.532 ;
			RECT	121.145 23.468 121.177 23.532 ;
			RECT	121.313 23.468 121.345 23.532 ;
			RECT	121.481 23.468 121.513 23.532 ;
			RECT	121.649 23.468 121.681 23.532 ;
			RECT	121.817 23.468 121.849 23.532 ;
			RECT	121.985 23.468 122.017 23.532 ;
			RECT	122.153 23.468 122.185 23.532 ;
			RECT	122.321 23.468 122.353 23.532 ;
			RECT	122.489 23.468 122.521 23.532 ;
			RECT	122.657 23.468 122.689 23.532 ;
			RECT	122.825 23.468 122.857 23.532 ;
			RECT	122.993 23.468 123.025 23.532 ;
			RECT	123.161 23.468 123.193 23.532 ;
			RECT	123.329 23.468 123.361 23.532 ;
			RECT	123.497 23.468 123.529 23.532 ;
			RECT	123.665 23.468 123.697 23.532 ;
			RECT	123.833 23.468 123.865 23.532 ;
			RECT	124.001 23.468 124.033 23.532 ;
			RECT	124.169 23.468 124.201 23.532 ;
			RECT	124.337 23.468 124.369 23.532 ;
			RECT	124.505 23.468 124.537 23.532 ;
			RECT	124.673 23.468 124.705 23.532 ;
			RECT	124.841 23.468 124.873 23.532 ;
			RECT	125.009 23.468 125.041 23.532 ;
			RECT	125.177 23.468 125.209 23.532 ;
			RECT	125.345 23.468 125.377 23.532 ;
			RECT	125.513 23.468 125.545 23.532 ;
			RECT	125.681 23.468 125.713 23.532 ;
			RECT	125.849 23.468 125.881 23.532 ;
			RECT	126.017 23.468 126.049 23.532 ;
			RECT	126.185 23.468 126.217 23.532 ;
			RECT	126.353 23.468 126.385 23.532 ;
			RECT	126.521 23.468 126.553 23.532 ;
			RECT	126.689 23.468 126.721 23.532 ;
			RECT	126.857 23.468 126.889 23.532 ;
			RECT	127.025 23.468 127.057 23.532 ;
			RECT	127.193 23.468 127.225 23.532 ;
			RECT	127.361 23.468 127.393 23.532 ;
			RECT	127.529 23.468 127.561 23.532 ;
			RECT	127.697 23.468 127.729 23.532 ;
			RECT	127.865 23.468 127.897 23.532 ;
			RECT	128.033 23.468 128.065 23.532 ;
			RECT	128.201 23.468 128.233 23.532 ;
			RECT	128.369 23.468 128.401 23.532 ;
			RECT	128.537 23.468 128.569 23.532 ;
			RECT	128.705 23.468 128.737 23.532 ;
			RECT	128.873 23.468 128.905 23.532 ;
			RECT	129.041 23.468 129.073 23.532 ;
			RECT	129.209 23.468 129.241 23.532 ;
			RECT	129.377 23.468 129.409 23.532 ;
			RECT	129.545 23.468 129.577 23.532 ;
			RECT	129.713 23.468 129.745 23.532 ;
			RECT	129.881 23.468 129.913 23.532 ;
			RECT	130.049 23.468 130.081 23.532 ;
			RECT	130.217 23.468 130.249 23.532 ;
			RECT	130.385 23.468 130.417 23.532 ;
			RECT	130.553 23.468 130.585 23.532 ;
			RECT	130.721 23.468 130.753 23.532 ;
			RECT	130.889 23.468 130.921 23.532 ;
			RECT	131.057 23.468 131.089 23.532 ;
			RECT	131.225 23.468 131.257 23.532 ;
			RECT	131.393 23.468 131.425 23.532 ;
			RECT	131.561 23.468 131.593 23.532 ;
			RECT	131.729 23.468 131.761 23.532 ;
			RECT	131.897 23.468 131.929 23.532 ;
			RECT	132.065 23.468 132.097 23.532 ;
			RECT	132.233 23.468 132.265 23.532 ;
			RECT	132.401 23.468 132.433 23.532 ;
			RECT	132.569 23.468 132.601 23.532 ;
			RECT	132.737 23.468 132.769 23.532 ;
			RECT	132.905 23.468 132.937 23.532 ;
			RECT	133.073 23.468 133.105 23.532 ;
			RECT	133.241 23.468 133.273 23.532 ;
			RECT	133.409 23.468 133.441 23.532 ;
			RECT	133.577 23.468 133.609 23.532 ;
			RECT	133.745 23.468 133.777 23.532 ;
			RECT	133.913 23.468 133.945 23.532 ;
			RECT	134.081 23.468 134.113 23.532 ;
			RECT	134.249 23.468 134.281 23.532 ;
			RECT	134.417 23.468 134.449 23.532 ;
			RECT	134.585 23.468 134.617 23.532 ;
			RECT	134.753 23.468 134.785 23.532 ;
			RECT	134.921 23.468 134.953 23.532 ;
			RECT	135.089 23.468 135.121 23.532 ;
			RECT	135.257 23.468 135.289 23.532 ;
			RECT	135.425 23.468 135.457 23.532 ;
			RECT	135.593 23.468 135.625 23.532 ;
			RECT	135.761 23.468 135.793 23.532 ;
			RECT	135.929 23.468 135.961 23.532 ;
			RECT	136.097 23.468 136.129 23.532 ;
			RECT	136.265 23.468 136.297 23.532 ;
			RECT	136.433 23.468 136.465 23.532 ;
			RECT	136.601 23.468 136.633 23.532 ;
			RECT	136.769 23.468 136.801 23.532 ;
			RECT	136.937 23.468 136.969 23.532 ;
			RECT	137.105 23.468 137.137 23.532 ;
			RECT	137.273 23.468 137.305 23.532 ;
			RECT	137.441 23.468 137.473 23.532 ;
			RECT	137.609 23.468 137.641 23.532 ;
			RECT	137.777 23.468 137.809 23.532 ;
			RECT	137.945 23.468 137.977 23.532 ;
			RECT	138.113 23.468 138.145 23.532 ;
			RECT	138.281 23.468 138.313 23.532 ;
			RECT	138.449 23.468 138.481 23.532 ;
			RECT	138.617 23.468 138.649 23.532 ;
			RECT	138.785 23.468 138.817 23.532 ;
			RECT	138.953 23.468 138.985 23.532 ;
			RECT	139.121 23.468 139.153 23.532 ;
			RECT	139.289 23.468 139.321 23.532 ;
			RECT	139.457 23.468 139.489 23.532 ;
			RECT	139.625 23.468 139.657 23.532 ;
			RECT	139.793 23.468 139.825 23.532 ;
			RECT	139.961 23.468 139.993 23.532 ;
			RECT	140.129 23.468 140.161 23.532 ;
			RECT	140.297 23.468 140.329 23.532 ;
			RECT	140.465 23.468 140.497 23.532 ;
			RECT	140.633 23.468 140.665 23.532 ;
			RECT	140.801 23.468 140.833 23.532 ;
			RECT	140.969 23.468 141.001 23.532 ;
			RECT	141.137 23.468 141.169 23.532 ;
			RECT	141.305 23.468 141.337 23.532 ;
			RECT	141.473 23.468 141.505 23.532 ;
			RECT	141.641 23.468 141.673 23.532 ;
			RECT	141.809 23.468 141.841 23.532 ;
			RECT	141.977 23.468 142.009 23.532 ;
			RECT	142.145 23.468 142.177 23.532 ;
			RECT	142.313 23.468 142.345 23.532 ;
			RECT	142.481 23.468 142.513 23.532 ;
			RECT	142.649 23.468 142.681 23.532 ;
			RECT	142.817 23.468 142.849 23.532 ;
			RECT	142.985 23.468 143.017 23.532 ;
			RECT	143.153 23.468 143.185 23.532 ;
			RECT	143.321 23.468 143.353 23.532 ;
			RECT	143.489 23.468 143.521 23.532 ;
			RECT	143.657 23.468 143.689 23.532 ;
			RECT	143.825 23.468 143.857 23.532 ;
			RECT	143.993 23.468 144.025 23.532 ;
			RECT	144.161 23.468 144.193 23.532 ;
			RECT	144.329 23.468 144.361 23.532 ;
			RECT	144.497 23.468 144.529 23.532 ;
			RECT	144.665 23.468 144.697 23.532 ;
			RECT	144.833 23.468 144.865 23.532 ;
			RECT	145.001 23.468 145.033 23.532 ;
			RECT	145.169 23.468 145.201 23.532 ;
			RECT	145.337 23.468 145.369 23.532 ;
			RECT	145.505 23.468 145.537 23.532 ;
			RECT	145.673 23.468 145.705 23.532 ;
			RECT	145.841 23.468 145.873 23.532 ;
			RECT	146.009 23.468 146.041 23.532 ;
			RECT	146.177 23.468 146.209 23.532 ;
			RECT	146.345 23.468 146.377 23.532 ;
			RECT	146.513 23.468 146.545 23.532 ;
			RECT	146.681 23.468 146.713 23.532 ;
			RECT	146.849 23.468 146.881 23.532 ;
			RECT	147.017 23.468 147.049 23.532 ;
			RECT	147.185 23.468 147.217 23.532 ;
			RECT	147.316 23.484 147.348 23.516 ;
			RECT	147.437 23.484 147.469 23.516 ;
			RECT	147.567 23.468 147.599 23.532 ;
			RECT	149.879 23.468 149.911 23.532 ;
			RECT	151.13 23.468 151.194 23.532 ;
			RECT	151.81 23.468 151.842 23.532 ;
			RECT	152.249 23.468 152.281 23.532 ;
			RECT	153.56 23.468 153.624 23.532 ;
			RECT	156.601 23.468 156.633 23.532 ;
			RECT	156.731 23.484 156.763 23.516 ;
			RECT	156.852 23.484 156.884 23.516 ;
			RECT	156.983 23.468 157.015 23.532 ;
			RECT	157.151 23.468 157.183 23.532 ;
			RECT	157.319 23.468 157.351 23.532 ;
			RECT	157.487 23.468 157.519 23.532 ;
			RECT	157.655 23.468 157.687 23.532 ;
			RECT	157.823 23.468 157.855 23.532 ;
			RECT	157.991 23.468 158.023 23.532 ;
			RECT	158.159 23.468 158.191 23.532 ;
			RECT	158.327 23.468 158.359 23.532 ;
			RECT	158.495 23.468 158.527 23.532 ;
			RECT	158.663 23.468 158.695 23.532 ;
			RECT	158.831 23.468 158.863 23.532 ;
			RECT	158.999 23.468 159.031 23.532 ;
			RECT	159.167 23.468 159.199 23.532 ;
			RECT	159.335 23.468 159.367 23.532 ;
			RECT	159.503 23.468 159.535 23.532 ;
			RECT	159.671 23.468 159.703 23.532 ;
			RECT	159.839 23.468 159.871 23.532 ;
			RECT	160.007 23.468 160.039 23.532 ;
			RECT	160.175 23.468 160.207 23.532 ;
			RECT	160.343 23.468 160.375 23.532 ;
			RECT	160.511 23.468 160.543 23.532 ;
			RECT	160.679 23.468 160.711 23.532 ;
			RECT	160.847 23.468 160.879 23.532 ;
			RECT	161.015 23.468 161.047 23.532 ;
			RECT	161.183 23.468 161.215 23.532 ;
			RECT	161.351 23.468 161.383 23.532 ;
			RECT	161.519 23.468 161.551 23.532 ;
			RECT	161.687 23.468 161.719 23.532 ;
			RECT	161.855 23.468 161.887 23.532 ;
			RECT	162.023 23.468 162.055 23.532 ;
			RECT	162.191 23.468 162.223 23.532 ;
			RECT	162.359 23.468 162.391 23.532 ;
			RECT	162.527 23.468 162.559 23.532 ;
			RECT	162.695 23.468 162.727 23.532 ;
			RECT	162.863 23.468 162.895 23.532 ;
			RECT	163.031 23.468 163.063 23.532 ;
			RECT	163.199 23.468 163.231 23.532 ;
			RECT	163.367 23.468 163.399 23.532 ;
			RECT	163.535 23.468 163.567 23.532 ;
			RECT	163.703 23.468 163.735 23.532 ;
			RECT	163.871 23.468 163.903 23.532 ;
			RECT	164.039 23.468 164.071 23.532 ;
			RECT	164.207 23.468 164.239 23.532 ;
			RECT	164.375 23.468 164.407 23.532 ;
			RECT	164.543 23.468 164.575 23.532 ;
			RECT	164.711 23.468 164.743 23.532 ;
			RECT	164.879 23.468 164.911 23.532 ;
			RECT	165.047 23.468 165.079 23.532 ;
			RECT	165.215 23.468 165.247 23.532 ;
			RECT	165.383 23.468 165.415 23.532 ;
			RECT	165.551 23.468 165.583 23.532 ;
			RECT	165.719 23.468 165.751 23.532 ;
			RECT	165.887 23.468 165.919 23.532 ;
			RECT	166.055 23.468 166.087 23.532 ;
			RECT	166.223 23.468 166.255 23.532 ;
			RECT	166.391 23.468 166.423 23.532 ;
			RECT	166.559 23.468 166.591 23.532 ;
			RECT	166.727 23.468 166.759 23.532 ;
			RECT	166.895 23.468 166.927 23.532 ;
			RECT	167.063 23.468 167.095 23.532 ;
			RECT	167.231 23.468 167.263 23.532 ;
			RECT	167.399 23.468 167.431 23.532 ;
			RECT	167.567 23.468 167.599 23.532 ;
			RECT	167.735 23.468 167.767 23.532 ;
			RECT	167.903 23.468 167.935 23.532 ;
			RECT	168.071 23.468 168.103 23.532 ;
			RECT	168.239 23.468 168.271 23.532 ;
			RECT	168.407 23.468 168.439 23.532 ;
			RECT	168.575 23.468 168.607 23.532 ;
			RECT	168.743 23.468 168.775 23.532 ;
			RECT	168.911 23.468 168.943 23.532 ;
			RECT	169.079 23.468 169.111 23.532 ;
			RECT	169.247 23.468 169.279 23.532 ;
			RECT	169.415 23.468 169.447 23.532 ;
			RECT	169.583 23.468 169.615 23.532 ;
			RECT	169.751 23.468 169.783 23.532 ;
			RECT	169.919 23.468 169.951 23.532 ;
			RECT	170.087 23.468 170.119 23.532 ;
			RECT	170.255 23.468 170.287 23.532 ;
			RECT	170.423 23.468 170.455 23.532 ;
			RECT	170.591 23.468 170.623 23.532 ;
			RECT	170.759 23.468 170.791 23.532 ;
			RECT	170.927 23.468 170.959 23.532 ;
			RECT	171.095 23.468 171.127 23.532 ;
			RECT	171.263 23.468 171.295 23.532 ;
			RECT	171.431 23.468 171.463 23.532 ;
			RECT	171.599 23.468 171.631 23.532 ;
			RECT	171.767 23.468 171.799 23.532 ;
			RECT	171.935 23.468 171.967 23.532 ;
			RECT	172.103 23.468 172.135 23.532 ;
			RECT	172.271 23.468 172.303 23.532 ;
			RECT	172.439 23.468 172.471 23.532 ;
			RECT	172.607 23.468 172.639 23.532 ;
			RECT	172.775 23.468 172.807 23.532 ;
			RECT	172.943 23.468 172.975 23.532 ;
			RECT	173.111 23.468 173.143 23.532 ;
			RECT	173.279 23.468 173.311 23.532 ;
			RECT	173.447 23.468 173.479 23.532 ;
			RECT	173.615 23.468 173.647 23.532 ;
			RECT	173.783 23.468 173.815 23.532 ;
			RECT	173.951 23.468 173.983 23.532 ;
			RECT	174.119 23.468 174.151 23.532 ;
			RECT	174.287 23.468 174.319 23.532 ;
			RECT	174.455 23.468 174.487 23.532 ;
			RECT	174.623 23.468 174.655 23.532 ;
			RECT	174.791 23.468 174.823 23.532 ;
			RECT	174.959 23.468 174.991 23.532 ;
			RECT	175.127 23.468 175.159 23.532 ;
			RECT	175.295 23.468 175.327 23.532 ;
			RECT	175.463 23.468 175.495 23.532 ;
			RECT	175.631 23.468 175.663 23.532 ;
			RECT	175.799 23.468 175.831 23.532 ;
			RECT	175.967 23.468 175.999 23.532 ;
			RECT	176.135 23.468 176.167 23.532 ;
			RECT	176.303 23.468 176.335 23.532 ;
			RECT	176.471 23.468 176.503 23.532 ;
			RECT	176.639 23.468 176.671 23.532 ;
			RECT	176.807 23.468 176.839 23.532 ;
			RECT	176.975 23.468 177.007 23.532 ;
			RECT	177.143 23.468 177.175 23.532 ;
			RECT	177.311 23.468 177.343 23.532 ;
			RECT	177.479 23.468 177.511 23.532 ;
			RECT	177.647 23.468 177.679 23.532 ;
			RECT	177.815 23.468 177.847 23.532 ;
			RECT	177.983 23.468 178.015 23.532 ;
			RECT	178.151 23.468 178.183 23.532 ;
			RECT	178.319 23.468 178.351 23.532 ;
			RECT	178.487 23.468 178.519 23.532 ;
			RECT	178.655 23.468 178.687 23.532 ;
			RECT	178.823 23.468 178.855 23.532 ;
			RECT	178.991 23.468 179.023 23.532 ;
			RECT	179.159 23.468 179.191 23.532 ;
			RECT	179.327 23.468 179.359 23.532 ;
			RECT	179.495 23.468 179.527 23.532 ;
			RECT	179.663 23.468 179.695 23.532 ;
			RECT	179.831 23.468 179.863 23.532 ;
			RECT	179.999 23.468 180.031 23.532 ;
			RECT	180.167 23.468 180.199 23.532 ;
			RECT	180.335 23.468 180.367 23.532 ;
			RECT	180.503 23.468 180.535 23.532 ;
			RECT	180.671 23.468 180.703 23.532 ;
			RECT	180.839 23.468 180.871 23.532 ;
			RECT	181.007 23.468 181.039 23.532 ;
			RECT	181.175 23.468 181.207 23.532 ;
			RECT	181.343 23.468 181.375 23.532 ;
			RECT	181.511 23.468 181.543 23.532 ;
			RECT	181.679 23.468 181.711 23.532 ;
			RECT	181.847 23.468 181.879 23.532 ;
			RECT	182.015 23.468 182.047 23.532 ;
			RECT	182.183 23.468 182.215 23.532 ;
			RECT	182.351 23.468 182.383 23.532 ;
			RECT	182.519 23.468 182.551 23.532 ;
			RECT	182.687 23.468 182.719 23.532 ;
			RECT	182.855 23.468 182.887 23.532 ;
			RECT	183.023 23.468 183.055 23.532 ;
			RECT	183.191 23.468 183.223 23.532 ;
			RECT	183.359 23.468 183.391 23.532 ;
			RECT	183.527 23.468 183.559 23.532 ;
			RECT	183.695 23.468 183.727 23.532 ;
			RECT	183.863 23.468 183.895 23.532 ;
			RECT	184.031 23.468 184.063 23.532 ;
			RECT	184.199 23.468 184.231 23.532 ;
			RECT	184.367 23.468 184.399 23.532 ;
			RECT	184.535 23.468 184.567 23.532 ;
			RECT	184.703 23.468 184.735 23.532 ;
			RECT	184.871 23.468 184.903 23.532 ;
			RECT	185.039 23.468 185.071 23.532 ;
			RECT	185.207 23.468 185.239 23.532 ;
			RECT	185.375 23.468 185.407 23.532 ;
			RECT	185.543 23.468 185.575 23.532 ;
			RECT	185.711 23.468 185.743 23.532 ;
			RECT	185.879 23.468 185.911 23.532 ;
			RECT	186.047 23.468 186.079 23.532 ;
			RECT	186.215 23.468 186.247 23.532 ;
			RECT	186.383 23.468 186.415 23.532 ;
			RECT	186.551 23.468 186.583 23.532 ;
			RECT	186.719 23.468 186.751 23.532 ;
			RECT	186.887 23.468 186.919 23.532 ;
			RECT	187.055 23.468 187.087 23.532 ;
			RECT	187.223 23.468 187.255 23.532 ;
			RECT	187.391 23.468 187.423 23.532 ;
			RECT	187.559 23.468 187.591 23.532 ;
			RECT	187.727 23.468 187.759 23.532 ;
			RECT	187.895 23.468 187.927 23.532 ;
			RECT	188.063 23.468 188.095 23.532 ;
			RECT	188.231 23.468 188.263 23.532 ;
			RECT	188.399 23.468 188.431 23.532 ;
			RECT	188.567 23.468 188.599 23.532 ;
			RECT	188.735 23.468 188.767 23.532 ;
			RECT	188.903 23.468 188.935 23.532 ;
			RECT	189.071 23.468 189.103 23.532 ;
			RECT	189.239 23.468 189.271 23.532 ;
			RECT	189.407 23.468 189.439 23.532 ;
			RECT	189.575 23.468 189.607 23.532 ;
			RECT	189.743 23.468 189.775 23.532 ;
			RECT	189.911 23.468 189.943 23.532 ;
			RECT	190.079 23.468 190.111 23.532 ;
			RECT	190.247 23.468 190.279 23.532 ;
			RECT	190.415 23.468 190.447 23.532 ;
			RECT	190.583 23.468 190.615 23.532 ;
			RECT	190.751 23.468 190.783 23.532 ;
			RECT	190.919 23.468 190.951 23.532 ;
			RECT	191.087 23.468 191.119 23.532 ;
			RECT	191.255 23.468 191.287 23.532 ;
			RECT	191.423 23.468 191.455 23.532 ;
			RECT	191.591 23.468 191.623 23.532 ;
			RECT	191.759 23.468 191.791 23.532 ;
			RECT	191.927 23.468 191.959 23.532 ;
			RECT	192.095 23.468 192.127 23.532 ;
			RECT	192.263 23.468 192.295 23.532 ;
			RECT	192.431 23.468 192.463 23.532 ;
			RECT	192.599 23.468 192.631 23.532 ;
			RECT	192.767 23.468 192.799 23.532 ;
			RECT	192.935 23.468 192.967 23.532 ;
			RECT	193.103 23.468 193.135 23.532 ;
			RECT	193.271 23.468 193.303 23.532 ;
			RECT	193.439 23.468 193.471 23.532 ;
			RECT	193.607 23.468 193.639 23.532 ;
			RECT	193.775 23.468 193.807 23.532 ;
			RECT	193.943 23.468 193.975 23.532 ;
			RECT	194.111 23.468 194.143 23.532 ;
			RECT	194.279 23.468 194.311 23.532 ;
			RECT	194.447 23.468 194.479 23.532 ;
			RECT	194.615 23.468 194.647 23.532 ;
			RECT	194.783 23.468 194.815 23.532 ;
			RECT	194.951 23.468 194.983 23.532 ;
			RECT	195.119 23.468 195.151 23.532 ;
			RECT	195.287 23.468 195.319 23.532 ;
			RECT	195.455 23.468 195.487 23.532 ;
			RECT	195.623 23.468 195.655 23.532 ;
			RECT	195.791 23.468 195.823 23.532 ;
			RECT	195.959 23.468 195.991 23.532 ;
			RECT	196.127 23.468 196.159 23.532 ;
			RECT	196.295 23.468 196.327 23.532 ;
			RECT	196.463 23.468 196.495 23.532 ;
			RECT	196.631 23.468 196.663 23.532 ;
			RECT	196.799 23.468 196.831 23.532 ;
			RECT	196.967 23.468 196.999 23.532 ;
			RECT	197.135 23.468 197.167 23.532 ;
			RECT	197.303 23.468 197.335 23.532 ;
			RECT	197.471 23.468 197.503 23.532 ;
			RECT	197.639 23.468 197.671 23.532 ;
			RECT	197.807 23.468 197.839 23.532 ;
			RECT	197.975 23.468 198.007 23.532 ;
			RECT	198.143 23.468 198.175 23.532 ;
			RECT	198.311 23.468 198.343 23.532 ;
			RECT	198.479 23.468 198.511 23.532 ;
			RECT	198.647 23.468 198.679 23.532 ;
			RECT	198.815 23.468 198.847 23.532 ;
			RECT	198.983 23.468 199.015 23.532 ;
			RECT	199.151 23.468 199.183 23.532 ;
			RECT	199.319 23.468 199.351 23.532 ;
			RECT	199.487 23.468 199.519 23.532 ;
			RECT	199.655 23.468 199.687 23.532 ;
			RECT	199.823 23.468 199.855 23.532 ;
			RECT	199.991 23.468 200.023 23.532 ;
			RECT	200.121 23.484 200.153 23.516 ;
			RECT	200.243 23.489 200.275 23.521 ;
			RECT	200.373 23.468 200.405 23.532 ;
			RECT	200.9 23.468 200.932 23.532 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 21.52 201.665 21.64 ;
			LAYER	J3 ;
			RECT	0.755 21.548 0.787 21.612 ;
			RECT	1.645 21.548 1.709 21.612 ;
			RECT	2.323 21.548 2.387 21.612 ;
			RECT	3.438 21.548 3.47 21.612 ;
			RECT	3.585 21.548 3.617 21.612 ;
			RECT	4.195 21.548 4.227 21.612 ;
			RECT	4.72 21.548 4.752 21.612 ;
			RECT	4.944 21.548 5.008 21.612 ;
			RECT	5.267 21.548 5.299 21.612 ;
			RECT	5.797 21.548 5.829 21.612 ;
			RECT	5.927 21.569 5.959 21.601 ;
			RECT	6.049 21.564 6.081 21.596 ;
			RECT	6.179 21.548 6.211 21.612 ;
			RECT	6.347 21.548 6.379 21.612 ;
			RECT	6.515 21.548 6.547 21.612 ;
			RECT	6.683 21.548 6.715 21.612 ;
			RECT	6.851 21.548 6.883 21.612 ;
			RECT	7.019 21.548 7.051 21.612 ;
			RECT	7.187 21.548 7.219 21.612 ;
			RECT	7.355 21.548 7.387 21.612 ;
			RECT	7.523 21.548 7.555 21.612 ;
			RECT	7.691 21.548 7.723 21.612 ;
			RECT	7.859 21.548 7.891 21.612 ;
			RECT	8.027 21.548 8.059 21.612 ;
			RECT	8.195 21.548 8.227 21.612 ;
			RECT	8.363 21.548 8.395 21.612 ;
			RECT	8.531 21.548 8.563 21.612 ;
			RECT	8.699 21.548 8.731 21.612 ;
			RECT	8.867 21.548 8.899 21.612 ;
			RECT	9.035 21.548 9.067 21.612 ;
			RECT	9.203 21.548 9.235 21.612 ;
			RECT	9.371 21.548 9.403 21.612 ;
			RECT	9.539 21.548 9.571 21.612 ;
			RECT	9.707 21.548 9.739 21.612 ;
			RECT	9.875 21.548 9.907 21.612 ;
			RECT	10.043 21.548 10.075 21.612 ;
			RECT	10.211 21.548 10.243 21.612 ;
			RECT	10.379 21.548 10.411 21.612 ;
			RECT	10.547 21.548 10.579 21.612 ;
			RECT	10.715 21.548 10.747 21.612 ;
			RECT	10.883 21.548 10.915 21.612 ;
			RECT	11.051 21.548 11.083 21.612 ;
			RECT	11.219 21.548 11.251 21.612 ;
			RECT	11.387 21.548 11.419 21.612 ;
			RECT	11.555 21.548 11.587 21.612 ;
			RECT	11.723 21.548 11.755 21.612 ;
			RECT	11.891 21.548 11.923 21.612 ;
			RECT	12.059 21.548 12.091 21.612 ;
			RECT	12.227 21.548 12.259 21.612 ;
			RECT	12.395 21.548 12.427 21.612 ;
			RECT	12.563 21.548 12.595 21.612 ;
			RECT	12.731 21.548 12.763 21.612 ;
			RECT	12.899 21.548 12.931 21.612 ;
			RECT	13.067 21.548 13.099 21.612 ;
			RECT	13.235 21.548 13.267 21.612 ;
			RECT	13.403 21.548 13.435 21.612 ;
			RECT	13.571 21.548 13.603 21.612 ;
			RECT	13.739 21.548 13.771 21.612 ;
			RECT	13.907 21.548 13.939 21.612 ;
			RECT	14.075 21.548 14.107 21.612 ;
			RECT	14.243 21.548 14.275 21.612 ;
			RECT	14.411 21.548 14.443 21.612 ;
			RECT	14.579 21.548 14.611 21.612 ;
			RECT	14.747 21.548 14.779 21.612 ;
			RECT	14.915 21.548 14.947 21.612 ;
			RECT	15.083 21.548 15.115 21.612 ;
			RECT	15.251 21.548 15.283 21.612 ;
			RECT	15.419 21.548 15.451 21.612 ;
			RECT	15.587 21.548 15.619 21.612 ;
			RECT	15.755 21.548 15.787 21.612 ;
			RECT	15.923 21.548 15.955 21.612 ;
			RECT	16.091 21.548 16.123 21.612 ;
			RECT	16.259 21.548 16.291 21.612 ;
			RECT	16.427 21.548 16.459 21.612 ;
			RECT	16.595 21.548 16.627 21.612 ;
			RECT	16.763 21.548 16.795 21.612 ;
			RECT	16.931 21.548 16.963 21.612 ;
			RECT	17.099 21.548 17.131 21.612 ;
			RECT	17.267 21.548 17.299 21.612 ;
			RECT	17.435 21.548 17.467 21.612 ;
			RECT	17.603 21.548 17.635 21.612 ;
			RECT	17.771 21.548 17.803 21.612 ;
			RECT	17.939 21.548 17.971 21.612 ;
			RECT	18.107 21.548 18.139 21.612 ;
			RECT	18.275 21.548 18.307 21.612 ;
			RECT	18.443 21.548 18.475 21.612 ;
			RECT	18.611 21.548 18.643 21.612 ;
			RECT	18.779 21.548 18.811 21.612 ;
			RECT	18.947 21.548 18.979 21.612 ;
			RECT	19.115 21.548 19.147 21.612 ;
			RECT	19.283 21.548 19.315 21.612 ;
			RECT	19.451 21.548 19.483 21.612 ;
			RECT	19.619 21.548 19.651 21.612 ;
			RECT	19.787 21.548 19.819 21.612 ;
			RECT	19.955 21.548 19.987 21.612 ;
			RECT	20.123 21.548 20.155 21.612 ;
			RECT	20.291 21.548 20.323 21.612 ;
			RECT	20.459 21.548 20.491 21.612 ;
			RECT	20.627 21.548 20.659 21.612 ;
			RECT	20.795 21.548 20.827 21.612 ;
			RECT	20.963 21.548 20.995 21.612 ;
			RECT	21.131 21.548 21.163 21.612 ;
			RECT	21.299 21.548 21.331 21.612 ;
			RECT	21.467 21.548 21.499 21.612 ;
			RECT	21.635 21.548 21.667 21.612 ;
			RECT	21.803 21.548 21.835 21.612 ;
			RECT	21.971 21.548 22.003 21.612 ;
			RECT	22.139 21.548 22.171 21.612 ;
			RECT	22.307 21.548 22.339 21.612 ;
			RECT	22.475 21.548 22.507 21.612 ;
			RECT	22.643 21.548 22.675 21.612 ;
			RECT	22.811 21.548 22.843 21.612 ;
			RECT	22.979 21.548 23.011 21.612 ;
			RECT	23.147 21.548 23.179 21.612 ;
			RECT	23.315 21.548 23.347 21.612 ;
			RECT	23.483 21.548 23.515 21.612 ;
			RECT	23.651 21.548 23.683 21.612 ;
			RECT	23.819 21.548 23.851 21.612 ;
			RECT	23.987 21.548 24.019 21.612 ;
			RECT	24.155 21.548 24.187 21.612 ;
			RECT	24.323 21.548 24.355 21.612 ;
			RECT	24.491 21.548 24.523 21.612 ;
			RECT	24.659 21.548 24.691 21.612 ;
			RECT	24.827 21.548 24.859 21.612 ;
			RECT	24.995 21.548 25.027 21.612 ;
			RECT	25.163 21.548 25.195 21.612 ;
			RECT	25.331 21.548 25.363 21.612 ;
			RECT	25.499 21.548 25.531 21.612 ;
			RECT	25.667 21.548 25.699 21.612 ;
			RECT	25.835 21.548 25.867 21.612 ;
			RECT	26.003 21.548 26.035 21.612 ;
			RECT	26.171 21.548 26.203 21.612 ;
			RECT	26.339 21.548 26.371 21.612 ;
			RECT	26.507 21.548 26.539 21.612 ;
			RECT	26.675 21.548 26.707 21.612 ;
			RECT	26.843 21.548 26.875 21.612 ;
			RECT	27.011 21.548 27.043 21.612 ;
			RECT	27.179 21.548 27.211 21.612 ;
			RECT	27.347 21.548 27.379 21.612 ;
			RECT	27.515 21.548 27.547 21.612 ;
			RECT	27.683 21.548 27.715 21.612 ;
			RECT	27.851 21.548 27.883 21.612 ;
			RECT	28.019 21.548 28.051 21.612 ;
			RECT	28.187 21.548 28.219 21.612 ;
			RECT	28.355 21.548 28.387 21.612 ;
			RECT	28.523 21.548 28.555 21.612 ;
			RECT	28.691 21.548 28.723 21.612 ;
			RECT	28.859 21.548 28.891 21.612 ;
			RECT	29.027 21.548 29.059 21.612 ;
			RECT	29.195 21.548 29.227 21.612 ;
			RECT	29.363 21.548 29.395 21.612 ;
			RECT	29.531 21.548 29.563 21.612 ;
			RECT	29.699 21.548 29.731 21.612 ;
			RECT	29.867 21.548 29.899 21.612 ;
			RECT	30.035 21.548 30.067 21.612 ;
			RECT	30.203 21.548 30.235 21.612 ;
			RECT	30.371 21.548 30.403 21.612 ;
			RECT	30.539 21.548 30.571 21.612 ;
			RECT	30.707 21.548 30.739 21.612 ;
			RECT	30.875 21.548 30.907 21.612 ;
			RECT	31.043 21.548 31.075 21.612 ;
			RECT	31.211 21.548 31.243 21.612 ;
			RECT	31.379 21.548 31.411 21.612 ;
			RECT	31.547 21.548 31.579 21.612 ;
			RECT	31.715 21.548 31.747 21.612 ;
			RECT	31.883 21.548 31.915 21.612 ;
			RECT	32.051 21.548 32.083 21.612 ;
			RECT	32.219 21.548 32.251 21.612 ;
			RECT	32.387 21.548 32.419 21.612 ;
			RECT	32.555 21.548 32.587 21.612 ;
			RECT	32.723 21.548 32.755 21.612 ;
			RECT	32.891 21.548 32.923 21.612 ;
			RECT	33.059 21.548 33.091 21.612 ;
			RECT	33.227 21.548 33.259 21.612 ;
			RECT	33.395 21.548 33.427 21.612 ;
			RECT	33.563 21.548 33.595 21.612 ;
			RECT	33.731 21.548 33.763 21.612 ;
			RECT	33.899 21.548 33.931 21.612 ;
			RECT	34.067 21.548 34.099 21.612 ;
			RECT	34.235 21.548 34.267 21.612 ;
			RECT	34.403 21.548 34.435 21.612 ;
			RECT	34.571 21.548 34.603 21.612 ;
			RECT	34.739 21.548 34.771 21.612 ;
			RECT	34.907 21.548 34.939 21.612 ;
			RECT	35.075 21.548 35.107 21.612 ;
			RECT	35.243 21.548 35.275 21.612 ;
			RECT	35.411 21.548 35.443 21.612 ;
			RECT	35.579 21.548 35.611 21.612 ;
			RECT	35.747 21.548 35.779 21.612 ;
			RECT	35.915 21.548 35.947 21.612 ;
			RECT	36.083 21.548 36.115 21.612 ;
			RECT	36.251 21.548 36.283 21.612 ;
			RECT	36.419 21.548 36.451 21.612 ;
			RECT	36.587 21.548 36.619 21.612 ;
			RECT	36.755 21.548 36.787 21.612 ;
			RECT	36.923 21.548 36.955 21.612 ;
			RECT	37.091 21.548 37.123 21.612 ;
			RECT	37.259 21.548 37.291 21.612 ;
			RECT	37.427 21.548 37.459 21.612 ;
			RECT	37.595 21.548 37.627 21.612 ;
			RECT	37.763 21.548 37.795 21.612 ;
			RECT	37.931 21.548 37.963 21.612 ;
			RECT	38.099 21.548 38.131 21.612 ;
			RECT	38.267 21.548 38.299 21.612 ;
			RECT	38.435 21.548 38.467 21.612 ;
			RECT	38.603 21.548 38.635 21.612 ;
			RECT	38.771 21.548 38.803 21.612 ;
			RECT	38.939 21.548 38.971 21.612 ;
			RECT	39.107 21.548 39.139 21.612 ;
			RECT	39.275 21.548 39.307 21.612 ;
			RECT	39.443 21.548 39.475 21.612 ;
			RECT	39.611 21.548 39.643 21.612 ;
			RECT	39.779 21.548 39.811 21.612 ;
			RECT	39.947 21.548 39.979 21.612 ;
			RECT	40.115 21.548 40.147 21.612 ;
			RECT	40.283 21.548 40.315 21.612 ;
			RECT	40.451 21.548 40.483 21.612 ;
			RECT	40.619 21.548 40.651 21.612 ;
			RECT	40.787 21.548 40.819 21.612 ;
			RECT	40.955 21.548 40.987 21.612 ;
			RECT	41.123 21.548 41.155 21.612 ;
			RECT	41.291 21.548 41.323 21.612 ;
			RECT	41.459 21.548 41.491 21.612 ;
			RECT	41.627 21.548 41.659 21.612 ;
			RECT	41.795 21.548 41.827 21.612 ;
			RECT	41.963 21.548 41.995 21.612 ;
			RECT	42.131 21.548 42.163 21.612 ;
			RECT	42.299 21.548 42.331 21.612 ;
			RECT	42.467 21.548 42.499 21.612 ;
			RECT	42.635 21.548 42.667 21.612 ;
			RECT	42.803 21.548 42.835 21.612 ;
			RECT	42.971 21.548 43.003 21.612 ;
			RECT	43.139 21.548 43.171 21.612 ;
			RECT	43.307 21.548 43.339 21.612 ;
			RECT	43.475 21.548 43.507 21.612 ;
			RECT	43.643 21.548 43.675 21.612 ;
			RECT	43.811 21.548 43.843 21.612 ;
			RECT	43.979 21.548 44.011 21.612 ;
			RECT	44.147 21.548 44.179 21.612 ;
			RECT	44.315 21.548 44.347 21.612 ;
			RECT	44.483 21.548 44.515 21.612 ;
			RECT	44.651 21.548 44.683 21.612 ;
			RECT	44.819 21.548 44.851 21.612 ;
			RECT	44.987 21.548 45.019 21.612 ;
			RECT	45.155 21.548 45.187 21.612 ;
			RECT	45.323 21.548 45.355 21.612 ;
			RECT	45.491 21.548 45.523 21.612 ;
			RECT	45.659 21.548 45.691 21.612 ;
			RECT	45.827 21.548 45.859 21.612 ;
			RECT	45.995 21.548 46.027 21.612 ;
			RECT	46.163 21.548 46.195 21.612 ;
			RECT	46.331 21.548 46.363 21.612 ;
			RECT	46.499 21.548 46.531 21.612 ;
			RECT	46.667 21.548 46.699 21.612 ;
			RECT	46.835 21.548 46.867 21.612 ;
			RECT	47.003 21.548 47.035 21.612 ;
			RECT	47.171 21.548 47.203 21.612 ;
			RECT	47.339 21.548 47.371 21.612 ;
			RECT	47.507 21.548 47.539 21.612 ;
			RECT	47.675 21.548 47.707 21.612 ;
			RECT	47.843 21.548 47.875 21.612 ;
			RECT	48.011 21.548 48.043 21.612 ;
			RECT	48.179 21.548 48.211 21.612 ;
			RECT	48.347 21.548 48.379 21.612 ;
			RECT	48.515 21.548 48.547 21.612 ;
			RECT	48.683 21.548 48.715 21.612 ;
			RECT	48.851 21.548 48.883 21.612 ;
			RECT	49.019 21.548 49.051 21.612 ;
			RECT	49.187 21.548 49.219 21.612 ;
			RECT	49.318 21.564 49.35 21.596 ;
			RECT	49.439 21.564 49.471 21.596 ;
			RECT	49.569 21.548 49.601 21.612 ;
			RECT	51.881 21.548 51.913 21.612 ;
			RECT	53.132 21.548 53.196 21.612 ;
			RECT	53.812 21.548 53.844 21.612 ;
			RECT	54.251 21.548 54.283 21.612 ;
			RECT	55.562 21.548 55.626 21.612 ;
			RECT	58.603 21.548 58.635 21.612 ;
			RECT	58.733 21.564 58.765 21.596 ;
			RECT	58.854 21.564 58.886 21.596 ;
			RECT	58.985 21.548 59.017 21.612 ;
			RECT	59.153 21.548 59.185 21.612 ;
			RECT	59.321 21.548 59.353 21.612 ;
			RECT	59.489 21.548 59.521 21.612 ;
			RECT	59.657 21.548 59.689 21.612 ;
			RECT	59.825 21.548 59.857 21.612 ;
			RECT	59.993 21.548 60.025 21.612 ;
			RECT	60.161 21.548 60.193 21.612 ;
			RECT	60.329 21.548 60.361 21.612 ;
			RECT	60.497 21.548 60.529 21.612 ;
			RECT	60.665 21.548 60.697 21.612 ;
			RECT	60.833 21.548 60.865 21.612 ;
			RECT	61.001 21.548 61.033 21.612 ;
			RECT	61.169 21.548 61.201 21.612 ;
			RECT	61.337 21.548 61.369 21.612 ;
			RECT	61.505 21.548 61.537 21.612 ;
			RECT	61.673 21.548 61.705 21.612 ;
			RECT	61.841 21.548 61.873 21.612 ;
			RECT	62.009 21.548 62.041 21.612 ;
			RECT	62.177 21.548 62.209 21.612 ;
			RECT	62.345 21.548 62.377 21.612 ;
			RECT	62.513 21.548 62.545 21.612 ;
			RECT	62.681 21.548 62.713 21.612 ;
			RECT	62.849 21.548 62.881 21.612 ;
			RECT	63.017 21.548 63.049 21.612 ;
			RECT	63.185 21.548 63.217 21.612 ;
			RECT	63.353 21.548 63.385 21.612 ;
			RECT	63.521 21.548 63.553 21.612 ;
			RECT	63.689 21.548 63.721 21.612 ;
			RECT	63.857 21.548 63.889 21.612 ;
			RECT	64.025 21.548 64.057 21.612 ;
			RECT	64.193 21.548 64.225 21.612 ;
			RECT	64.361 21.548 64.393 21.612 ;
			RECT	64.529 21.548 64.561 21.612 ;
			RECT	64.697 21.548 64.729 21.612 ;
			RECT	64.865 21.548 64.897 21.612 ;
			RECT	65.033 21.548 65.065 21.612 ;
			RECT	65.201 21.548 65.233 21.612 ;
			RECT	65.369 21.548 65.401 21.612 ;
			RECT	65.537 21.548 65.569 21.612 ;
			RECT	65.705 21.548 65.737 21.612 ;
			RECT	65.873 21.548 65.905 21.612 ;
			RECT	66.041 21.548 66.073 21.612 ;
			RECT	66.209 21.548 66.241 21.612 ;
			RECT	66.377 21.548 66.409 21.612 ;
			RECT	66.545 21.548 66.577 21.612 ;
			RECT	66.713 21.548 66.745 21.612 ;
			RECT	66.881 21.548 66.913 21.612 ;
			RECT	67.049 21.548 67.081 21.612 ;
			RECT	67.217 21.548 67.249 21.612 ;
			RECT	67.385 21.548 67.417 21.612 ;
			RECT	67.553 21.548 67.585 21.612 ;
			RECT	67.721 21.548 67.753 21.612 ;
			RECT	67.889 21.548 67.921 21.612 ;
			RECT	68.057 21.548 68.089 21.612 ;
			RECT	68.225 21.548 68.257 21.612 ;
			RECT	68.393 21.548 68.425 21.612 ;
			RECT	68.561 21.548 68.593 21.612 ;
			RECT	68.729 21.548 68.761 21.612 ;
			RECT	68.897 21.548 68.929 21.612 ;
			RECT	69.065 21.548 69.097 21.612 ;
			RECT	69.233 21.548 69.265 21.612 ;
			RECT	69.401 21.548 69.433 21.612 ;
			RECT	69.569 21.548 69.601 21.612 ;
			RECT	69.737 21.548 69.769 21.612 ;
			RECT	69.905 21.548 69.937 21.612 ;
			RECT	70.073 21.548 70.105 21.612 ;
			RECT	70.241 21.548 70.273 21.612 ;
			RECT	70.409 21.548 70.441 21.612 ;
			RECT	70.577 21.548 70.609 21.612 ;
			RECT	70.745 21.548 70.777 21.612 ;
			RECT	70.913 21.548 70.945 21.612 ;
			RECT	71.081 21.548 71.113 21.612 ;
			RECT	71.249 21.548 71.281 21.612 ;
			RECT	71.417 21.548 71.449 21.612 ;
			RECT	71.585 21.548 71.617 21.612 ;
			RECT	71.753 21.548 71.785 21.612 ;
			RECT	71.921 21.548 71.953 21.612 ;
			RECT	72.089 21.548 72.121 21.612 ;
			RECT	72.257 21.548 72.289 21.612 ;
			RECT	72.425 21.548 72.457 21.612 ;
			RECT	72.593 21.548 72.625 21.612 ;
			RECT	72.761 21.548 72.793 21.612 ;
			RECT	72.929 21.548 72.961 21.612 ;
			RECT	73.097 21.548 73.129 21.612 ;
			RECT	73.265 21.548 73.297 21.612 ;
			RECT	73.433 21.548 73.465 21.612 ;
			RECT	73.601 21.548 73.633 21.612 ;
			RECT	73.769 21.548 73.801 21.612 ;
			RECT	73.937 21.548 73.969 21.612 ;
			RECT	74.105 21.548 74.137 21.612 ;
			RECT	74.273 21.548 74.305 21.612 ;
			RECT	74.441 21.548 74.473 21.612 ;
			RECT	74.609 21.548 74.641 21.612 ;
			RECT	74.777 21.548 74.809 21.612 ;
			RECT	74.945 21.548 74.977 21.612 ;
			RECT	75.113 21.548 75.145 21.612 ;
			RECT	75.281 21.548 75.313 21.612 ;
			RECT	75.449 21.548 75.481 21.612 ;
			RECT	75.617 21.548 75.649 21.612 ;
			RECT	75.785 21.548 75.817 21.612 ;
			RECT	75.953 21.548 75.985 21.612 ;
			RECT	76.121 21.548 76.153 21.612 ;
			RECT	76.289 21.548 76.321 21.612 ;
			RECT	76.457 21.548 76.489 21.612 ;
			RECT	76.625 21.548 76.657 21.612 ;
			RECT	76.793 21.548 76.825 21.612 ;
			RECT	76.961 21.548 76.993 21.612 ;
			RECT	77.129 21.548 77.161 21.612 ;
			RECT	77.297 21.548 77.329 21.612 ;
			RECT	77.465 21.548 77.497 21.612 ;
			RECT	77.633 21.548 77.665 21.612 ;
			RECT	77.801 21.548 77.833 21.612 ;
			RECT	77.969 21.548 78.001 21.612 ;
			RECT	78.137 21.548 78.169 21.612 ;
			RECT	78.305 21.548 78.337 21.612 ;
			RECT	78.473 21.548 78.505 21.612 ;
			RECT	78.641 21.548 78.673 21.612 ;
			RECT	78.809 21.548 78.841 21.612 ;
			RECT	78.977 21.548 79.009 21.612 ;
			RECT	79.145 21.548 79.177 21.612 ;
			RECT	79.313 21.548 79.345 21.612 ;
			RECT	79.481 21.548 79.513 21.612 ;
			RECT	79.649 21.548 79.681 21.612 ;
			RECT	79.817 21.548 79.849 21.612 ;
			RECT	79.985 21.548 80.017 21.612 ;
			RECT	80.153 21.548 80.185 21.612 ;
			RECT	80.321 21.548 80.353 21.612 ;
			RECT	80.489 21.548 80.521 21.612 ;
			RECT	80.657 21.548 80.689 21.612 ;
			RECT	80.825 21.548 80.857 21.612 ;
			RECT	80.993 21.548 81.025 21.612 ;
			RECT	81.161 21.548 81.193 21.612 ;
			RECT	81.329 21.548 81.361 21.612 ;
			RECT	81.497 21.548 81.529 21.612 ;
			RECT	81.665 21.548 81.697 21.612 ;
			RECT	81.833 21.548 81.865 21.612 ;
			RECT	82.001 21.548 82.033 21.612 ;
			RECT	82.169 21.548 82.201 21.612 ;
			RECT	82.337 21.548 82.369 21.612 ;
			RECT	82.505 21.548 82.537 21.612 ;
			RECT	82.673 21.548 82.705 21.612 ;
			RECT	82.841 21.548 82.873 21.612 ;
			RECT	83.009 21.548 83.041 21.612 ;
			RECT	83.177 21.548 83.209 21.612 ;
			RECT	83.345 21.548 83.377 21.612 ;
			RECT	83.513 21.548 83.545 21.612 ;
			RECT	83.681 21.548 83.713 21.612 ;
			RECT	83.849 21.548 83.881 21.612 ;
			RECT	84.017 21.548 84.049 21.612 ;
			RECT	84.185 21.548 84.217 21.612 ;
			RECT	84.353 21.548 84.385 21.612 ;
			RECT	84.521 21.548 84.553 21.612 ;
			RECT	84.689 21.548 84.721 21.612 ;
			RECT	84.857 21.548 84.889 21.612 ;
			RECT	85.025 21.548 85.057 21.612 ;
			RECT	85.193 21.548 85.225 21.612 ;
			RECT	85.361 21.548 85.393 21.612 ;
			RECT	85.529 21.548 85.561 21.612 ;
			RECT	85.697 21.548 85.729 21.612 ;
			RECT	85.865 21.548 85.897 21.612 ;
			RECT	86.033 21.548 86.065 21.612 ;
			RECT	86.201 21.548 86.233 21.612 ;
			RECT	86.369 21.548 86.401 21.612 ;
			RECT	86.537 21.548 86.569 21.612 ;
			RECT	86.705 21.548 86.737 21.612 ;
			RECT	86.873 21.548 86.905 21.612 ;
			RECT	87.041 21.548 87.073 21.612 ;
			RECT	87.209 21.548 87.241 21.612 ;
			RECT	87.377 21.548 87.409 21.612 ;
			RECT	87.545 21.548 87.577 21.612 ;
			RECT	87.713 21.548 87.745 21.612 ;
			RECT	87.881 21.548 87.913 21.612 ;
			RECT	88.049 21.548 88.081 21.612 ;
			RECT	88.217 21.548 88.249 21.612 ;
			RECT	88.385 21.548 88.417 21.612 ;
			RECT	88.553 21.548 88.585 21.612 ;
			RECT	88.721 21.548 88.753 21.612 ;
			RECT	88.889 21.548 88.921 21.612 ;
			RECT	89.057 21.548 89.089 21.612 ;
			RECT	89.225 21.548 89.257 21.612 ;
			RECT	89.393 21.548 89.425 21.612 ;
			RECT	89.561 21.548 89.593 21.612 ;
			RECT	89.729 21.548 89.761 21.612 ;
			RECT	89.897 21.548 89.929 21.612 ;
			RECT	90.065 21.548 90.097 21.612 ;
			RECT	90.233 21.548 90.265 21.612 ;
			RECT	90.401 21.548 90.433 21.612 ;
			RECT	90.569 21.548 90.601 21.612 ;
			RECT	90.737 21.548 90.769 21.612 ;
			RECT	90.905 21.548 90.937 21.612 ;
			RECT	91.073 21.548 91.105 21.612 ;
			RECT	91.241 21.548 91.273 21.612 ;
			RECT	91.409 21.548 91.441 21.612 ;
			RECT	91.577 21.548 91.609 21.612 ;
			RECT	91.745 21.548 91.777 21.612 ;
			RECT	91.913 21.548 91.945 21.612 ;
			RECT	92.081 21.548 92.113 21.612 ;
			RECT	92.249 21.548 92.281 21.612 ;
			RECT	92.417 21.548 92.449 21.612 ;
			RECT	92.585 21.548 92.617 21.612 ;
			RECT	92.753 21.548 92.785 21.612 ;
			RECT	92.921 21.548 92.953 21.612 ;
			RECT	93.089 21.548 93.121 21.612 ;
			RECT	93.257 21.548 93.289 21.612 ;
			RECT	93.425 21.548 93.457 21.612 ;
			RECT	93.593 21.548 93.625 21.612 ;
			RECT	93.761 21.548 93.793 21.612 ;
			RECT	93.929 21.548 93.961 21.612 ;
			RECT	94.097 21.548 94.129 21.612 ;
			RECT	94.265 21.548 94.297 21.612 ;
			RECT	94.433 21.548 94.465 21.612 ;
			RECT	94.601 21.548 94.633 21.612 ;
			RECT	94.769 21.548 94.801 21.612 ;
			RECT	94.937 21.548 94.969 21.612 ;
			RECT	95.105 21.548 95.137 21.612 ;
			RECT	95.273 21.548 95.305 21.612 ;
			RECT	95.441 21.548 95.473 21.612 ;
			RECT	95.609 21.548 95.641 21.612 ;
			RECT	95.777 21.548 95.809 21.612 ;
			RECT	95.945 21.548 95.977 21.612 ;
			RECT	96.113 21.548 96.145 21.612 ;
			RECT	96.281 21.548 96.313 21.612 ;
			RECT	96.449 21.548 96.481 21.612 ;
			RECT	96.617 21.548 96.649 21.612 ;
			RECT	96.785 21.548 96.817 21.612 ;
			RECT	96.953 21.548 96.985 21.612 ;
			RECT	97.121 21.548 97.153 21.612 ;
			RECT	97.289 21.548 97.321 21.612 ;
			RECT	97.457 21.548 97.489 21.612 ;
			RECT	97.625 21.548 97.657 21.612 ;
			RECT	97.793 21.548 97.825 21.612 ;
			RECT	97.961 21.548 97.993 21.612 ;
			RECT	98.129 21.548 98.161 21.612 ;
			RECT	98.297 21.548 98.329 21.612 ;
			RECT	98.465 21.548 98.497 21.612 ;
			RECT	98.633 21.548 98.665 21.612 ;
			RECT	98.801 21.548 98.833 21.612 ;
			RECT	98.969 21.548 99.001 21.612 ;
			RECT	99.137 21.548 99.169 21.612 ;
			RECT	99.305 21.548 99.337 21.612 ;
			RECT	99.473 21.548 99.505 21.612 ;
			RECT	99.641 21.548 99.673 21.612 ;
			RECT	99.809 21.548 99.841 21.612 ;
			RECT	99.977 21.548 100.009 21.612 ;
			RECT	100.145 21.548 100.177 21.612 ;
			RECT	100.313 21.548 100.345 21.612 ;
			RECT	100.481 21.548 100.513 21.612 ;
			RECT	100.649 21.548 100.681 21.612 ;
			RECT	100.817 21.548 100.849 21.612 ;
			RECT	100.985 21.548 101.017 21.612 ;
			RECT	101.153 21.548 101.185 21.612 ;
			RECT	101.321 21.548 101.353 21.612 ;
			RECT	101.489 21.548 101.521 21.612 ;
			RECT	101.657 21.548 101.689 21.612 ;
			RECT	101.825 21.548 101.857 21.612 ;
			RECT	101.993 21.548 102.025 21.612 ;
			RECT	102.123 21.564 102.155 21.596 ;
			RECT	102.245 21.569 102.277 21.601 ;
			RECT	102.375 21.548 102.407 21.612 ;
			RECT	103.795 21.548 103.827 21.612 ;
			RECT	103.925 21.569 103.957 21.601 ;
			RECT	104.047 21.564 104.079 21.596 ;
			RECT	104.177 21.548 104.209 21.612 ;
			RECT	104.345 21.548 104.377 21.612 ;
			RECT	104.513 21.548 104.545 21.612 ;
			RECT	104.681 21.548 104.713 21.612 ;
			RECT	104.849 21.548 104.881 21.612 ;
			RECT	105.017 21.548 105.049 21.612 ;
			RECT	105.185 21.548 105.217 21.612 ;
			RECT	105.353 21.548 105.385 21.612 ;
			RECT	105.521 21.548 105.553 21.612 ;
			RECT	105.689 21.548 105.721 21.612 ;
			RECT	105.857 21.548 105.889 21.612 ;
			RECT	106.025 21.548 106.057 21.612 ;
			RECT	106.193 21.548 106.225 21.612 ;
			RECT	106.361 21.548 106.393 21.612 ;
			RECT	106.529 21.548 106.561 21.612 ;
			RECT	106.697 21.548 106.729 21.612 ;
			RECT	106.865 21.548 106.897 21.612 ;
			RECT	107.033 21.548 107.065 21.612 ;
			RECT	107.201 21.548 107.233 21.612 ;
			RECT	107.369 21.548 107.401 21.612 ;
			RECT	107.537 21.548 107.569 21.612 ;
			RECT	107.705 21.548 107.737 21.612 ;
			RECT	107.873 21.548 107.905 21.612 ;
			RECT	108.041 21.548 108.073 21.612 ;
			RECT	108.209 21.548 108.241 21.612 ;
			RECT	108.377 21.548 108.409 21.612 ;
			RECT	108.545 21.548 108.577 21.612 ;
			RECT	108.713 21.548 108.745 21.612 ;
			RECT	108.881 21.548 108.913 21.612 ;
			RECT	109.049 21.548 109.081 21.612 ;
			RECT	109.217 21.548 109.249 21.612 ;
			RECT	109.385 21.548 109.417 21.612 ;
			RECT	109.553 21.548 109.585 21.612 ;
			RECT	109.721 21.548 109.753 21.612 ;
			RECT	109.889 21.548 109.921 21.612 ;
			RECT	110.057 21.548 110.089 21.612 ;
			RECT	110.225 21.548 110.257 21.612 ;
			RECT	110.393 21.548 110.425 21.612 ;
			RECT	110.561 21.548 110.593 21.612 ;
			RECT	110.729 21.548 110.761 21.612 ;
			RECT	110.897 21.548 110.929 21.612 ;
			RECT	111.065 21.548 111.097 21.612 ;
			RECT	111.233 21.548 111.265 21.612 ;
			RECT	111.401 21.548 111.433 21.612 ;
			RECT	111.569 21.548 111.601 21.612 ;
			RECT	111.737 21.548 111.769 21.612 ;
			RECT	111.905 21.548 111.937 21.612 ;
			RECT	112.073 21.548 112.105 21.612 ;
			RECT	112.241 21.548 112.273 21.612 ;
			RECT	112.409 21.548 112.441 21.612 ;
			RECT	112.577 21.548 112.609 21.612 ;
			RECT	112.745 21.548 112.777 21.612 ;
			RECT	112.913 21.548 112.945 21.612 ;
			RECT	113.081 21.548 113.113 21.612 ;
			RECT	113.249 21.548 113.281 21.612 ;
			RECT	113.417 21.548 113.449 21.612 ;
			RECT	113.585 21.548 113.617 21.612 ;
			RECT	113.753 21.548 113.785 21.612 ;
			RECT	113.921 21.548 113.953 21.612 ;
			RECT	114.089 21.548 114.121 21.612 ;
			RECT	114.257 21.548 114.289 21.612 ;
			RECT	114.425 21.548 114.457 21.612 ;
			RECT	114.593 21.548 114.625 21.612 ;
			RECT	114.761 21.548 114.793 21.612 ;
			RECT	114.929 21.548 114.961 21.612 ;
			RECT	115.097 21.548 115.129 21.612 ;
			RECT	115.265 21.548 115.297 21.612 ;
			RECT	115.433 21.548 115.465 21.612 ;
			RECT	115.601 21.548 115.633 21.612 ;
			RECT	115.769 21.548 115.801 21.612 ;
			RECT	115.937 21.548 115.969 21.612 ;
			RECT	116.105 21.548 116.137 21.612 ;
			RECT	116.273 21.548 116.305 21.612 ;
			RECT	116.441 21.548 116.473 21.612 ;
			RECT	116.609 21.548 116.641 21.612 ;
			RECT	116.777 21.548 116.809 21.612 ;
			RECT	116.945 21.548 116.977 21.612 ;
			RECT	117.113 21.548 117.145 21.612 ;
			RECT	117.281 21.548 117.313 21.612 ;
			RECT	117.449 21.548 117.481 21.612 ;
			RECT	117.617 21.548 117.649 21.612 ;
			RECT	117.785 21.548 117.817 21.612 ;
			RECT	117.953 21.548 117.985 21.612 ;
			RECT	118.121 21.548 118.153 21.612 ;
			RECT	118.289 21.548 118.321 21.612 ;
			RECT	118.457 21.548 118.489 21.612 ;
			RECT	118.625 21.548 118.657 21.612 ;
			RECT	118.793 21.548 118.825 21.612 ;
			RECT	118.961 21.548 118.993 21.612 ;
			RECT	119.129 21.548 119.161 21.612 ;
			RECT	119.297 21.548 119.329 21.612 ;
			RECT	119.465 21.548 119.497 21.612 ;
			RECT	119.633 21.548 119.665 21.612 ;
			RECT	119.801 21.548 119.833 21.612 ;
			RECT	119.969 21.548 120.001 21.612 ;
			RECT	120.137 21.548 120.169 21.612 ;
			RECT	120.305 21.548 120.337 21.612 ;
			RECT	120.473 21.548 120.505 21.612 ;
			RECT	120.641 21.548 120.673 21.612 ;
			RECT	120.809 21.548 120.841 21.612 ;
			RECT	120.977 21.548 121.009 21.612 ;
			RECT	121.145 21.548 121.177 21.612 ;
			RECT	121.313 21.548 121.345 21.612 ;
			RECT	121.481 21.548 121.513 21.612 ;
			RECT	121.649 21.548 121.681 21.612 ;
			RECT	121.817 21.548 121.849 21.612 ;
			RECT	121.985 21.548 122.017 21.612 ;
			RECT	122.153 21.548 122.185 21.612 ;
			RECT	122.321 21.548 122.353 21.612 ;
			RECT	122.489 21.548 122.521 21.612 ;
			RECT	122.657 21.548 122.689 21.612 ;
			RECT	122.825 21.548 122.857 21.612 ;
			RECT	122.993 21.548 123.025 21.612 ;
			RECT	123.161 21.548 123.193 21.612 ;
			RECT	123.329 21.548 123.361 21.612 ;
			RECT	123.497 21.548 123.529 21.612 ;
			RECT	123.665 21.548 123.697 21.612 ;
			RECT	123.833 21.548 123.865 21.612 ;
			RECT	124.001 21.548 124.033 21.612 ;
			RECT	124.169 21.548 124.201 21.612 ;
			RECT	124.337 21.548 124.369 21.612 ;
			RECT	124.505 21.548 124.537 21.612 ;
			RECT	124.673 21.548 124.705 21.612 ;
			RECT	124.841 21.548 124.873 21.612 ;
			RECT	125.009 21.548 125.041 21.612 ;
			RECT	125.177 21.548 125.209 21.612 ;
			RECT	125.345 21.548 125.377 21.612 ;
			RECT	125.513 21.548 125.545 21.612 ;
			RECT	125.681 21.548 125.713 21.612 ;
			RECT	125.849 21.548 125.881 21.612 ;
			RECT	126.017 21.548 126.049 21.612 ;
			RECT	126.185 21.548 126.217 21.612 ;
			RECT	126.353 21.548 126.385 21.612 ;
			RECT	126.521 21.548 126.553 21.612 ;
			RECT	126.689 21.548 126.721 21.612 ;
			RECT	126.857 21.548 126.889 21.612 ;
			RECT	127.025 21.548 127.057 21.612 ;
			RECT	127.193 21.548 127.225 21.612 ;
			RECT	127.361 21.548 127.393 21.612 ;
			RECT	127.529 21.548 127.561 21.612 ;
			RECT	127.697 21.548 127.729 21.612 ;
			RECT	127.865 21.548 127.897 21.612 ;
			RECT	128.033 21.548 128.065 21.612 ;
			RECT	128.201 21.548 128.233 21.612 ;
			RECT	128.369 21.548 128.401 21.612 ;
			RECT	128.537 21.548 128.569 21.612 ;
			RECT	128.705 21.548 128.737 21.612 ;
			RECT	128.873 21.548 128.905 21.612 ;
			RECT	129.041 21.548 129.073 21.612 ;
			RECT	129.209 21.548 129.241 21.612 ;
			RECT	129.377 21.548 129.409 21.612 ;
			RECT	129.545 21.548 129.577 21.612 ;
			RECT	129.713 21.548 129.745 21.612 ;
			RECT	129.881 21.548 129.913 21.612 ;
			RECT	130.049 21.548 130.081 21.612 ;
			RECT	130.217 21.548 130.249 21.612 ;
			RECT	130.385 21.548 130.417 21.612 ;
			RECT	130.553 21.548 130.585 21.612 ;
			RECT	130.721 21.548 130.753 21.612 ;
			RECT	130.889 21.548 130.921 21.612 ;
			RECT	131.057 21.548 131.089 21.612 ;
			RECT	131.225 21.548 131.257 21.612 ;
			RECT	131.393 21.548 131.425 21.612 ;
			RECT	131.561 21.548 131.593 21.612 ;
			RECT	131.729 21.548 131.761 21.612 ;
			RECT	131.897 21.548 131.929 21.612 ;
			RECT	132.065 21.548 132.097 21.612 ;
			RECT	132.233 21.548 132.265 21.612 ;
			RECT	132.401 21.548 132.433 21.612 ;
			RECT	132.569 21.548 132.601 21.612 ;
			RECT	132.737 21.548 132.769 21.612 ;
			RECT	132.905 21.548 132.937 21.612 ;
			RECT	133.073 21.548 133.105 21.612 ;
			RECT	133.241 21.548 133.273 21.612 ;
			RECT	133.409 21.548 133.441 21.612 ;
			RECT	133.577 21.548 133.609 21.612 ;
			RECT	133.745 21.548 133.777 21.612 ;
			RECT	133.913 21.548 133.945 21.612 ;
			RECT	134.081 21.548 134.113 21.612 ;
			RECT	134.249 21.548 134.281 21.612 ;
			RECT	134.417 21.548 134.449 21.612 ;
			RECT	134.585 21.548 134.617 21.612 ;
			RECT	134.753 21.548 134.785 21.612 ;
			RECT	134.921 21.548 134.953 21.612 ;
			RECT	135.089 21.548 135.121 21.612 ;
			RECT	135.257 21.548 135.289 21.612 ;
			RECT	135.425 21.548 135.457 21.612 ;
			RECT	135.593 21.548 135.625 21.612 ;
			RECT	135.761 21.548 135.793 21.612 ;
			RECT	135.929 21.548 135.961 21.612 ;
			RECT	136.097 21.548 136.129 21.612 ;
			RECT	136.265 21.548 136.297 21.612 ;
			RECT	136.433 21.548 136.465 21.612 ;
			RECT	136.601 21.548 136.633 21.612 ;
			RECT	136.769 21.548 136.801 21.612 ;
			RECT	136.937 21.548 136.969 21.612 ;
			RECT	137.105 21.548 137.137 21.612 ;
			RECT	137.273 21.548 137.305 21.612 ;
			RECT	137.441 21.548 137.473 21.612 ;
			RECT	137.609 21.548 137.641 21.612 ;
			RECT	137.777 21.548 137.809 21.612 ;
			RECT	137.945 21.548 137.977 21.612 ;
			RECT	138.113 21.548 138.145 21.612 ;
			RECT	138.281 21.548 138.313 21.612 ;
			RECT	138.449 21.548 138.481 21.612 ;
			RECT	138.617 21.548 138.649 21.612 ;
			RECT	138.785 21.548 138.817 21.612 ;
			RECT	138.953 21.548 138.985 21.612 ;
			RECT	139.121 21.548 139.153 21.612 ;
			RECT	139.289 21.548 139.321 21.612 ;
			RECT	139.457 21.548 139.489 21.612 ;
			RECT	139.625 21.548 139.657 21.612 ;
			RECT	139.793 21.548 139.825 21.612 ;
			RECT	139.961 21.548 139.993 21.612 ;
			RECT	140.129 21.548 140.161 21.612 ;
			RECT	140.297 21.548 140.329 21.612 ;
			RECT	140.465 21.548 140.497 21.612 ;
			RECT	140.633 21.548 140.665 21.612 ;
			RECT	140.801 21.548 140.833 21.612 ;
			RECT	140.969 21.548 141.001 21.612 ;
			RECT	141.137 21.548 141.169 21.612 ;
			RECT	141.305 21.548 141.337 21.612 ;
			RECT	141.473 21.548 141.505 21.612 ;
			RECT	141.641 21.548 141.673 21.612 ;
			RECT	141.809 21.548 141.841 21.612 ;
			RECT	141.977 21.548 142.009 21.612 ;
			RECT	142.145 21.548 142.177 21.612 ;
			RECT	142.313 21.548 142.345 21.612 ;
			RECT	142.481 21.548 142.513 21.612 ;
			RECT	142.649 21.548 142.681 21.612 ;
			RECT	142.817 21.548 142.849 21.612 ;
			RECT	142.985 21.548 143.017 21.612 ;
			RECT	143.153 21.548 143.185 21.612 ;
			RECT	143.321 21.548 143.353 21.612 ;
			RECT	143.489 21.548 143.521 21.612 ;
			RECT	143.657 21.548 143.689 21.612 ;
			RECT	143.825 21.548 143.857 21.612 ;
			RECT	143.993 21.548 144.025 21.612 ;
			RECT	144.161 21.548 144.193 21.612 ;
			RECT	144.329 21.548 144.361 21.612 ;
			RECT	144.497 21.548 144.529 21.612 ;
			RECT	144.665 21.548 144.697 21.612 ;
			RECT	144.833 21.548 144.865 21.612 ;
			RECT	145.001 21.548 145.033 21.612 ;
			RECT	145.169 21.548 145.201 21.612 ;
			RECT	145.337 21.548 145.369 21.612 ;
			RECT	145.505 21.548 145.537 21.612 ;
			RECT	145.673 21.548 145.705 21.612 ;
			RECT	145.841 21.548 145.873 21.612 ;
			RECT	146.009 21.548 146.041 21.612 ;
			RECT	146.177 21.548 146.209 21.612 ;
			RECT	146.345 21.548 146.377 21.612 ;
			RECT	146.513 21.548 146.545 21.612 ;
			RECT	146.681 21.548 146.713 21.612 ;
			RECT	146.849 21.548 146.881 21.612 ;
			RECT	147.017 21.548 147.049 21.612 ;
			RECT	147.185 21.548 147.217 21.612 ;
			RECT	147.316 21.564 147.348 21.596 ;
			RECT	147.437 21.564 147.469 21.596 ;
			RECT	147.567 21.548 147.599 21.612 ;
			RECT	149.879 21.548 149.911 21.612 ;
			RECT	151.13 21.548 151.194 21.612 ;
			RECT	151.81 21.548 151.842 21.612 ;
			RECT	152.249 21.548 152.281 21.612 ;
			RECT	153.56 21.548 153.624 21.612 ;
			RECT	156.601 21.548 156.633 21.612 ;
			RECT	156.731 21.564 156.763 21.596 ;
			RECT	156.852 21.564 156.884 21.596 ;
			RECT	156.983 21.548 157.015 21.612 ;
			RECT	157.151 21.548 157.183 21.612 ;
			RECT	157.319 21.548 157.351 21.612 ;
			RECT	157.487 21.548 157.519 21.612 ;
			RECT	157.655 21.548 157.687 21.612 ;
			RECT	157.823 21.548 157.855 21.612 ;
			RECT	157.991 21.548 158.023 21.612 ;
			RECT	158.159 21.548 158.191 21.612 ;
			RECT	158.327 21.548 158.359 21.612 ;
			RECT	158.495 21.548 158.527 21.612 ;
			RECT	158.663 21.548 158.695 21.612 ;
			RECT	158.831 21.548 158.863 21.612 ;
			RECT	158.999 21.548 159.031 21.612 ;
			RECT	159.167 21.548 159.199 21.612 ;
			RECT	159.335 21.548 159.367 21.612 ;
			RECT	159.503 21.548 159.535 21.612 ;
			RECT	159.671 21.548 159.703 21.612 ;
			RECT	159.839 21.548 159.871 21.612 ;
			RECT	160.007 21.548 160.039 21.612 ;
			RECT	160.175 21.548 160.207 21.612 ;
			RECT	160.343 21.548 160.375 21.612 ;
			RECT	160.511 21.548 160.543 21.612 ;
			RECT	160.679 21.548 160.711 21.612 ;
			RECT	160.847 21.548 160.879 21.612 ;
			RECT	161.015 21.548 161.047 21.612 ;
			RECT	161.183 21.548 161.215 21.612 ;
			RECT	161.351 21.548 161.383 21.612 ;
			RECT	161.519 21.548 161.551 21.612 ;
			RECT	161.687 21.548 161.719 21.612 ;
			RECT	161.855 21.548 161.887 21.612 ;
			RECT	162.023 21.548 162.055 21.612 ;
			RECT	162.191 21.548 162.223 21.612 ;
			RECT	162.359 21.548 162.391 21.612 ;
			RECT	162.527 21.548 162.559 21.612 ;
			RECT	162.695 21.548 162.727 21.612 ;
			RECT	162.863 21.548 162.895 21.612 ;
			RECT	163.031 21.548 163.063 21.612 ;
			RECT	163.199 21.548 163.231 21.612 ;
			RECT	163.367 21.548 163.399 21.612 ;
			RECT	163.535 21.548 163.567 21.612 ;
			RECT	163.703 21.548 163.735 21.612 ;
			RECT	163.871 21.548 163.903 21.612 ;
			RECT	164.039 21.548 164.071 21.612 ;
			RECT	164.207 21.548 164.239 21.612 ;
			RECT	164.375 21.548 164.407 21.612 ;
			RECT	164.543 21.548 164.575 21.612 ;
			RECT	164.711 21.548 164.743 21.612 ;
			RECT	164.879 21.548 164.911 21.612 ;
			RECT	165.047 21.548 165.079 21.612 ;
			RECT	165.215 21.548 165.247 21.612 ;
			RECT	165.383 21.548 165.415 21.612 ;
			RECT	165.551 21.548 165.583 21.612 ;
			RECT	165.719 21.548 165.751 21.612 ;
			RECT	165.887 21.548 165.919 21.612 ;
			RECT	166.055 21.548 166.087 21.612 ;
			RECT	166.223 21.548 166.255 21.612 ;
			RECT	166.391 21.548 166.423 21.612 ;
			RECT	166.559 21.548 166.591 21.612 ;
			RECT	166.727 21.548 166.759 21.612 ;
			RECT	166.895 21.548 166.927 21.612 ;
			RECT	167.063 21.548 167.095 21.612 ;
			RECT	167.231 21.548 167.263 21.612 ;
			RECT	167.399 21.548 167.431 21.612 ;
			RECT	167.567 21.548 167.599 21.612 ;
			RECT	167.735 21.548 167.767 21.612 ;
			RECT	167.903 21.548 167.935 21.612 ;
			RECT	168.071 21.548 168.103 21.612 ;
			RECT	168.239 21.548 168.271 21.612 ;
			RECT	168.407 21.548 168.439 21.612 ;
			RECT	168.575 21.548 168.607 21.612 ;
			RECT	168.743 21.548 168.775 21.612 ;
			RECT	168.911 21.548 168.943 21.612 ;
			RECT	169.079 21.548 169.111 21.612 ;
			RECT	169.247 21.548 169.279 21.612 ;
			RECT	169.415 21.548 169.447 21.612 ;
			RECT	169.583 21.548 169.615 21.612 ;
			RECT	169.751 21.548 169.783 21.612 ;
			RECT	169.919 21.548 169.951 21.612 ;
			RECT	170.087 21.548 170.119 21.612 ;
			RECT	170.255 21.548 170.287 21.612 ;
			RECT	170.423 21.548 170.455 21.612 ;
			RECT	170.591 21.548 170.623 21.612 ;
			RECT	170.759 21.548 170.791 21.612 ;
			RECT	170.927 21.548 170.959 21.612 ;
			RECT	171.095 21.548 171.127 21.612 ;
			RECT	171.263 21.548 171.295 21.612 ;
			RECT	171.431 21.548 171.463 21.612 ;
			RECT	171.599 21.548 171.631 21.612 ;
			RECT	171.767 21.548 171.799 21.612 ;
			RECT	171.935 21.548 171.967 21.612 ;
			RECT	172.103 21.548 172.135 21.612 ;
			RECT	172.271 21.548 172.303 21.612 ;
			RECT	172.439 21.548 172.471 21.612 ;
			RECT	172.607 21.548 172.639 21.612 ;
			RECT	172.775 21.548 172.807 21.612 ;
			RECT	172.943 21.548 172.975 21.612 ;
			RECT	173.111 21.548 173.143 21.612 ;
			RECT	173.279 21.548 173.311 21.612 ;
			RECT	173.447 21.548 173.479 21.612 ;
			RECT	173.615 21.548 173.647 21.612 ;
			RECT	173.783 21.548 173.815 21.612 ;
			RECT	173.951 21.548 173.983 21.612 ;
			RECT	174.119 21.548 174.151 21.612 ;
			RECT	174.287 21.548 174.319 21.612 ;
			RECT	174.455 21.548 174.487 21.612 ;
			RECT	174.623 21.548 174.655 21.612 ;
			RECT	174.791 21.548 174.823 21.612 ;
			RECT	174.959 21.548 174.991 21.612 ;
			RECT	175.127 21.548 175.159 21.612 ;
			RECT	175.295 21.548 175.327 21.612 ;
			RECT	175.463 21.548 175.495 21.612 ;
			RECT	175.631 21.548 175.663 21.612 ;
			RECT	175.799 21.548 175.831 21.612 ;
			RECT	175.967 21.548 175.999 21.612 ;
			RECT	176.135 21.548 176.167 21.612 ;
			RECT	176.303 21.548 176.335 21.612 ;
			RECT	176.471 21.548 176.503 21.612 ;
			RECT	176.639 21.548 176.671 21.612 ;
			RECT	176.807 21.548 176.839 21.612 ;
			RECT	176.975 21.548 177.007 21.612 ;
			RECT	177.143 21.548 177.175 21.612 ;
			RECT	177.311 21.548 177.343 21.612 ;
			RECT	177.479 21.548 177.511 21.612 ;
			RECT	177.647 21.548 177.679 21.612 ;
			RECT	177.815 21.548 177.847 21.612 ;
			RECT	177.983 21.548 178.015 21.612 ;
			RECT	178.151 21.548 178.183 21.612 ;
			RECT	178.319 21.548 178.351 21.612 ;
			RECT	178.487 21.548 178.519 21.612 ;
			RECT	178.655 21.548 178.687 21.612 ;
			RECT	178.823 21.548 178.855 21.612 ;
			RECT	178.991 21.548 179.023 21.612 ;
			RECT	179.159 21.548 179.191 21.612 ;
			RECT	179.327 21.548 179.359 21.612 ;
			RECT	179.495 21.548 179.527 21.612 ;
			RECT	179.663 21.548 179.695 21.612 ;
			RECT	179.831 21.548 179.863 21.612 ;
			RECT	179.999 21.548 180.031 21.612 ;
			RECT	180.167 21.548 180.199 21.612 ;
			RECT	180.335 21.548 180.367 21.612 ;
			RECT	180.503 21.548 180.535 21.612 ;
			RECT	180.671 21.548 180.703 21.612 ;
			RECT	180.839 21.548 180.871 21.612 ;
			RECT	181.007 21.548 181.039 21.612 ;
			RECT	181.175 21.548 181.207 21.612 ;
			RECT	181.343 21.548 181.375 21.612 ;
			RECT	181.511 21.548 181.543 21.612 ;
			RECT	181.679 21.548 181.711 21.612 ;
			RECT	181.847 21.548 181.879 21.612 ;
			RECT	182.015 21.548 182.047 21.612 ;
			RECT	182.183 21.548 182.215 21.612 ;
			RECT	182.351 21.548 182.383 21.612 ;
			RECT	182.519 21.548 182.551 21.612 ;
			RECT	182.687 21.548 182.719 21.612 ;
			RECT	182.855 21.548 182.887 21.612 ;
			RECT	183.023 21.548 183.055 21.612 ;
			RECT	183.191 21.548 183.223 21.612 ;
			RECT	183.359 21.548 183.391 21.612 ;
			RECT	183.527 21.548 183.559 21.612 ;
			RECT	183.695 21.548 183.727 21.612 ;
			RECT	183.863 21.548 183.895 21.612 ;
			RECT	184.031 21.548 184.063 21.612 ;
			RECT	184.199 21.548 184.231 21.612 ;
			RECT	184.367 21.548 184.399 21.612 ;
			RECT	184.535 21.548 184.567 21.612 ;
			RECT	184.703 21.548 184.735 21.612 ;
			RECT	184.871 21.548 184.903 21.612 ;
			RECT	185.039 21.548 185.071 21.612 ;
			RECT	185.207 21.548 185.239 21.612 ;
			RECT	185.375 21.548 185.407 21.612 ;
			RECT	185.543 21.548 185.575 21.612 ;
			RECT	185.711 21.548 185.743 21.612 ;
			RECT	185.879 21.548 185.911 21.612 ;
			RECT	186.047 21.548 186.079 21.612 ;
			RECT	186.215 21.548 186.247 21.612 ;
			RECT	186.383 21.548 186.415 21.612 ;
			RECT	186.551 21.548 186.583 21.612 ;
			RECT	186.719 21.548 186.751 21.612 ;
			RECT	186.887 21.548 186.919 21.612 ;
			RECT	187.055 21.548 187.087 21.612 ;
			RECT	187.223 21.548 187.255 21.612 ;
			RECT	187.391 21.548 187.423 21.612 ;
			RECT	187.559 21.548 187.591 21.612 ;
			RECT	187.727 21.548 187.759 21.612 ;
			RECT	187.895 21.548 187.927 21.612 ;
			RECT	188.063 21.548 188.095 21.612 ;
			RECT	188.231 21.548 188.263 21.612 ;
			RECT	188.399 21.548 188.431 21.612 ;
			RECT	188.567 21.548 188.599 21.612 ;
			RECT	188.735 21.548 188.767 21.612 ;
			RECT	188.903 21.548 188.935 21.612 ;
			RECT	189.071 21.548 189.103 21.612 ;
			RECT	189.239 21.548 189.271 21.612 ;
			RECT	189.407 21.548 189.439 21.612 ;
			RECT	189.575 21.548 189.607 21.612 ;
			RECT	189.743 21.548 189.775 21.612 ;
			RECT	189.911 21.548 189.943 21.612 ;
			RECT	190.079 21.548 190.111 21.612 ;
			RECT	190.247 21.548 190.279 21.612 ;
			RECT	190.415 21.548 190.447 21.612 ;
			RECT	190.583 21.548 190.615 21.612 ;
			RECT	190.751 21.548 190.783 21.612 ;
			RECT	190.919 21.548 190.951 21.612 ;
			RECT	191.087 21.548 191.119 21.612 ;
			RECT	191.255 21.548 191.287 21.612 ;
			RECT	191.423 21.548 191.455 21.612 ;
			RECT	191.591 21.548 191.623 21.612 ;
			RECT	191.759 21.548 191.791 21.612 ;
			RECT	191.927 21.548 191.959 21.612 ;
			RECT	192.095 21.548 192.127 21.612 ;
			RECT	192.263 21.548 192.295 21.612 ;
			RECT	192.431 21.548 192.463 21.612 ;
			RECT	192.599 21.548 192.631 21.612 ;
			RECT	192.767 21.548 192.799 21.612 ;
			RECT	192.935 21.548 192.967 21.612 ;
			RECT	193.103 21.548 193.135 21.612 ;
			RECT	193.271 21.548 193.303 21.612 ;
			RECT	193.439 21.548 193.471 21.612 ;
			RECT	193.607 21.548 193.639 21.612 ;
			RECT	193.775 21.548 193.807 21.612 ;
			RECT	193.943 21.548 193.975 21.612 ;
			RECT	194.111 21.548 194.143 21.612 ;
			RECT	194.279 21.548 194.311 21.612 ;
			RECT	194.447 21.548 194.479 21.612 ;
			RECT	194.615 21.548 194.647 21.612 ;
			RECT	194.783 21.548 194.815 21.612 ;
			RECT	194.951 21.548 194.983 21.612 ;
			RECT	195.119 21.548 195.151 21.612 ;
			RECT	195.287 21.548 195.319 21.612 ;
			RECT	195.455 21.548 195.487 21.612 ;
			RECT	195.623 21.548 195.655 21.612 ;
			RECT	195.791 21.548 195.823 21.612 ;
			RECT	195.959 21.548 195.991 21.612 ;
			RECT	196.127 21.548 196.159 21.612 ;
			RECT	196.295 21.548 196.327 21.612 ;
			RECT	196.463 21.548 196.495 21.612 ;
			RECT	196.631 21.548 196.663 21.612 ;
			RECT	196.799 21.548 196.831 21.612 ;
			RECT	196.967 21.548 196.999 21.612 ;
			RECT	197.135 21.548 197.167 21.612 ;
			RECT	197.303 21.548 197.335 21.612 ;
			RECT	197.471 21.548 197.503 21.612 ;
			RECT	197.639 21.548 197.671 21.612 ;
			RECT	197.807 21.548 197.839 21.612 ;
			RECT	197.975 21.548 198.007 21.612 ;
			RECT	198.143 21.548 198.175 21.612 ;
			RECT	198.311 21.548 198.343 21.612 ;
			RECT	198.479 21.548 198.511 21.612 ;
			RECT	198.647 21.548 198.679 21.612 ;
			RECT	198.815 21.548 198.847 21.612 ;
			RECT	198.983 21.548 199.015 21.612 ;
			RECT	199.151 21.548 199.183 21.612 ;
			RECT	199.319 21.548 199.351 21.612 ;
			RECT	199.487 21.548 199.519 21.612 ;
			RECT	199.655 21.548 199.687 21.612 ;
			RECT	199.823 21.548 199.855 21.612 ;
			RECT	199.991 21.548 200.023 21.612 ;
			RECT	200.121 21.564 200.153 21.596 ;
			RECT	200.243 21.569 200.275 21.601 ;
			RECT	200.373 21.548 200.405 21.612 ;
			RECT	200.9 21.548 200.932 21.612 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 19.6 201.665 19.72 ;
			LAYER	J3 ;
			RECT	0.755 19.628 0.787 19.692 ;
			RECT	1.645 19.628 1.709 19.692 ;
			RECT	2.323 19.628 2.387 19.692 ;
			RECT	3.438 19.628 3.47 19.692 ;
			RECT	3.585 19.628 3.617 19.692 ;
			RECT	4.195 19.628 4.227 19.692 ;
			RECT	4.72 19.628 4.752 19.692 ;
			RECT	4.944 19.628 5.008 19.692 ;
			RECT	5.267 19.628 5.299 19.692 ;
			RECT	5.797 19.628 5.829 19.692 ;
			RECT	5.927 19.649 5.959 19.681 ;
			RECT	6.049 19.644 6.081 19.676 ;
			RECT	6.179 19.628 6.211 19.692 ;
			RECT	6.347 19.628 6.379 19.692 ;
			RECT	6.515 19.628 6.547 19.692 ;
			RECT	6.683 19.628 6.715 19.692 ;
			RECT	6.851 19.628 6.883 19.692 ;
			RECT	7.019 19.628 7.051 19.692 ;
			RECT	7.187 19.628 7.219 19.692 ;
			RECT	7.355 19.628 7.387 19.692 ;
			RECT	7.523 19.628 7.555 19.692 ;
			RECT	7.691 19.628 7.723 19.692 ;
			RECT	7.859 19.628 7.891 19.692 ;
			RECT	8.027 19.628 8.059 19.692 ;
			RECT	8.195 19.628 8.227 19.692 ;
			RECT	8.363 19.628 8.395 19.692 ;
			RECT	8.531 19.628 8.563 19.692 ;
			RECT	8.699 19.628 8.731 19.692 ;
			RECT	8.867 19.628 8.899 19.692 ;
			RECT	9.035 19.628 9.067 19.692 ;
			RECT	9.203 19.628 9.235 19.692 ;
			RECT	9.371 19.628 9.403 19.692 ;
			RECT	9.539 19.628 9.571 19.692 ;
			RECT	9.707 19.628 9.739 19.692 ;
			RECT	9.875 19.628 9.907 19.692 ;
			RECT	10.043 19.628 10.075 19.692 ;
			RECT	10.211 19.628 10.243 19.692 ;
			RECT	10.379 19.628 10.411 19.692 ;
			RECT	10.547 19.628 10.579 19.692 ;
			RECT	10.715 19.628 10.747 19.692 ;
			RECT	10.883 19.628 10.915 19.692 ;
			RECT	11.051 19.628 11.083 19.692 ;
			RECT	11.219 19.628 11.251 19.692 ;
			RECT	11.387 19.628 11.419 19.692 ;
			RECT	11.555 19.628 11.587 19.692 ;
			RECT	11.723 19.628 11.755 19.692 ;
			RECT	11.891 19.628 11.923 19.692 ;
			RECT	12.059 19.628 12.091 19.692 ;
			RECT	12.227 19.628 12.259 19.692 ;
			RECT	12.395 19.628 12.427 19.692 ;
			RECT	12.563 19.628 12.595 19.692 ;
			RECT	12.731 19.628 12.763 19.692 ;
			RECT	12.899 19.628 12.931 19.692 ;
			RECT	13.067 19.628 13.099 19.692 ;
			RECT	13.235 19.628 13.267 19.692 ;
			RECT	13.403 19.628 13.435 19.692 ;
			RECT	13.571 19.628 13.603 19.692 ;
			RECT	13.739 19.628 13.771 19.692 ;
			RECT	13.907 19.628 13.939 19.692 ;
			RECT	14.075 19.628 14.107 19.692 ;
			RECT	14.243 19.628 14.275 19.692 ;
			RECT	14.411 19.628 14.443 19.692 ;
			RECT	14.579 19.628 14.611 19.692 ;
			RECT	14.747 19.628 14.779 19.692 ;
			RECT	14.915 19.628 14.947 19.692 ;
			RECT	15.083 19.628 15.115 19.692 ;
			RECT	15.251 19.628 15.283 19.692 ;
			RECT	15.419 19.628 15.451 19.692 ;
			RECT	15.587 19.628 15.619 19.692 ;
			RECT	15.755 19.628 15.787 19.692 ;
			RECT	15.923 19.628 15.955 19.692 ;
			RECT	16.091 19.628 16.123 19.692 ;
			RECT	16.259 19.628 16.291 19.692 ;
			RECT	16.427 19.628 16.459 19.692 ;
			RECT	16.595 19.628 16.627 19.692 ;
			RECT	16.763 19.628 16.795 19.692 ;
			RECT	16.931 19.628 16.963 19.692 ;
			RECT	17.099 19.628 17.131 19.692 ;
			RECT	17.267 19.628 17.299 19.692 ;
			RECT	17.435 19.628 17.467 19.692 ;
			RECT	17.603 19.628 17.635 19.692 ;
			RECT	17.771 19.628 17.803 19.692 ;
			RECT	17.939 19.628 17.971 19.692 ;
			RECT	18.107 19.628 18.139 19.692 ;
			RECT	18.275 19.628 18.307 19.692 ;
			RECT	18.443 19.628 18.475 19.692 ;
			RECT	18.611 19.628 18.643 19.692 ;
			RECT	18.779 19.628 18.811 19.692 ;
			RECT	18.947 19.628 18.979 19.692 ;
			RECT	19.115 19.628 19.147 19.692 ;
			RECT	19.283 19.628 19.315 19.692 ;
			RECT	19.451 19.628 19.483 19.692 ;
			RECT	19.619 19.628 19.651 19.692 ;
			RECT	19.787 19.628 19.819 19.692 ;
			RECT	19.955 19.628 19.987 19.692 ;
			RECT	20.123 19.628 20.155 19.692 ;
			RECT	20.291 19.628 20.323 19.692 ;
			RECT	20.459 19.628 20.491 19.692 ;
			RECT	20.627 19.628 20.659 19.692 ;
			RECT	20.795 19.628 20.827 19.692 ;
			RECT	20.963 19.628 20.995 19.692 ;
			RECT	21.131 19.628 21.163 19.692 ;
			RECT	21.299 19.628 21.331 19.692 ;
			RECT	21.467 19.628 21.499 19.692 ;
			RECT	21.635 19.628 21.667 19.692 ;
			RECT	21.803 19.628 21.835 19.692 ;
			RECT	21.971 19.628 22.003 19.692 ;
			RECT	22.139 19.628 22.171 19.692 ;
			RECT	22.307 19.628 22.339 19.692 ;
			RECT	22.475 19.628 22.507 19.692 ;
			RECT	22.643 19.628 22.675 19.692 ;
			RECT	22.811 19.628 22.843 19.692 ;
			RECT	22.979 19.628 23.011 19.692 ;
			RECT	23.147 19.628 23.179 19.692 ;
			RECT	23.315 19.628 23.347 19.692 ;
			RECT	23.483 19.628 23.515 19.692 ;
			RECT	23.651 19.628 23.683 19.692 ;
			RECT	23.819 19.628 23.851 19.692 ;
			RECT	23.987 19.628 24.019 19.692 ;
			RECT	24.155 19.628 24.187 19.692 ;
			RECT	24.323 19.628 24.355 19.692 ;
			RECT	24.491 19.628 24.523 19.692 ;
			RECT	24.659 19.628 24.691 19.692 ;
			RECT	24.827 19.628 24.859 19.692 ;
			RECT	24.995 19.628 25.027 19.692 ;
			RECT	25.163 19.628 25.195 19.692 ;
			RECT	25.331 19.628 25.363 19.692 ;
			RECT	25.499 19.628 25.531 19.692 ;
			RECT	25.667 19.628 25.699 19.692 ;
			RECT	25.835 19.628 25.867 19.692 ;
			RECT	26.003 19.628 26.035 19.692 ;
			RECT	26.171 19.628 26.203 19.692 ;
			RECT	26.339 19.628 26.371 19.692 ;
			RECT	26.507 19.628 26.539 19.692 ;
			RECT	26.675 19.628 26.707 19.692 ;
			RECT	26.843 19.628 26.875 19.692 ;
			RECT	27.011 19.628 27.043 19.692 ;
			RECT	27.179 19.628 27.211 19.692 ;
			RECT	27.347 19.628 27.379 19.692 ;
			RECT	27.515 19.628 27.547 19.692 ;
			RECT	27.683 19.628 27.715 19.692 ;
			RECT	27.851 19.628 27.883 19.692 ;
			RECT	28.019 19.628 28.051 19.692 ;
			RECT	28.187 19.628 28.219 19.692 ;
			RECT	28.355 19.628 28.387 19.692 ;
			RECT	28.523 19.628 28.555 19.692 ;
			RECT	28.691 19.628 28.723 19.692 ;
			RECT	28.859 19.628 28.891 19.692 ;
			RECT	29.027 19.628 29.059 19.692 ;
			RECT	29.195 19.628 29.227 19.692 ;
			RECT	29.363 19.628 29.395 19.692 ;
			RECT	29.531 19.628 29.563 19.692 ;
			RECT	29.699 19.628 29.731 19.692 ;
			RECT	29.867 19.628 29.899 19.692 ;
			RECT	30.035 19.628 30.067 19.692 ;
			RECT	30.203 19.628 30.235 19.692 ;
			RECT	30.371 19.628 30.403 19.692 ;
			RECT	30.539 19.628 30.571 19.692 ;
			RECT	30.707 19.628 30.739 19.692 ;
			RECT	30.875 19.628 30.907 19.692 ;
			RECT	31.043 19.628 31.075 19.692 ;
			RECT	31.211 19.628 31.243 19.692 ;
			RECT	31.379 19.628 31.411 19.692 ;
			RECT	31.547 19.628 31.579 19.692 ;
			RECT	31.715 19.628 31.747 19.692 ;
			RECT	31.883 19.628 31.915 19.692 ;
			RECT	32.051 19.628 32.083 19.692 ;
			RECT	32.219 19.628 32.251 19.692 ;
			RECT	32.387 19.628 32.419 19.692 ;
			RECT	32.555 19.628 32.587 19.692 ;
			RECT	32.723 19.628 32.755 19.692 ;
			RECT	32.891 19.628 32.923 19.692 ;
			RECT	33.059 19.628 33.091 19.692 ;
			RECT	33.227 19.628 33.259 19.692 ;
			RECT	33.395 19.628 33.427 19.692 ;
			RECT	33.563 19.628 33.595 19.692 ;
			RECT	33.731 19.628 33.763 19.692 ;
			RECT	33.899 19.628 33.931 19.692 ;
			RECT	34.067 19.628 34.099 19.692 ;
			RECT	34.235 19.628 34.267 19.692 ;
			RECT	34.403 19.628 34.435 19.692 ;
			RECT	34.571 19.628 34.603 19.692 ;
			RECT	34.739 19.628 34.771 19.692 ;
			RECT	34.907 19.628 34.939 19.692 ;
			RECT	35.075 19.628 35.107 19.692 ;
			RECT	35.243 19.628 35.275 19.692 ;
			RECT	35.411 19.628 35.443 19.692 ;
			RECT	35.579 19.628 35.611 19.692 ;
			RECT	35.747 19.628 35.779 19.692 ;
			RECT	35.915 19.628 35.947 19.692 ;
			RECT	36.083 19.628 36.115 19.692 ;
			RECT	36.251 19.628 36.283 19.692 ;
			RECT	36.419 19.628 36.451 19.692 ;
			RECT	36.587 19.628 36.619 19.692 ;
			RECT	36.755 19.628 36.787 19.692 ;
			RECT	36.923 19.628 36.955 19.692 ;
			RECT	37.091 19.628 37.123 19.692 ;
			RECT	37.259 19.628 37.291 19.692 ;
			RECT	37.427 19.628 37.459 19.692 ;
			RECT	37.595 19.628 37.627 19.692 ;
			RECT	37.763 19.628 37.795 19.692 ;
			RECT	37.931 19.628 37.963 19.692 ;
			RECT	38.099 19.628 38.131 19.692 ;
			RECT	38.267 19.628 38.299 19.692 ;
			RECT	38.435 19.628 38.467 19.692 ;
			RECT	38.603 19.628 38.635 19.692 ;
			RECT	38.771 19.628 38.803 19.692 ;
			RECT	38.939 19.628 38.971 19.692 ;
			RECT	39.107 19.628 39.139 19.692 ;
			RECT	39.275 19.628 39.307 19.692 ;
			RECT	39.443 19.628 39.475 19.692 ;
			RECT	39.611 19.628 39.643 19.692 ;
			RECT	39.779 19.628 39.811 19.692 ;
			RECT	39.947 19.628 39.979 19.692 ;
			RECT	40.115 19.628 40.147 19.692 ;
			RECT	40.283 19.628 40.315 19.692 ;
			RECT	40.451 19.628 40.483 19.692 ;
			RECT	40.619 19.628 40.651 19.692 ;
			RECT	40.787 19.628 40.819 19.692 ;
			RECT	40.955 19.628 40.987 19.692 ;
			RECT	41.123 19.628 41.155 19.692 ;
			RECT	41.291 19.628 41.323 19.692 ;
			RECT	41.459 19.628 41.491 19.692 ;
			RECT	41.627 19.628 41.659 19.692 ;
			RECT	41.795 19.628 41.827 19.692 ;
			RECT	41.963 19.628 41.995 19.692 ;
			RECT	42.131 19.628 42.163 19.692 ;
			RECT	42.299 19.628 42.331 19.692 ;
			RECT	42.467 19.628 42.499 19.692 ;
			RECT	42.635 19.628 42.667 19.692 ;
			RECT	42.803 19.628 42.835 19.692 ;
			RECT	42.971 19.628 43.003 19.692 ;
			RECT	43.139 19.628 43.171 19.692 ;
			RECT	43.307 19.628 43.339 19.692 ;
			RECT	43.475 19.628 43.507 19.692 ;
			RECT	43.643 19.628 43.675 19.692 ;
			RECT	43.811 19.628 43.843 19.692 ;
			RECT	43.979 19.628 44.011 19.692 ;
			RECT	44.147 19.628 44.179 19.692 ;
			RECT	44.315 19.628 44.347 19.692 ;
			RECT	44.483 19.628 44.515 19.692 ;
			RECT	44.651 19.628 44.683 19.692 ;
			RECT	44.819 19.628 44.851 19.692 ;
			RECT	44.987 19.628 45.019 19.692 ;
			RECT	45.155 19.628 45.187 19.692 ;
			RECT	45.323 19.628 45.355 19.692 ;
			RECT	45.491 19.628 45.523 19.692 ;
			RECT	45.659 19.628 45.691 19.692 ;
			RECT	45.827 19.628 45.859 19.692 ;
			RECT	45.995 19.628 46.027 19.692 ;
			RECT	46.163 19.628 46.195 19.692 ;
			RECT	46.331 19.628 46.363 19.692 ;
			RECT	46.499 19.628 46.531 19.692 ;
			RECT	46.667 19.628 46.699 19.692 ;
			RECT	46.835 19.628 46.867 19.692 ;
			RECT	47.003 19.628 47.035 19.692 ;
			RECT	47.171 19.628 47.203 19.692 ;
			RECT	47.339 19.628 47.371 19.692 ;
			RECT	47.507 19.628 47.539 19.692 ;
			RECT	47.675 19.628 47.707 19.692 ;
			RECT	47.843 19.628 47.875 19.692 ;
			RECT	48.011 19.628 48.043 19.692 ;
			RECT	48.179 19.628 48.211 19.692 ;
			RECT	48.347 19.628 48.379 19.692 ;
			RECT	48.515 19.628 48.547 19.692 ;
			RECT	48.683 19.628 48.715 19.692 ;
			RECT	48.851 19.628 48.883 19.692 ;
			RECT	49.019 19.628 49.051 19.692 ;
			RECT	49.187 19.628 49.219 19.692 ;
			RECT	49.318 19.644 49.35 19.676 ;
			RECT	49.439 19.644 49.471 19.676 ;
			RECT	49.569 19.628 49.601 19.692 ;
			RECT	51.881 19.628 51.913 19.692 ;
			RECT	53.132 19.628 53.196 19.692 ;
			RECT	53.812 19.628 53.844 19.692 ;
			RECT	54.251 19.628 54.283 19.692 ;
			RECT	55.562 19.628 55.626 19.692 ;
			RECT	58.603 19.628 58.635 19.692 ;
			RECT	58.733 19.644 58.765 19.676 ;
			RECT	58.854 19.644 58.886 19.676 ;
			RECT	58.985 19.628 59.017 19.692 ;
			RECT	59.153 19.628 59.185 19.692 ;
			RECT	59.321 19.628 59.353 19.692 ;
			RECT	59.489 19.628 59.521 19.692 ;
			RECT	59.657 19.628 59.689 19.692 ;
			RECT	59.825 19.628 59.857 19.692 ;
			RECT	59.993 19.628 60.025 19.692 ;
			RECT	60.161 19.628 60.193 19.692 ;
			RECT	60.329 19.628 60.361 19.692 ;
			RECT	60.497 19.628 60.529 19.692 ;
			RECT	60.665 19.628 60.697 19.692 ;
			RECT	60.833 19.628 60.865 19.692 ;
			RECT	61.001 19.628 61.033 19.692 ;
			RECT	61.169 19.628 61.201 19.692 ;
			RECT	61.337 19.628 61.369 19.692 ;
			RECT	61.505 19.628 61.537 19.692 ;
			RECT	61.673 19.628 61.705 19.692 ;
			RECT	61.841 19.628 61.873 19.692 ;
			RECT	62.009 19.628 62.041 19.692 ;
			RECT	62.177 19.628 62.209 19.692 ;
			RECT	62.345 19.628 62.377 19.692 ;
			RECT	62.513 19.628 62.545 19.692 ;
			RECT	62.681 19.628 62.713 19.692 ;
			RECT	62.849 19.628 62.881 19.692 ;
			RECT	63.017 19.628 63.049 19.692 ;
			RECT	63.185 19.628 63.217 19.692 ;
			RECT	63.353 19.628 63.385 19.692 ;
			RECT	63.521 19.628 63.553 19.692 ;
			RECT	63.689 19.628 63.721 19.692 ;
			RECT	63.857 19.628 63.889 19.692 ;
			RECT	64.025 19.628 64.057 19.692 ;
			RECT	64.193 19.628 64.225 19.692 ;
			RECT	64.361 19.628 64.393 19.692 ;
			RECT	64.529 19.628 64.561 19.692 ;
			RECT	64.697 19.628 64.729 19.692 ;
			RECT	64.865 19.628 64.897 19.692 ;
			RECT	65.033 19.628 65.065 19.692 ;
			RECT	65.201 19.628 65.233 19.692 ;
			RECT	65.369 19.628 65.401 19.692 ;
			RECT	65.537 19.628 65.569 19.692 ;
			RECT	65.705 19.628 65.737 19.692 ;
			RECT	65.873 19.628 65.905 19.692 ;
			RECT	66.041 19.628 66.073 19.692 ;
			RECT	66.209 19.628 66.241 19.692 ;
			RECT	66.377 19.628 66.409 19.692 ;
			RECT	66.545 19.628 66.577 19.692 ;
			RECT	66.713 19.628 66.745 19.692 ;
			RECT	66.881 19.628 66.913 19.692 ;
			RECT	67.049 19.628 67.081 19.692 ;
			RECT	67.217 19.628 67.249 19.692 ;
			RECT	67.385 19.628 67.417 19.692 ;
			RECT	67.553 19.628 67.585 19.692 ;
			RECT	67.721 19.628 67.753 19.692 ;
			RECT	67.889 19.628 67.921 19.692 ;
			RECT	68.057 19.628 68.089 19.692 ;
			RECT	68.225 19.628 68.257 19.692 ;
			RECT	68.393 19.628 68.425 19.692 ;
			RECT	68.561 19.628 68.593 19.692 ;
			RECT	68.729 19.628 68.761 19.692 ;
			RECT	68.897 19.628 68.929 19.692 ;
			RECT	69.065 19.628 69.097 19.692 ;
			RECT	69.233 19.628 69.265 19.692 ;
			RECT	69.401 19.628 69.433 19.692 ;
			RECT	69.569 19.628 69.601 19.692 ;
			RECT	69.737 19.628 69.769 19.692 ;
			RECT	69.905 19.628 69.937 19.692 ;
			RECT	70.073 19.628 70.105 19.692 ;
			RECT	70.241 19.628 70.273 19.692 ;
			RECT	70.409 19.628 70.441 19.692 ;
			RECT	70.577 19.628 70.609 19.692 ;
			RECT	70.745 19.628 70.777 19.692 ;
			RECT	70.913 19.628 70.945 19.692 ;
			RECT	71.081 19.628 71.113 19.692 ;
			RECT	71.249 19.628 71.281 19.692 ;
			RECT	71.417 19.628 71.449 19.692 ;
			RECT	71.585 19.628 71.617 19.692 ;
			RECT	71.753 19.628 71.785 19.692 ;
			RECT	71.921 19.628 71.953 19.692 ;
			RECT	72.089 19.628 72.121 19.692 ;
			RECT	72.257 19.628 72.289 19.692 ;
			RECT	72.425 19.628 72.457 19.692 ;
			RECT	72.593 19.628 72.625 19.692 ;
			RECT	72.761 19.628 72.793 19.692 ;
			RECT	72.929 19.628 72.961 19.692 ;
			RECT	73.097 19.628 73.129 19.692 ;
			RECT	73.265 19.628 73.297 19.692 ;
			RECT	73.433 19.628 73.465 19.692 ;
			RECT	73.601 19.628 73.633 19.692 ;
			RECT	73.769 19.628 73.801 19.692 ;
			RECT	73.937 19.628 73.969 19.692 ;
			RECT	74.105 19.628 74.137 19.692 ;
			RECT	74.273 19.628 74.305 19.692 ;
			RECT	74.441 19.628 74.473 19.692 ;
			RECT	74.609 19.628 74.641 19.692 ;
			RECT	74.777 19.628 74.809 19.692 ;
			RECT	74.945 19.628 74.977 19.692 ;
			RECT	75.113 19.628 75.145 19.692 ;
			RECT	75.281 19.628 75.313 19.692 ;
			RECT	75.449 19.628 75.481 19.692 ;
			RECT	75.617 19.628 75.649 19.692 ;
			RECT	75.785 19.628 75.817 19.692 ;
			RECT	75.953 19.628 75.985 19.692 ;
			RECT	76.121 19.628 76.153 19.692 ;
			RECT	76.289 19.628 76.321 19.692 ;
			RECT	76.457 19.628 76.489 19.692 ;
			RECT	76.625 19.628 76.657 19.692 ;
			RECT	76.793 19.628 76.825 19.692 ;
			RECT	76.961 19.628 76.993 19.692 ;
			RECT	77.129 19.628 77.161 19.692 ;
			RECT	77.297 19.628 77.329 19.692 ;
			RECT	77.465 19.628 77.497 19.692 ;
			RECT	77.633 19.628 77.665 19.692 ;
			RECT	77.801 19.628 77.833 19.692 ;
			RECT	77.969 19.628 78.001 19.692 ;
			RECT	78.137 19.628 78.169 19.692 ;
			RECT	78.305 19.628 78.337 19.692 ;
			RECT	78.473 19.628 78.505 19.692 ;
			RECT	78.641 19.628 78.673 19.692 ;
			RECT	78.809 19.628 78.841 19.692 ;
			RECT	78.977 19.628 79.009 19.692 ;
			RECT	79.145 19.628 79.177 19.692 ;
			RECT	79.313 19.628 79.345 19.692 ;
			RECT	79.481 19.628 79.513 19.692 ;
			RECT	79.649 19.628 79.681 19.692 ;
			RECT	79.817 19.628 79.849 19.692 ;
			RECT	79.985 19.628 80.017 19.692 ;
			RECT	80.153 19.628 80.185 19.692 ;
			RECT	80.321 19.628 80.353 19.692 ;
			RECT	80.489 19.628 80.521 19.692 ;
			RECT	80.657 19.628 80.689 19.692 ;
			RECT	80.825 19.628 80.857 19.692 ;
			RECT	80.993 19.628 81.025 19.692 ;
			RECT	81.161 19.628 81.193 19.692 ;
			RECT	81.329 19.628 81.361 19.692 ;
			RECT	81.497 19.628 81.529 19.692 ;
			RECT	81.665 19.628 81.697 19.692 ;
			RECT	81.833 19.628 81.865 19.692 ;
			RECT	82.001 19.628 82.033 19.692 ;
			RECT	82.169 19.628 82.201 19.692 ;
			RECT	82.337 19.628 82.369 19.692 ;
			RECT	82.505 19.628 82.537 19.692 ;
			RECT	82.673 19.628 82.705 19.692 ;
			RECT	82.841 19.628 82.873 19.692 ;
			RECT	83.009 19.628 83.041 19.692 ;
			RECT	83.177 19.628 83.209 19.692 ;
			RECT	83.345 19.628 83.377 19.692 ;
			RECT	83.513 19.628 83.545 19.692 ;
			RECT	83.681 19.628 83.713 19.692 ;
			RECT	83.849 19.628 83.881 19.692 ;
			RECT	84.017 19.628 84.049 19.692 ;
			RECT	84.185 19.628 84.217 19.692 ;
			RECT	84.353 19.628 84.385 19.692 ;
			RECT	84.521 19.628 84.553 19.692 ;
			RECT	84.689 19.628 84.721 19.692 ;
			RECT	84.857 19.628 84.889 19.692 ;
			RECT	85.025 19.628 85.057 19.692 ;
			RECT	85.193 19.628 85.225 19.692 ;
			RECT	85.361 19.628 85.393 19.692 ;
			RECT	85.529 19.628 85.561 19.692 ;
			RECT	85.697 19.628 85.729 19.692 ;
			RECT	85.865 19.628 85.897 19.692 ;
			RECT	86.033 19.628 86.065 19.692 ;
			RECT	86.201 19.628 86.233 19.692 ;
			RECT	86.369 19.628 86.401 19.692 ;
			RECT	86.537 19.628 86.569 19.692 ;
			RECT	86.705 19.628 86.737 19.692 ;
			RECT	86.873 19.628 86.905 19.692 ;
			RECT	87.041 19.628 87.073 19.692 ;
			RECT	87.209 19.628 87.241 19.692 ;
			RECT	87.377 19.628 87.409 19.692 ;
			RECT	87.545 19.628 87.577 19.692 ;
			RECT	87.713 19.628 87.745 19.692 ;
			RECT	87.881 19.628 87.913 19.692 ;
			RECT	88.049 19.628 88.081 19.692 ;
			RECT	88.217 19.628 88.249 19.692 ;
			RECT	88.385 19.628 88.417 19.692 ;
			RECT	88.553 19.628 88.585 19.692 ;
			RECT	88.721 19.628 88.753 19.692 ;
			RECT	88.889 19.628 88.921 19.692 ;
			RECT	89.057 19.628 89.089 19.692 ;
			RECT	89.225 19.628 89.257 19.692 ;
			RECT	89.393 19.628 89.425 19.692 ;
			RECT	89.561 19.628 89.593 19.692 ;
			RECT	89.729 19.628 89.761 19.692 ;
			RECT	89.897 19.628 89.929 19.692 ;
			RECT	90.065 19.628 90.097 19.692 ;
			RECT	90.233 19.628 90.265 19.692 ;
			RECT	90.401 19.628 90.433 19.692 ;
			RECT	90.569 19.628 90.601 19.692 ;
			RECT	90.737 19.628 90.769 19.692 ;
			RECT	90.905 19.628 90.937 19.692 ;
			RECT	91.073 19.628 91.105 19.692 ;
			RECT	91.241 19.628 91.273 19.692 ;
			RECT	91.409 19.628 91.441 19.692 ;
			RECT	91.577 19.628 91.609 19.692 ;
			RECT	91.745 19.628 91.777 19.692 ;
			RECT	91.913 19.628 91.945 19.692 ;
			RECT	92.081 19.628 92.113 19.692 ;
			RECT	92.249 19.628 92.281 19.692 ;
			RECT	92.417 19.628 92.449 19.692 ;
			RECT	92.585 19.628 92.617 19.692 ;
			RECT	92.753 19.628 92.785 19.692 ;
			RECT	92.921 19.628 92.953 19.692 ;
			RECT	93.089 19.628 93.121 19.692 ;
			RECT	93.257 19.628 93.289 19.692 ;
			RECT	93.425 19.628 93.457 19.692 ;
			RECT	93.593 19.628 93.625 19.692 ;
			RECT	93.761 19.628 93.793 19.692 ;
			RECT	93.929 19.628 93.961 19.692 ;
			RECT	94.097 19.628 94.129 19.692 ;
			RECT	94.265 19.628 94.297 19.692 ;
			RECT	94.433 19.628 94.465 19.692 ;
			RECT	94.601 19.628 94.633 19.692 ;
			RECT	94.769 19.628 94.801 19.692 ;
			RECT	94.937 19.628 94.969 19.692 ;
			RECT	95.105 19.628 95.137 19.692 ;
			RECT	95.273 19.628 95.305 19.692 ;
			RECT	95.441 19.628 95.473 19.692 ;
			RECT	95.609 19.628 95.641 19.692 ;
			RECT	95.777 19.628 95.809 19.692 ;
			RECT	95.945 19.628 95.977 19.692 ;
			RECT	96.113 19.628 96.145 19.692 ;
			RECT	96.281 19.628 96.313 19.692 ;
			RECT	96.449 19.628 96.481 19.692 ;
			RECT	96.617 19.628 96.649 19.692 ;
			RECT	96.785 19.628 96.817 19.692 ;
			RECT	96.953 19.628 96.985 19.692 ;
			RECT	97.121 19.628 97.153 19.692 ;
			RECT	97.289 19.628 97.321 19.692 ;
			RECT	97.457 19.628 97.489 19.692 ;
			RECT	97.625 19.628 97.657 19.692 ;
			RECT	97.793 19.628 97.825 19.692 ;
			RECT	97.961 19.628 97.993 19.692 ;
			RECT	98.129 19.628 98.161 19.692 ;
			RECT	98.297 19.628 98.329 19.692 ;
			RECT	98.465 19.628 98.497 19.692 ;
			RECT	98.633 19.628 98.665 19.692 ;
			RECT	98.801 19.628 98.833 19.692 ;
			RECT	98.969 19.628 99.001 19.692 ;
			RECT	99.137 19.628 99.169 19.692 ;
			RECT	99.305 19.628 99.337 19.692 ;
			RECT	99.473 19.628 99.505 19.692 ;
			RECT	99.641 19.628 99.673 19.692 ;
			RECT	99.809 19.628 99.841 19.692 ;
			RECT	99.977 19.628 100.009 19.692 ;
			RECT	100.145 19.628 100.177 19.692 ;
			RECT	100.313 19.628 100.345 19.692 ;
			RECT	100.481 19.628 100.513 19.692 ;
			RECT	100.649 19.628 100.681 19.692 ;
			RECT	100.817 19.628 100.849 19.692 ;
			RECT	100.985 19.628 101.017 19.692 ;
			RECT	101.153 19.628 101.185 19.692 ;
			RECT	101.321 19.628 101.353 19.692 ;
			RECT	101.489 19.628 101.521 19.692 ;
			RECT	101.657 19.628 101.689 19.692 ;
			RECT	101.825 19.628 101.857 19.692 ;
			RECT	101.993 19.628 102.025 19.692 ;
			RECT	102.123 19.644 102.155 19.676 ;
			RECT	102.245 19.649 102.277 19.681 ;
			RECT	102.375 19.628 102.407 19.692 ;
			RECT	103.795 19.628 103.827 19.692 ;
			RECT	103.925 19.649 103.957 19.681 ;
			RECT	104.047 19.644 104.079 19.676 ;
			RECT	104.177 19.628 104.209 19.692 ;
			RECT	104.345 19.628 104.377 19.692 ;
			RECT	104.513 19.628 104.545 19.692 ;
			RECT	104.681 19.628 104.713 19.692 ;
			RECT	104.849 19.628 104.881 19.692 ;
			RECT	105.017 19.628 105.049 19.692 ;
			RECT	105.185 19.628 105.217 19.692 ;
			RECT	105.353 19.628 105.385 19.692 ;
			RECT	105.521 19.628 105.553 19.692 ;
			RECT	105.689 19.628 105.721 19.692 ;
			RECT	105.857 19.628 105.889 19.692 ;
			RECT	106.025 19.628 106.057 19.692 ;
			RECT	106.193 19.628 106.225 19.692 ;
			RECT	106.361 19.628 106.393 19.692 ;
			RECT	106.529 19.628 106.561 19.692 ;
			RECT	106.697 19.628 106.729 19.692 ;
			RECT	106.865 19.628 106.897 19.692 ;
			RECT	107.033 19.628 107.065 19.692 ;
			RECT	107.201 19.628 107.233 19.692 ;
			RECT	107.369 19.628 107.401 19.692 ;
			RECT	107.537 19.628 107.569 19.692 ;
			RECT	107.705 19.628 107.737 19.692 ;
			RECT	107.873 19.628 107.905 19.692 ;
			RECT	108.041 19.628 108.073 19.692 ;
			RECT	108.209 19.628 108.241 19.692 ;
			RECT	108.377 19.628 108.409 19.692 ;
			RECT	108.545 19.628 108.577 19.692 ;
			RECT	108.713 19.628 108.745 19.692 ;
			RECT	108.881 19.628 108.913 19.692 ;
			RECT	109.049 19.628 109.081 19.692 ;
			RECT	109.217 19.628 109.249 19.692 ;
			RECT	109.385 19.628 109.417 19.692 ;
			RECT	109.553 19.628 109.585 19.692 ;
			RECT	109.721 19.628 109.753 19.692 ;
			RECT	109.889 19.628 109.921 19.692 ;
			RECT	110.057 19.628 110.089 19.692 ;
			RECT	110.225 19.628 110.257 19.692 ;
			RECT	110.393 19.628 110.425 19.692 ;
			RECT	110.561 19.628 110.593 19.692 ;
			RECT	110.729 19.628 110.761 19.692 ;
			RECT	110.897 19.628 110.929 19.692 ;
			RECT	111.065 19.628 111.097 19.692 ;
			RECT	111.233 19.628 111.265 19.692 ;
			RECT	111.401 19.628 111.433 19.692 ;
			RECT	111.569 19.628 111.601 19.692 ;
			RECT	111.737 19.628 111.769 19.692 ;
			RECT	111.905 19.628 111.937 19.692 ;
			RECT	112.073 19.628 112.105 19.692 ;
			RECT	112.241 19.628 112.273 19.692 ;
			RECT	112.409 19.628 112.441 19.692 ;
			RECT	112.577 19.628 112.609 19.692 ;
			RECT	112.745 19.628 112.777 19.692 ;
			RECT	112.913 19.628 112.945 19.692 ;
			RECT	113.081 19.628 113.113 19.692 ;
			RECT	113.249 19.628 113.281 19.692 ;
			RECT	113.417 19.628 113.449 19.692 ;
			RECT	113.585 19.628 113.617 19.692 ;
			RECT	113.753 19.628 113.785 19.692 ;
			RECT	113.921 19.628 113.953 19.692 ;
			RECT	114.089 19.628 114.121 19.692 ;
			RECT	114.257 19.628 114.289 19.692 ;
			RECT	114.425 19.628 114.457 19.692 ;
			RECT	114.593 19.628 114.625 19.692 ;
			RECT	114.761 19.628 114.793 19.692 ;
			RECT	114.929 19.628 114.961 19.692 ;
			RECT	115.097 19.628 115.129 19.692 ;
			RECT	115.265 19.628 115.297 19.692 ;
			RECT	115.433 19.628 115.465 19.692 ;
			RECT	115.601 19.628 115.633 19.692 ;
			RECT	115.769 19.628 115.801 19.692 ;
			RECT	115.937 19.628 115.969 19.692 ;
			RECT	116.105 19.628 116.137 19.692 ;
			RECT	116.273 19.628 116.305 19.692 ;
			RECT	116.441 19.628 116.473 19.692 ;
			RECT	116.609 19.628 116.641 19.692 ;
			RECT	116.777 19.628 116.809 19.692 ;
			RECT	116.945 19.628 116.977 19.692 ;
			RECT	117.113 19.628 117.145 19.692 ;
			RECT	117.281 19.628 117.313 19.692 ;
			RECT	117.449 19.628 117.481 19.692 ;
			RECT	117.617 19.628 117.649 19.692 ;
			RECT	117.785 19.628 117.817 19.692 ;
			RECT	117.953 19.628 117.985 19.692 ;
			RECT	118.121 19.628 118.153 19.692 ;
			RECT	118.289 19.628 118.321 19.692 ;
			RECT	118.457 19.628 118.489 19.692 ;
			RECT	118.625 19.628 118.657 19.692 ;
			RECT	118.793 19.628 118.825 19.692 ;
			RECT	118.961 19.628 118.993 19.692 ;
			RECT	119.129 19.628 119.161 19.692 ;
			RECT	119.297 19.628 119.329 19.692 ;
			RECT	119.465 19.628 119.497 19.692 ;
			RECT	119.633 19.628 119.665 19.692 ;
			RECT	119.801 19.628 119.833 19.692 ;
			RECT	119.969 19.628 120.001 19.692 ;
			RECT	120.137 19.628 120.169 19.692 ;
			RECT	120.305 19.628 120.337 19.692 ;
			RECT	120.473 19.628 120.505 19.692 ;
			RECT	120.641 19.628 120.673 19.692 ;
			RECT	120.809 19.628 120.841 19.692 ;
			RECT	120.977 19.628 121.009 19.692 ;
			RECT	121.145 19.628 121.177 19.692 ;
			RECT	121.313 19.628 121.345 19.692 ;
			RECT	121.481 19.628 121.513 19.692 ;
			RECT	121.649 19.628 121.681 19.692 ;
			RECT	121.817 19.628 121.849 19.692 ;
			RECT	121.985 19.628 122.017 19.692 ;
			RECT	122.153 19.628 122.185 19.692 ;
			RECT	122.321 19.628 122.353 19.692 ;
			RECT	122.489 19.628 122.521 19.692 ;
			RECT	122.657 19.628 122.689 19.692 ;
			RECT	122.825 19.628 122.857 19.692 ;
			RECT	122.993 19.628 123.025 19.692 ;
			RECT	123.161 19.628 123.193 19.692 ;
			RECT	123.329 19.628 123.361 19.692 ;
			RECT	123.497 19.628 123.529 19.692 ;
			RECT	123.665 19.628 123.697 19.692 ;
			RECT	123.833 19.628 123.865 19.692 ;
			RECT	124.001 19.628 124.033 19.692 ;
			RECT	124.169 19.628 124.201 19.692 ;
			RECT	124.337 19.628 124.369 19.692 ;
			RECT	124.505 19.628 124.537 19.692 ;
			RECT	124.673 19.628 124.705 19.692 ;
			RECT	124.841 19.628 124.873 19.692 ;
			RECT	125.009 19.628 125.041 19.692 ;
			RECT	125.177 19.628 125.209 19.692 ;
			RECT	125.345 19.628 125.377 19.692 ;
			RECT	125.513 19.628 125.545 19.692 ;
			RECT	125.681 19.628 125.713 19.692 ;
			RECT	125.849 19.628 125.881 19.692 ;
			RECT	126.017 19.628 126.049 19.692 ;
			RECT	126.185 19.628 126.217 19.692 ;
			RECT	126.353 19.628 126.385 19.692 ;
			RECT	126.521 19.628 126.553 19.692 ;
			RECT	126.689 19.628 126.721 19.692 ;
			RECT	126.857 19.628 126.889 19.692 ;
			RECT	127.025 19.628 127.057 19.692 ;
			RECT	127.193 19.628 127.225 19.692 ;
			RECT	127.361 19.628 127.393 19.692 ;
			RECT	127.529 19.628 127.561 19.692 ;
			RECT	127.697 19.628 127.729 19.692 ;
			RECT	127.865 19.628 127.897 19.692 ;
			RECT	128.033 19.628 128.065 19.692 ;
			RECT	128.201 19.628 128.233 19.692 ;
			RECT	128.369 19.628 128.401 19.692 ;
			RECT	128.537 19.628 128.569 19.692 ;
			RECT	128.705 19.628 128.737 19.692 ;
			RECT	128.873 19.628 128.905 19.692 ;
			RECT	129.041 19.628 129.073 19.692 ;
			RECT	129.209 19.628 129.241 19.692 ;
			RECT	129.377 19.628 129.409 19.692 ;
			RECT	129.545 19.628 129.577 19.692 ;
			RECT	129.713 19.628 129.745 19.692 ;
			RECT	129.881 19.628 129.913 19.692 ;
			RECT	130.049 19.628 130.081 19.692 ;
			RECT	130.217 19.628 130.249 19.692 ;
			RECT	130.385 19.628 130.417 19.692 ;
			RECT	130.553 19.628 130.585 19.692 ;
			RECT	130.721 19.628 130.753 19.692 ;
			RECT	130.889 19.628 130.921 19.692 ;
			RECT	131.057 19.628 131.089 19.692 ;
			RECT	131.225 19.628 131.257 19.692 ;
			RECT	131.393 19.628 131.425 19.692 ;
			RECT	131.561 19.628 131.593 19.692 ;
			RECT	131.729 19.628 131.761 19.692 ;
			RECT	131.897 19.628 131.929 19.692 ;
			RECT	132.065 19.628 132.097 19.692 ;
			RECT	132.233 19.628 132.265 19.692 ;
			RECT	132.401 19.628 132.433 19.692 ;
			RECT	132.569 19.628 132.601 19.692 ;
			RECT	132.737 19.628 132.769 19.692 ;
			RECT	132.905 19.628 132.937 19.692 ;
			RECT	133.073 19.628 133.105 19.692 ;
			RECT	133.241 19.628 133.273 19.692 ;
			RECT	133.409 19.628 133.441 19.692 ;
			RECT	133.577 19.628 133.609 19.692 ;
			RECT	133.745 19.628 133.777 19.692 ;
			RECT	133.913 19.628 133.945 19.692 ;
			RECT	134.081 19.628 134.113 19.692 ;
			RECT	134.249 19.628 134.281 19.692 ;
			RECT	134.417 19.628 134.449 19.692 ;
			RECT	134.585 19.628 134.617 19.692 ;
			RECT	134.753 19.628 134.785 19.692 ;
			RECT	134.921 19.628 134.953 19.692 ;
			RECT	135.089 19.628 135.121 19.692 ;
			RECT	135.257 19.628 135.289 19.692 ;
			RECT	135.425 19.628 135.457 19.692 ;
			RECT	135.593 19.628 135.625 19.692 ;
			RECT	135.761 19.628 135.793 19.692 ;
			RECT	135.929 19.628 135.961 19.692 ;
			RECT	136.097 19.628 136.129 19.692 ;
			RECT	136.265 19.628 136.297 19.692 ;
			RECT	136.433 19.628 136.465 19.692 ;
			RECT	136.601 19.628 136.633 19.692 ;
			RECT	136.769 19.628 136.801 19.692 ;
			RECT	136.937 19.628 136.969 19.692 ;
			RECT	137.105 19.628 137.137 19.692 ;
			RECT	137.273 19.628 137.305 19.692 ;
			RECT	137.441 19.628 137.473 19.692 ;
			RECT	137.609 19.628 137.641 19.692 ;
			RECT	137.777 19.628 137.809 19.692 ;
			RECT	137.945 19.628 137.977 19.692 ;
			RECT	138.113 19.628 138.145 19.692 ;
			RECT	138.281 19.628 138.313 19.692 ;
			RECT	138.449 19.628 138.481 19.692 ;
			RECT	138.617 19.628 138.649 19.692 ;
			RECT	138.785 19.628 138.817 19.692 ;
			RECT	138.953 19.628 138.985 19.692 ;
			RECT	139.121 19.628 139.153 19.692 ;
			RECT	139.289 19.628 139.321 19.692 ;
			RECT	139.457 19.628 139.489 19.692 ;
			RECT	139.625 19.628 139.657 19.692 ;
			RECT	139.793 19.628 139.825 19.692 ;
			RECT	139.961 19.628 139.993 19.692 ;
			RECT	140.129 19.628 140.161 19.692 ;
			RECT	140.297 19.628 140.329 19.692 ;
			RECT	140.465 19.628 140.497 19.692 ;
			RECT	140.633 19.628 140.665 19.692 ;
			RECT	140.801 19.628 140.833 19.692 ;
			RECT	140.969 19.628 141.001 19.692 ;
			RECT	141.137 19.628 141.169 19.692 ;
			RECT	141.305 19.628 141.337 19.692 ;
			RECT	141.473 19.628 141.505 19.692 ;
			RECT	141.641 19.628 141.673 19.692 ;
			RECT	141.809 19.628 141.841 19.692 ;
			RECT	141.977 19.628 142.009 19.692 ;
			RECT	142.145 19.628 142.177 19.692 ;
			RECT	142.313 19.628 142.345 19.692 ;
			RECT	142.481 19.628 142.513 19.692 ;
			RECT	142.649 19.628 142.681 19.692 ;
			RECT	142.817 19.628 142.849 19.692 ;
			RECT	142.985 19.628 143.017 19.692 ;
			RECT	143.153 19.628 143.185 19.692 ;
			RECT	143.321 19.628 143.353 19.692 ;
			RECT	143.489 19.628 143.521 19.692 ;
			RECT	143.657 19.628 143.689 19.692 ;
			RECT	143.825 19.628 143.857 19.692 ;
			RECT	143.993 19.628 144.025 19.692 ;
			RECT	144.161 19.628 144.193 19.692 ;
			RECT	144.329 19.628 144.361 19.692 ;
			RECT	144.497 19.628 144.529 19.692 ;
			RECT	144.665 19.628 144.697 19.692 ;
			RECT	144.833 19.628 144.865 19.692 ;
			RECT	145.001 19.628 145.033 19.692 ;
			RECT	145.169 19.628 145.201 19.692 ;
			RECT	145.337 19.628 145.369 19.692 ;
			RECT	145.505 19.628 145.537 19.692 ;
			RECT	145.673 19.628 145.705 19.692 ;
			RECT	145.841 19.628 145.873 19.692 ;
			RECT	146.009 19.628 146.041 19.692 ;
			RECT	146.177 19.628 146.209 19.692 ;
			RECT	146.345 19.628 146.377 19.692 ;
			RECT	146.513 19.628 146.545 19.692 ;
			RECT	146.681 19.628 146.713 19.692 ;
			RECT	146.849 19.628 146.881 19.692 ;
			RECT	147.017 19.628 147.049 19.692 ;
			RECT	147.185 19.628 147.217 19.692 ;
			RECT	147.316 19.644 147.348 19.676 ;
			RECT	147.437 19.644 147.469 19.676 ;
			RECT	147.567 19.628 147.599 19.692 ;
			RECT	149.879 19.628 149.911 19.692 ;
			RECT	151.13 19.628 151.194 19.692 ;
			RECT	151.81 19.628 151.842 19.692 ;
			RECT	152.249 19.628 152.281 19.692 ;
			RECT	153.56 19.628 153.624 19.692 ;
			RECT	156.601 19.628 156.633 19.692 ;
			RECT	156.731 19.644 156.763 19.676 ;
			RECT	156.852 19.644 156.884 19.676 ;
			RECT	156.983 19.628 157.015 19.692 ;
			RECT	157.151 19.628 157.183 19.692 ;
			RECT	157.319 19.628 157.351 19.692 ;
			RECT	157.487 19.628 157.519 19.692 ;
			RECT	157.655 19.628 157.687 19.692 ;
			RECT	157.823 19.628 157.855 19.692 ;
			RECT	157.991 19.628 158.023 19.692 ;
			RECT	158.159 19.628 158.191 19.692 ;
			RECT	158.327 19.628 158.359 19.692 ;
			RECT	158.495 19.628 158.527 19.692 ;
			RECT	158.663 19.628 158.695 19.692 ;
			RECT	158.831 19.628 158.863 19.692 ;
			RECT	158.999 19.628 159.031 19.692 ;
			RECT	159.167 19.628 159.199 19.692 ;
			RECT	159.335 19.628 159.367 19.692 ;
			RECT	159.503 19.628 159.535 19.692 ;
			RECT	159.671 19.628 159.703 19.692 ;
			RECT	159.839 19.628 159.871 19.692 ;
			RECT	160.007 19.628 160.039 19.692 ;
			RECT	160.175 19.628 160.207 19.692 ;
			RECT	160.343 19.628 160.375 19.692 ;
			RECT	160.511 19.628 160.543 19.692 ;
			RECT	160.679 19.628 160.711 19.692 ;
			RECT	160.847 19.628 160.879 19.692 ;
			RECT	161.015 19.628 161.047 19.692 ;
			RECT	161.183 19.628 161.215 19.692 ;
			RECT	161.351 19.628 161.383 19.692 ;
			RECT	161.519 19.628 161.551 19.692 ;
			RECT	161.687 19.628 161.719 19.692 ;
			RECT	161.855 19.628 161.887 19.692 ;
			RECT	162.023 19.628 162.055 19.692 ;
			RECT	162.191 19.628 162.223 19.692 ;
			RECT	162.359 19.628 162.391 19.692 ;
			RECT	162.527 19.628 162.559 19.692 ;
			RECT	162.695 19.628 162.727 19.692 ;
			RECT	162.863 19.628 162.895 19.692 ;
			RECT	163.031 19.628 163.063 19.692 ;
			RECT	163.199 19.628 163.231 19.692 ;
			RECT	163.367 19.628 163.399 19.692 ;
			RECT	163.535 19.628 163.567 19.692 ;
			RECT	163.703 19.628 163.735 19.692 ;
			RECT	163.871 19.628 163.903 19.692 ;
			RECT	164.039 19.628 164.071 19.692 ;
			RECT	164.207 19.628 164.239 19.692 ;
			RECT	164.375 19.628 164.407 19.692 ;
			RECT	164.543 19.628 164.575 19.692 ;
			RECT	164.711 19.628 164.743 19.692 ;
			RECT	164.879 19.628 164.911 19.692 ;
			RECT	165.047 19.628 165.079 19.692 ;
			RECT	165.215 19.628 165.247 19.692 ;
			RECT	165.383 19.628 165.415 19.692 ;
			RECT	165.551 19.628 165.583 19.692 ;
			RECT	165.719 19.628 165.751 19.692 ;
			RECT	165.887 19.628 165.919 19.692 ;
			RECT	166.055 19.628 166.087 19.692 ;
			RECT	166.223 19.628 166.255 19.692 ;
			RECT	166.391 19.628 166.423 19.692 ;
			RECT	166.559 19.628 166.591 19.692 ;
			RECT	166.727 19.628 166.759 19.692 ;
			RECT	166.895 19.628 166.927 19.692 ;
			RECT	167.063 19.628 167.095 19.692 ;
			RECT	167.231 19.628 167.263 19.692 ;
			RECT	167.399 19.628 167.431 19.692 ;
			RECT	167.567 19.628 167.599 19.692 ;
			RECT	167.735 19.628 167.767 19.692 ;
			RECT	167.903 19.628 167.935 19.692 ;
			RECT	168.071 19.628 168.103 19.692 ;
			RECT	168.239 19.628 168.271 19.692 ;
			RECT	168.407 19.628 168.439 19.692 ;
			RECT	168.575 19.628 168.607 19.692 ;
			RECT	168.743 19.628 168.775 19.692 ;
			RECT	168.911 19.628 168.943 19.692 ;
			RECT	169.079 19.628 169.111 19.692 ;
			RECT	169.247 19.628 169.279 19.692 ;
			RECT	169.415 19.628 169.447 19.692 ;
			RECT	169.583 19.628 169.615 19.692 ;
			RECT	169.751 19.628 169.783 19.692 ;
			RECT	169.919 19.628 169.951 19.692 ;
			RECT	170.087 19.628 170.119 19.692 ;
			RECT	170.255 19.628 170.287 19.692 ;
			RECT	170.423 19.628 170.455 19.692 ;
			RECT	170.591 19.628 170.623 19.692 ;
			RECT	170.759 19.628 170.791 19.692 ;
			RECT	170.927 19.628 170.959 19.692 ;
			RECT	171.095 19.628 171.127 19.692 ;
			RECT	171.263 19.628 171.295 19.692 ;
			RECT	171.431 19.628 171.463 19.692 ;
			RECT	171.599 19.628 171.631 19.692 ;
			RECT	171.767 19.628 171.799 19.692 ;
			RECT	171.935 19.628 171.967 19.692 ;
			RECT	172.103 19.628 172.135 19.692 ;
			RECT	172.271 19.628 172.303 19.692 ;
			RECT	172.439 19.628 172.471 19.692 ;
			RECT	172.607 19.628 172.639 19.692 ;
			RECT	172.775 19.628 172.807 19.692 ;
			RECT	172.943 19.628 172.975 19.692 ;
			RECT	173.111 19.628 173.143 19.692 ;
			RECT	173.279 19.628 173.311 19.692 ;
			RECT	173.447 19.628 173.479 19.692 ;
			RECT	173.615 19.628 173.647 19.692 ;
			RECT	173.783 19.628 173.815 19.692 ;
			RECT	173.951 19.628 173.983 19.692 ;
			RECT	174.119 19.628 174.151 19.692 ;
			RECT	174.287 19.628 174.319 19.692 ;
			RECT	174.455 19.628 174.487 19.692 ;
			RECT	174.623 19.628 174.655 19.692 ;
			RECT	174.791 19.628 174.823 19.692 ;
			RECT	174.959 19.628 174.991 19.692 ;
			RECT	175.127 19.628 175.159 19.692 ;
			RECT	175.295 19.628 175.327 19.692 ;
			RECT	175.463 19.628 175.495 19.692 ;
			RECT	175.631 19.628 175.663 19.692 ;
			RECT	175.799 19.628 175.831 19.692 ;
			RECT	175.967 19.628 175.999 19.692 ;
			RECT	176.135 19.628 176.167 19.692 ;
			RECT	176.303 19.628 176.335 19.692 ;
			RECT	176.471 19.628 176.503 19.692 ;
			RECT	176.639 19.628 176.671 19.692 ;
			RECT	176.807 19.628 176.839 19.692 ;
			RECT	176.975 19.628 177.007 19.692 ;
			RECT	177.143 19.628 177.175 19.692 ;
			RECT	177.311 19.628 177.343 19.692 ;
			RECT	177.479 19.628 177.511 19.692 ;
			RECT	177.647 19.628 177.679 19.692 ;
			RECT	177.815 19.628 177.847 19.692 ;
			RECT	177.983 19.628 178.015 19.692 ;
			RECT	178.151 19.628 178.183 19.692 ;
			RECT	178.319 19.628 178.351 19.692 ;
			RECT	178.487 19.628 178.519 19.692 ;
			RECT	178.655 19.628 178.687 19.692 ;
			RECT	178.823 19.628 178.855 19.692 ;
			RECT	178.991 19.628 179.023 19.692 ;
			RECT	179.159 19.628 179.191 19.692 ;
			RECT	179.327 19.628 179.359 19.692 ;
			RECT	179.495 19.628 179.527 19.692 ;
			RECT	179.663 19.628 179.695 19.692 ;
			RECT	179.831 19.628 179.863 19.692 ;
			RECT	179.999 19.628 180.031 19.692 ;
			RECT	180.167 19.628 180.199 19.692 ;
			RECT	180.335 19.628 180.367 19.692 ;
			RECT	180.503 19.628 180.535 19.692 ;
			RECT	180.671 19.628 180.703 19.692 ;
			RECT	180.839 19.628 180.871 19.692 ;
			RECT	181.007 19.628 181.039 19.692 ;
			RECT	181.175 19.628 181.207 19.692 ;
			RECT	181.343 19.628 181.375 19.692 ;
			RECT	181.511 19.628 181.543 19.692 ;
			RECT	181.679 19.628 181.711 19.692 ;
			RECT	181.847 19.628 181.879 19.692 ;
			RECT	182.015 19.628 182.047 19.692 ;
			RECT	182.183 19.628 182.215 19.692 ;
			RECT	182.351 19.628 182.383 19.692 ;
			RECT	182.519 19.628 182.551 19.692 ;
			RECT	182.687 19.628 182.719 19.692 ;
			RECT	182.855 19.628 182.887 19.692 ;
			RECT	183.023 19.628 183.055 19.692 ;
			RECT	183.191 19.628 183.223 19.692 ;
			RECT	183.359 19.628 183.391 19.692 ;
			RECT	183.527 19.628 183.559 19.692 ;
			RECT	183.695 19.628 183.727 19.692 ;
			RECT	183.863 19.628 183.895 19.692 ;
			RECT	184.031 19.628 184.063 19.692 ;
			RECT	184.199 19.628 184.231 19.692 ;
			RECT	184.367 19.628 184.399 19.692 ;
			RECT	184.535 19.628 184.567 19.692 ;
			RECT	184.703 19.628 184.735 19.692 ;
			RECT	184.871 19.628 184.903 19.692 ;
			RECT	185.039 19.628 185.071 19.692 ;
			RECT	185.207 19.628 185.239 19.692 ;
			RECT	185.375 19.628 185.407 19.692 ;
			RECT	185.543 19.628 185.575 19.692 ;
			RECT	185.711 19.628 185.743 19.692 ;
			RECT	185.879 19.628 185.911 19.692 ;
			RECT	186.047 19.628 186.079 19.692 ;
			RECT	186.215 19.628 186.247 19.692 ;
			RECT	186.383 19.628 186.415 19.692 ;
			RECT	186.551 19.628 186.583 19.692 ;
			RECT	186.719 19.628 186.751 19.692 ;
			RECT	186.887 19.628 186.919 19.692 ;
			RECT	187.055 19.628 187.087 19.692 ;
			RECT	187.223 19.628 187.255 19.692 ;
			RECT	187.391 19.628 187.423 19.692 ;
			RECT	187.559 19.628 187.591 19.692 ;
			RECT	187.727 19.628 187.759 19.692 ;
			RECT	187.895 19.628 187.927 19.692 ;
			RECT	188.063 19.628 188.095 19.692 ;
			RECT	188.231 19.628 188.263 19.692 ;
			RECT	188.399 19.628 188.431 19.692 ;
			RECT	188.567 19.628 188.599 19.692 ;
			RECT	188.735 19.628 188.767 19.692 ;
			RECT	188.903 19.628 188.935 19.692 ;
			RECT	189.071 19.628 189.103 19.692 ;
			RECT	189.239 19.628 189.271 19.692 ;
			RECT	189.407 19.628 189.439 19.692 ;
			RECT	189.575 19.628 189.607 19.692 ;
			RECT	189.743 19.628 189.775 19.692 ;
			RECT	189.911 19.628 189.943 19.692 ;
			RECT	190.079 19.628 190.111 19.692 ;
			RECT	190.247 19.628 190.279 19.692 ;
			RECT	190.415 19.628 190.447 19.692 ;
			RECT	190.583 19.628 190.615 19.692 ;
			RECT	190.751 19.628 190.783 19.692 ;
			RECT	190.919 19.628 190.951 19.692 ;
			RECT	191.087 19.628 191.119 19.692 ;
			RECT	191.255 19.628 191.287 19.692 ;
			RECT	191.423 19.628 191.455 19.692 ;
			RECT	191.591 19.628 191.623 19.692 ;
			RECT	191.759 19.628 191.791 19.692 ;
			RECT	191.927 19.628 191.959 19.692 ;
			RECT	192.095 19.628 192.127 19.692 ;
			RECT	192.263 19.628 192.295 19.692 ;
			RECT	192.431 19.628 192.463 19.692 ;
			RECT	192.599 19.628 192.631 19.692 ;
			RECT	192.767 19.628 192.799 19.692 ;
			RECT	192.935 19.628 192.967 19.692 ;
			RECT	193.103 19.628 193.135 19.692 ;
			RECT	193.271 19.628 193.303 19.692 ;
			RECT	193.439 19.628 193.471 19.692 ;
			RECT	193.607 19.628 193.639 19.692 ;
			RECT	193.775 19.628 193.807 19.692 ;
			RECT	193.943 19.628 193.975 19.692 ;
			RECT	194.111 19.628 194.143 19.692 ;
			RECT	194.279 19.628 194.311 19.692 ;
			RECT	194.447 19.628 194.479 19.692 ;
			RECT	194.615 19.628 194.647 19.692 ;
			RECT	194.783 19.628 194.815 19.692 ;
			RECT	194.951 19.628 194.983 19.692 ;
			RECT	195.119 19.628 195.151 19.692 ;
			RECT	195.287 19.628 195.319 19.692 ;
			RECT	195.455 19.628 195.487 19.692 ;
			RECT	195.623 19.628 195.655 19.692 ;
			RECT	195.791 19.628 195.823 19.692 ;
			RECT	195.959 19.628 195.991 19.692 ;
			RECT	196.127 19.628 196.159 19.692 ;
			RECT	196.295 19.628 196.327 19.692 ;
			RECT	196.463 19.628 196.495 19.692 ;
			RECT	196.631 19.628 196.663 19.692 ;
			RECT	196.799 19.628 196.831 19.692 ;
			RECT	196.967 19.628 196.999 19.692 ;
			RECT	197.135 19.628 197.167 19.692 ;
			RECT	197.303 19.628 197.335 19.692 ;
			RECT	197.471 19.628 197.503 19.692 ;
			RECT	197.639 19.628 197.671 19.692 ;
			RECT	197.807 19.628 197.839 19.692 ;
			RECT	197.975 19.628 198.007 19.692 ;
			RECT	198.143 19.628 198.175 19.692 ;
			RECT	198.311 19.628 198.343 19.692 ;
			RECT	198.479 19.628 198.511 19.692 ;
			RECT	198.647 19.628 198.679 19.692 ;
			RECT	198.815 19.628 198.847 19.692 ;
			RECT	198.983 19.628 199.015 19.692 ;
			RECT	199.151 19.628 199.183 19.692 ;
			RECT	199.319 19.628 199.351 19.692 ;
			RECT	199.487 19.628 199.519 19.692 ;
			RECT	199.655 19.628 199.687 19.692 ;
			RECT	199.823 19.628 199.855 19.692 ;
			RECT	199.991 19.628 200.023 19.692 ;
			RECT	200.121 19.644 200.153 19.676 ;
			RECT	200.243 19.649 200.275 19.681 ;
			RECT	200.373 19.628 200.405 19.692 ;
			RECT	200.9 19.628 200.932 19.692 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 17.68 201.665 17.8 ;
			LAYER	J3 ;
			RECT	0.755 17.708 0.787 17.772 ;
			RECT	1.645 17.708 1.709 17.772 ;
			RECT	2.323 17.708 2.387 17.772 ;
			RECT	3.438 17.708 3.47 17.772 ;
			RECT	3.585 17.708 3.617 17.772 ;
			RECT	4.195 17.708 4.227 17.772 ;
			RECT	4.72 17.708 4.752 17.772 ;
			RECT	4.944 17.708 5.008 17.772 ;
			RECT	5.267 17.708 5.299 17.772 ;
			RECT	5.797 17.708 5.829 17.772 ;
			RECT	5.927 17.729 5.959 17.761 ;
			RECT	6.049 17.724 6.081 17.756 ;
			RECT	6.179 17.708 6.211 17.772 ;
			RECT	6.347 17.708 6.379 17.772 ;
			RECT	6.515 17.708 6.547 17.772 ;
			RECT	6.683 17.708 6.715 17.772 ;
			RECT	6.851 17.708 6.883 17.772 ;
			RECT	7.019 17.708 7.051 17.772 ;
			RECT	7.187 17.708 7.219 17.772 ;
			RECT	7.355 17.708 7.387 17.772 ;
			RECT	7.523 17.708 7.555 17.772 ;
			RECT	7.691 17.708 7.723 17.772 ;
			RECT	7.859 17.708 7.891 17.772 ;
			RECT	8.027 17.708 8.059 17.772 ;
			RECT	8.195 17.708 8.227 17.772 ;
			RECT	8.363 17.708 8.395 17.772 ;
			RECT	8.531 17.708 8.563 17.772 ;
			RECT	8.699 17.708 8.731 17.772 ;
			RECT	8.867 17.708 8.899 17.772 ;
			RECT	9.035 17.708 9.067 17.772 ;
			RECT	9.203 17.708 9.235 17.772 ;
			RECT	9.371 17.708 9.403 17.772 ;
			RECT	9.539 17.708 9.571 17.772 ;
			RECT	9.707 17.708 9.739 17.772 ;
			RECT	9.875 17.708 9.907 17.772 ;
			RECT	10.043 17.708 10.075 17.772 ;
			RECT	10.211 17.708 10.243 17.772 ;
			RECT	10.379 17.708 10.411 17.772 ;
			RECT	10.547 17.708 10.579 17.772 ;
			RECT	10.715 17.708 10.747 17.772 ;
			RECT	10.883 17.708 10.915 17.772 ;
			RECT	11.051 17.708 11.083 17.772 ;
			RECT	11.219 17.708 11.251 17.772 ;
			RECT	11.387 17.708 11.419 17.772 ;
			RECT	11.555 17.708 11.587 17.772 ;
			RECT	11.723 17.708 11.755 17.772 ;
			RECT	11.891 17.708 11.923 17.772 ;
			RECT	12.059 17.708 12.091 17.772 ;
			RECT	12.227 17.708 12.259 17.772 ;
			RECT	12.395 17.708 12.427 17.772 ;
			RECT	12.563 17.708 12.595 17.772 ;
			RECT	12.731 17.708 12.763 17.772 ;
			RECT	12.899 17.708 12.931 17.772 ;
			RECT	13.067 17.708 13.099 17.772 ;
			RECT	13.235 17.708 13.267 17.772 ;
			RECT	13.403 17.708 13.435 17.772 ;
			RECT	13.571 17.708 13.603 17.772 ;
			RECT	13.739 17.708 13.771 17.772 ;
			RECT	13.907 17.708 13.939 17.772 ;
			RECT	14.075 17.708 14.107 17.772 ;
			RECT	14.243 17.708 14.275 17.772 ;
			RECT	14.411 17.708 14.443 17.772 ;
			RECT	14.579 17.708 14.611 17.772 ;
			RECT	14.747 17.708 14.779 17.772 ;
			RECT	14.915 17.708 14.947 17.772 ;
			RECT	15.083 17.708 15.115 17.772 ;
			RECT	15.251 17.708 15.283 17.772 ;
			RECT	15.419 17.708 15.451 17.772 ;
			RECT	15.587 17.708 15.619 17.772 ;
			RECT	15.755 17.708 15.787 17.772 ;
			RECT	15.923 17.708 15.955 17.772 ;
			RECT	16.091 17.708 16.123 17.772 ;
			RECT	16.259 17.708 16.291 17.772 ;
			RECT	16.427 17.708 16.459 17.772 ;
			RECT	16.595 17.708 16.627 17.772 ;
			RECT	16.763 17.708 16.795 17.772 ;
			RECT	16.931 17.708 16.963 17.772 ;
			RECT	17.099 17.708 17.131 17.772 ;
			RECT	17.267 17.708 17.299 17.772 ;
			RECT	17.435 17.708 17.467 17.772 ;
			RECT	17.603 17.708 17.635 17.772 ;
			RECT	17.771 17.708 17.803 17.772 ;
			RECT	17.939 17.708 17.971 17.772 ;
			RECT	18.107 17.708 18.139 17.772 ;
			RECT	18.275 17.708 18.307 17.772 ;
			RECT	18.443 17.708 18.475 17.772 ;
			RECT	18.611 17.708 18.643 17.772 ;
			RECT	18.779 17.708 18.811 17.772 ;
			RECT	18.947 17.708 18.979 17.772 ;
			RECT	19.115 17.708 19.147 17.772 ;
			RECT	19.283 17.708 19.315 17.772 ;
			RECT	19.451 17.708 19.483 17.772 ;
			RECT	19.619 17.708 19.651 17.772 ;
			RECT	19.787 17.708 19.819 17.772 ;
			RECT	19.955 17.708 19.987 17.772 ;
			RECT	20.123 17.708 20.155 17.772 ;
			RECT	20.291 17.708 20.323 17.772 ;
			RECT	20.459 17.708 20.491 17.772 ;
			RECT	20.627 17.708 20.659 17.772 ;
			RECT	20.795 17.708 20.827 17.772 ;
			RECT	20.963 17.708 20.995 17.772 ;
			RECT	21.131 17.708 21.163 17.772 ;
			RECT	21.299 17.708 21.331 17.772 ;
			RECT	21.467 17.708 21.499 17.772 ;
			RECT	21.635 17.708 21.667 17.772 ;
			RECT	21.803 17.708 21.835 17.772 ;
			RECT	21.971 17.708 22.003 17.772 ;
			RECT	22.139 17.708 22.171 17.772 ;
			RECT	22.307 17.708 22.339 17.772 ;
			RECT	22.475 17.708 22.507 17.772 ;
			RECT	22.643 17.708 22.675 17.772 ;
			RECT	22.811 17.708 22.843 17.772 ;
			RECT	22.979 17.708 23.011 17.772 ;
			RECT	23.147 17.708 23.179 17.772 ;
			RECT	23.315 17.708 23.347 17.772 ;
			RECT	23.483 17.708 23.515 17.772 ;
			RECT	23.651 17.708 23.683 17.772 ;
			RECT	23.819 17.708 23.851 17.772 ;
			RECT	23.987 17.708 24.019 17.772 ;
			RECT	24.155 17.708 24.187 17.772 ;
			RECT	24.323 17.708 24.355 17.772 ;
			RECT	24.491 17.708 24.523 17.772 ;
			RECT	24.659 17.708 24.691 17.772 ;
			RECT	24.827 17.708 24.859 17.772 ;
			RECT	24.995 17.708 25.027 17.772 ;
			RECT	25.163 17.708 25.195 17.772 ;
			RECT	25.331 17.708 25.363 17.772 ;
			RECT	25.499 17.708 25.531 17.772 ;
			RECT	25.667 17.708 25.699 17.772 ;
			RECT	25.835 17.708 25.867 17.772 ;
			RECT	26.003 17.708 26.035 17.772 ;
			RECT	26.171 17.708 26.203 17.772 ;
			RECT	26.339 17.708 26.371 17.772 ;
			RECT	26.507 17.708 26.539 17.772 ;
			RECT	26.675 17.708 26.707 17.772 ;
			RECT	26.843 17.708 26.875 17.772 ;
			RECT	27.011 17.708 27.043 17.772 ;
			RECT	27.179 17.708 27.211 17.772 ;
			RECT	27.347 17.708 27.379 17.772 ;
			RECT	27.515 17.708 27.547 17.772 ;
			RECT	27.683 17.708 27.715 17.772 ;
			RECT	27.851 17.708 27.883 17.772 ;
			RECT	28.019 17.708 28.051 17.772 ;
			RECT	28.187 17.708 28.219 17.772 ;
			RECT	28.355 17.708 28.387 17.772 ;
			RECT	28.523 17.708 28.555 17.772 ;
			RECT	28.691 17.708 28.723 17.772 ;
			RECT	28.859 17.708 28.891 17.772 ;
			RECT	29.027 17.708 29.059 17.772 ;
			RECT	29.195 17.708 29.227 17.772 ;
			RECT	29.363 17.708 29.395 17.772 ;
			RECT	29.531 17.708 29.563 17.772 ;
			RECT	29.699 17.708 29.731 17.772 ;
			RECT	29.867 17.708 29.899 17.772 ;
			RECT	30.035 17.708 30.067 17.772 ;
			RECT	30.203 17.708 30.235 17.772 ;
			RECT	30.371 17.708 30.403 17.772 ;
			RECT	30.539 17.708 30.571 17.772 ;
			RECT	30.707 17.708 30.739 17.772 ;
			RECT	30.875 17.708 30.907 17.772 ;
			RECT	31.043 17.708 31.075 17.772 ;
			RECT	31.211 17.708 31.243 17.772 ;
			RECT	31.379 17.708 31.411 17.772 ;
			RECT	31.547 17.708 31.579 17.772 ;
			RECT	31.715 17.708 31.747 17.772 ;
			RECT	31.883 17.708 31.915 17.772 ;
			RECT	32.051 17.708 32.083 17.772 ;
			RECT	32.219 17.708 32.251 17.772 ;
			RECT	32.387 17.708 32.419 17.772 ;
			RECT	32.555 17.708 32.587 17.772 ;
			RECT	32.723 17.708 32.755 17.772 ;
			RECT	32.891 17.708 32.923 17.772 ;
			RECT	33.059 17.708 33.091 17.772 ;
			RECT	33.227 17.708 33.259 17.772 ;
			RECT	33.395 17.708 33.427 17.772 ;
			RECT	33.563 17.708 33.595 17.772 ;
			RECT	33.731 17.708 33.763 17.772 ;
			RECT	33.899 17.708 33.931 17.772 ;
			RECT	34.067 17.708 34.099 17.772 ;
			RECT	34.235 17.708 34.267 17.772 ;
			RECT	34.403 17.708 34.435 17.772 ;
			RECT	34.571 17.708 34.603 17.772 ;
			RECT	34.739 17.708 34.771 17.772 ;
			RECT	34.907 17.708 34.939 17.772 ;
			RECT	35.075 17.708 35.107 17.772 ;
			RECT	35.243 17.708 35.275 17.772 ;
			RECT	35.411 17.708 35.443 17.772 ;
			RECT	35.579 17.708 35.611 17.772 ;
			RECT	35.747 17.708 35.779 17.772 ;
			RECT	35.915 17.708 35.947 17.772 ;
			RECT	36.083 17.708 36.115 17.772 ;
			RECT	36.251 17.708 36.283 17.772 ;
			RECT	36.419 17.708 36.451 17.772 ;
			RECT	36.587 17.708 36.619 17.772 ;
			RECT	36.755 17.708 36.787 17.772 ;
			RECT	36.923 17.708 36.955 17.772 ;
			RECT	37.091 17.708 37.123 17.772 ;
			RECT	37.259 17.708 37.291 17.772 ;
			RECT	37.427 17.708 37.459 17.772 ;
			RECT	37.595 17.708 37.627 17.772 ;
			RECT	37.763 17.708 37.795 17.772 ;
			RECT	37.931 17.708 37.963 17.772 ;
			RECT	38.099 17.708 38.131 17.772 ;
			RECT	38.267 17.708 38.299 17.772 ;
			RECT	38.435 17.708 38.467 17.772 ;
			RECT	38.603 17.708 38.635 17.772 ;
			RECT	38.771 17.708 38.803 17.772 ;
			RECT	38.939 17.708 38.971 17.772 ;
			RECT	39.107 17.708 39.139 17.772 ;
			RECT	39.275 17.708 39.307 17.772 ;
			RECT	39.443 17.708 39.475 17.772 ;
			RECT	39.611 17.708 39.643 17.772 ;
			RECT	39.779 17.708 39.811 17.772 ;
			RECT	39.947 17.708 39.979 17.772 ;
			RECT	40.115 17.708 40.147 17.772 ;
			RECT	40.283 17.708 40.315 17.772 ;
			RECT	40.451 17.708 40.483 17.772 ;
			RECT	40.619 17.708 40.651 17.772 ;
			RECT	40.787 17.708 40.819 17.772 ;
			RECT	40.955 17.708 40.987 17.772 ;
			RECT	41.123 17.708 41.155 17.772 ;
			RECT	41.291 17.708 41.323 17.772 ;
			RECT	41.459 17.708 41.491 17.772 ;
			RECT	41.627 17.708 41.659 17.772 ;
			RECT	41.795 17.708 41.827 17.772 ;
			RECT	41.963 17.708 41.995 17.772 ;
			RECT	42.131 17.708 42.163 17.772 ;
			RECT	42.299 17.708 42.331 17.772 ;
			RECT	42.467 17.708 42.499 17.772 ;
			RECT	42.635 17.708 42.667 17.772 ;
			RECT	42.803 17.708 42.835 17.772 ;
			RECT	42.971 17.708 43.003 17.772 ;
			RECT	43.139 17.708 43.171 17.772 ;
			RECT	43.307 17.708 43.339 17.772 ;
			RECT	43.475 17.708 43.507 17.772 ;
			RECT	43.643 17.708 43.675 17.772 ;
			RECT	43.811 17.708 43.843 17.772 ;
			RECT	43.979 17.708 44.011 17.772 ;
			RECT	44.147 17.708 44.179 17.772 ;
			RECT	44.315 17.708 44.347 17.772 ;
			RECT	44.483 17.708 44.515 17.772 ;
			RECT	44.651 17.708 44.683 17.772 ;
			RECT	44.819 17.708 44.851 17.772 ;
			RECT	44.987 17.708 45.019 17.772 ;
			RECT	45.155 17.708 45.187 17.772 ;
			RECT	45.323 17.708 45.355 17.772 ;
			RECT	45.491 17.708 45.523 17.772 ;
			RECT	45.659 17.708 45.691 17.772 ;
			RECT	45.827 17.708 45.859 17.772 ;
			RECT	45.995 17.708 46.027 17.772 ;
			RECT	46.163 17.708 46.195 17.772 ;
			RECT	46.331 17.708 46.363 17.772 ;
			RECT	46.499 17.708 46.531 17.772 ;
			RECT	46.667 17.708 46.699 17.772 ;
			RECT	46.835 17.708 46.867 17.772 ;
			RECT	47.003 17.708 47.035 17.772 ;
			RECT	47.171 17.708 47.203 17.772 ;
			RECT	47.339 17.708 47.371 17.772 ;
			RECT	47.507 17.708 47.539 17.772 ;
			RECT	47.675 17.708 47.707 17.772 ;
			RECT	47.843 17.708 47.875 17.772 ;
			RECT	48.011 17.708 48.043 17.772 ;
			RECT	48.179 17.708 48.211 17.772 ;
			RECT	48.347 17.708 48.379 17.772 ;
			RECT	48.515 17.708 48.547 17.772 ;
			RECT	48.683 17.708 48.715 17.772 ;
			RECT	48.851 17.708 48.883 17.772 ;
			RECT	49.019 17.708 49.051 17.772 ;
			RECT	49.187 17.708 49.219 17.772 ;
			RECT	49.318 17.724 49.35 17.756 ;
			RECT	49.439 17.724 49.471 17.756 ;
			RECT	49.569 17.708 49.601 17.772 ;
			RECT	51.881 17.708 51.913 17.772 ;
			RECT	53.132 17.708 53.196 17.772 ;
			RECT	53.812 17.708 53.844 17.772 ;
			RECT	54.251 17.708 54.283 17.772 ;
			RECT	55.562 17.708 55.626 17.772 ;
			RECT	58.603 17.708 58.635 17.772 ;
			RECT	58.733 17.724 58.765 17.756 ;
			RECT	58.854 17.724 58.886 17.756 ;
			RECT	58.985 17.708 59.017 17.772 ;
			RECT	59.153 17.708 59.185 17.772 ;
			RECT	59.321 17.708 59.353 17.772 ;
			RECT	59.489 17.708 59.521 17.772 ;
			RECT	59.657 17.708 59.689 17.772 ;
			RECT	59.825 17.708 59.857 17.772 ;
			RECT	59.993 17.708 60.025 17.772 ;
			RECT	60.161 17.708 60.193 17.772 ;
			RECT	60.329 17.708 60.361 17.772 ;
			RECT	60.497 17.708 60.529 17.772 ;
			RECT	60.665 17.708 60.697 17.772 ;
			RECT	60.833 17.708 60.865 17.772 ;
			RECT	61.001 17.708 61.033 17.772 ;
			RECT	61.169 17.708 61.201 17.772 ;
			RECT	61.337 17.708 61.369 17.772 ;
			RECT	61.505 17.708 61.537 17.772 ;
			RECT	61.673 17.708 61.705 17.772 ;
			RECT	61.841 17.708 61.873 17.772 ;
			RECT	62.009 17.708 62.041 17.772 ;
			RECT	62.177 17.708 62.209 17.772 ;
			RECT	62.345 17.708 62.377 17.772 ;
			RECT	62.513 17.708 62.545 17.772 ;
			RECT	62.681 17.708 62.713 17.772 ;
			RECT	62.849 17.708 62.881 17.772 ;
			RECT	63.017 17.708 63.049 17.772 ;
			RECT	63.185 17.708 63.217 17.772 ;
			RECT	63.353 17.708 63.385 17.772 ;
			RECT	63.521 17.708 63.553 17.772 ;
			RECT	63.689 17.708 63.721 17.772 ;
			RECT	63.857 17.708 63.889 17.772 ;
			RECT	64.025 17.708 64.057 17.772 ;
			RECT	64.193 17.708 64.225 17.772 ;
			RECT	64.361 17.708 64.393 17.772 ;
			RECT	64.529 17.708 64.561 17.772 ;
			RECT	64.697 17.708 64.729 17.772 ;
			RECT	64.865 17.708 64.897 17.772 ;
			RECT	65.033 17.708 65.065 17.772 ;
			RECT	65.201 17.708 65.233 17.772 ;
			RECT	65.369 17.708 65.401 17.772 ;
			RECT	65.537 17.708 65.569 17.772 ;
			RECT	65.705 17.708 65.737 17.772 ;
			RECT	65.873 17.708 65.905 17.772 ;
			RECT	66.041 17.708 66.073 17.772 ;
			RECT	66.209 17.708 66.241 17.772 ;
			RECT	66.377 17.708 66.409 17.772 ;
			RECT	66.545 17.708 66.577 17.772 ;
			RECT	66.713 17.708 66.745 17.772 ;
			RECT	66.881 17.708 66.913 17.772 ;
			RECT	67.049 17.708 67.081 17.772 ;
			RECT	67.217 17.708 67.249 17.772 ;
			RECT	67.385 17.708 67.417 17.772 ;
			RECT	67.553 17.708 67.585 17.772 ;
			RECT	67.721 17.708 67.753 17.772 ;
			RECT	67.889 17.708 67.921 17.772 ;
			RECT	68.057 17.708 68.089 17.772 ;
			RECT	68.225 17.708 68.257 17.772 ;
			RECT	68.393 17.708 68.425 17.772 ;
			RECT	68.561 17.708 68.593 17.772 ;
			RECT	68.729 17.708 68.761 17.772 ;
			RECT	68.897 17.708 68.929 17.772 ;
			RECT	69.065 17.708 69.097 17.772 ;
			RECT	69.233 17.708 69.265 17.772 ;
			RECT	69.401 17.708 69.433 17.772 ;
			RECT	69.569 17.708 69.601 17.772 ;
			RECT	69.737 17.708 69.769 17.772 ;
			RECT	69.905 17.708 69.937 17.772 ;
			RECT	70.073 17.708 70.105 17.772 ;
			RECT	70.241 17.708 70.273 17.772 ;
			RECT	70.409 17.708 70.441 17.772 ;
			RECT	70.577 17.708 70.609 17.772 ;
			RECT	70.745 17.708 70.777 17.772 ;
			RECT	70.913 17.708 70.945 17.772 ;
			RECT	71.081 17.708 71.113 17.772 ;
			RECT	71.249 17.708 71.281 17.772 ;
			RECT	71.417 17.708 71.449 17.772 ;
			RECT	71.585 17.708 71.617 17.772 ;
			RECT	71.753 17.708 71.785 17.772 ;
			RECT	71.921 17.708 71.953 17.772 ;
			RECT	72.089 17.708 72.121 17.772 ;
			RECT	72.257 17.708 72.289 17.772 ;
			RECT	72.425 17.708 72.457 17.772 ;
			RECT	72.593 17.708 72.625 17.772 ;
			RECT	72.761 17.708 72.793 17.772 ;
			RECT	72.929 17.708 72.961 17.772 ;
			RECT	73.097 17.708 73.129 17.772 ;
			RECT	73.265 17.708 73.297 17.772 ;
			RECT	73.433 17.708 73.465 17.772 ;
			RECT	73.601 17.708 73.633 17.772 ;
			RECT	73.769 17.708 73.801 17.772 ;
			RECT	73.937 17.708 73.969 17.772 ;
			RECT	74.105 17.708 74.137 17.772 ;
			RECT	74.273 17.708 74.305 17.772 ;
			RECT	74.441 17.708 74.473 17.772 ;
			RECT	74.609 17.708 74.641 17.772 ;
			RECT	74.777 17.708 74.809 17.772 ;
			RECT	74.945 17.708 74.977 17.772 ;
			RECT	75.113 17.708 75.145 17.772 ;
			RECT	75.281 17.708 75.313 17.772 ;
			RECT	75.449 17.708 75.481 17.772 ;
			RECT	75.617 17.708 75.649 17.772 ;
			RECT	75.785 17.708 75.817 17.772 ;
			RECT	75.953 17.708 75.985 17.772 ;
			RECT	76.121 17.708 76.153 17.772 ;
			RECT	76.289 17.708 76.321 17.772 ;
			RECT	76.457 17.708 76.489 17.772 ;
			RECT	76.625 17.708 76.657 17.772 ;
			RECT	76.793 17.708 76.825 17.772 ;
			RECT	76.961 17.708 76.993 17.772 ;
			RECT	77.129 17.708 77.161 17.772 ;
			RECT	77.297 17.708 77.329 17.772 ;
			RECT	77.465 17.708 77.497 17.772 ;
			RECT	77.633 17.708 77.665 17.772 ;
			RECT	77.801 17.708 77.833 17.772 ;
			RECT	77.969 17.708 78.001 17.772 ;
			RECT	78.137 17.708 78.169 17.772 ;
			RECT	78.305 17.708 78.337 17.772 ;
			RECT	78.473 17.708 78.505 17.772 ;
			RECT	78.641 17.708 78.673 17.772 ;
			RECT	78.809 17.708 78.841 17.772 ;
			RECT	78.977 17.708 79.009 17.772 ;
			RECT	79.145 17.708 79.177 17.772 ;
			RECT	79.313 17.708 79.345 17.772 ;
			RECT	79.481 17.708 79.513 17.772 ;
			RECT	79.649 17.708 79.681 17.772 ;
			RECT	79.817 17.708 79.849 17.772 ;
			RECT	79.985 17.708 80.017 17.772 ;
			RECT	80.153 17.708 80.185 17.772 ;
			RECT	80.321 17.708 80.353 17.772 ;
			RECT	80.489 17.708 80.521 17.772 ;
			RECT	80.657 17.708 80.689 17.772 ;
			RECT	80.825 17.708 80.857 17.772 ;
			RECT	80.993 17.708 81.025 17.772 ;
			RECT	81.161 17.708 81.193 17.772 ;
			RECT	81.329 17.708 81.361 17.772 ;
			RECT	81.497 17.708 81.529 17.772 ;
			RECT	81.665 17.708 81.697 17.772 ;
			RECT	81.833 17.708 81.865 17.772 ;
			RECT	82.001 17.708 82.033 17.772 ;
			RECT	82.169 17.708 82.201 17.772 ;
			RECT	82.337 17.708 82.369 17.772 ;
			RECT	82.505 17.708 82.537 17.772 ;
			RECT	82.673 17.708 82.705 17.772 ;
			RECT	82.841 17.708 82.873 17.772 ;
			RECT	83.009 17.708 83.041 17.772 ;
			RECT	83.177 17.708 83.209 17.772 ;
			RECT	83.345 17.708 83.377 17.772 ;
			RECT	83.513 17.708 83.545 17.772 ;
			RECT	83.681 17.708 83.713 17.772 ;
			RECT	83.849 17.708 83.881 17.772 ;
			RECT	84.017 17.708 84.049 17.772 ;
			RECT	84.185 17.708 84.217 17.772 ;
			RECT	84.353 17.708 84.385 17.772 ;
			RECT	84.521 17.708 84.553 17.772 ;
			RECT	84.689 17.708 84.721 17.772 ;
			RECT	84.857 17.708 84.889 17.772 ;
			RECT	85.025 17.708 85.057 17.772 ;
			RECT	85.193 17.708 85.225 17.772 ;
			RECT	85.361 17.708 85.393 17.772 ;
			RECT	85.529 17.708 85.561 17.772 ;
			RECT	85.697 17.708 85.729 17.772 ;
			RECT	85.865 17.708 85.897 17.772 ;
			RECT	86.033 17.708 86.065 17.772 ;
			RECT	86.201 17.708 86.233 17.772 ;
			RECT	86.369 17.708 86.401 17.772 ;
			RECT	86.537 17.708 86.569 17.772 ;
			RECT	86.705 17.708 86.737 17.772 ;
			RECT	86.873 17.708 86.905 17.772 ;
			RECT	87.041 17.708 87.073 17.772 ;
			RECT	87.209 17.708 87.241 17.772 ;
			RECT	87.377 17.708 87.409 17.772 ;
			RECT	87.545 17.708 87.577 17.772 ;
			RECT	87.713 17.708 87.745 17.772 ;
			RECT	87.881 17.708 87.913 17.772 ;
			RECT	88.049 17.708 88.081 17.772 ;
			RECT	88.217 17.708 88.249 17.772 ;
			RECT	88.385 17.708 88.417 17.772 ;
			RECT	88.553 17.708 88.585 17.772 ;
			RECT	88.721 17.708 88.753 17.772 ;
			RECT	88.889 17.708 88.921 17.772 ;
			RECT	89.057 17.708 89.089 17.772 ;
			RECT	89.225 17.708 89.257 17.772 ;
			RECT	89.393 17.708 89.425 17.772 ;
			RECT	89.561 17.708 89.593 17.772 ;
			RECT	89.729 17.708 89.761 17.772 ;
			RECT	89.897 17.708 89.929 17.772 ;
			RECT	90.065 17.708 90.097 17.772 ;
			RECT	90.233 17.708 90.265 17.772 ;
			RECT	90.401 17.708 90.433 17.772 ;
			RECT	90.569 17.708 90.601 17.772 ;
			RECT	90.737 17.708 90.769 17.772 ;
			RECT	90.905 17.708 90.937 17.772 ;
			RECT	91.073 17.708 91.105 17.772 ;
			RECT	91.241 17.708 91.273 17.772 ;
			RECT	91.409 17.708 91.441 17.772 ;
			RECT	91.577 17.708 91.609 17.772 ;
			RECT	91.745 17.708 91.777 17.772 ;
			RECT	91.913 17.708 91.945 17.772 ;
			RECT	92.081 17.708 92.113 17.772 ;
			RECT	92.249 17.708 92.281 17.772 ;
			RECT	92.417 17.708 92.449 17.772 ;
			RECT	92.585 17.708 92.617 17.772 ;
			RECT	92.753 17.708 92.785 17.772 ;
			RECT	92.921 17.708 92.953 17.772 ;
			RECT	93.089 17.708 93.121 17.772 ;
			RECT	93.257 17.708 93.289 17.772 ;
			RECT	93.425 17.708 93.457 17.772 ;
			RECT	93.593 17.708 93.625 17.772 ;
			RECT	93.761 17.708 93.793 17.772 ;
			RECT	93.929 17.708 93.961 17.772 ;
			RECT	94.097 17.708 94.129 17.772 ;
			RECT	94.265 17.708 94.297 17.772 ;
			RECT	94.433 17.708 94.465 17.772 ;
			RECT	94.601 17.708 94.633 17.772 ;
			RECT	94.769 17.708 94.801 17.772 ;
			RECT	94.937 17.708 94.969 17.772 ;
			RECT	95.105 17.708 95.137 17.772 ;
			RECT	95.273 17.708 95.305 17.772 ;
			RECT	95.441 17.708 95.473 17.772 ;
			RECT	95.609 17.708 95.641 17.772 ;
			RECT	95.777 17.708 95.809 17.772 ;
			RECT	95.945 17.708 95.977 17.772 ;
			RECT	96.113 17.708 96.145 17.772 ;
			RECT	96.281 17.708 96.313 17.772 ;
			RECT	96.449 17.708 96.481 17.772 ;
			RECT	96.617 17.708 96.649 17.772 ;
			RECT	96.785 17.708 96.817 17.772 ;
			RECT	96.953 17.708 96.985 17.772 ;
			RECT	97.121 17.708 97.153 17.772 ;
			RECT	97.289 17.708 97.321 17.772 ;
			RECT	97.457 17.708 97.489 17.772 ;
			RECT	97.625 17.708 97.657 17.772 ;
			RECT	97.793 17.708 97.825 17.772 ;
			RECT	97.961 17.708 97.993 17.772 ;
			RECT	98.129 17.708 98.161 17.772 ;
			RECT	98.297 17.708 98.329 17.772 ;
			RECT	98.465 17.708 98.497 17.772 ;
			RECT	98.633 17.708 98.665 17.772 ;
			RECT	98.801 17.708 98.833 17.772 ;
			RECT	98.969 17.708 99.001 17.772 ;
			RECT	99.137 17.708 99.169 17.772 ;
			RECT	99.305 17.708 99.337 17.772 ;
			RECT	99.473 17.708 99.505 17.772 ;
			RECT	99.641 17.708 99.673 17.772 ;
			RECT	99.809 17.708 99.841 17.772 ;
			RECT	99.977 17.708 100.009 17.772 ;
			RECT	100.145 17.708 100.177 17.772 ;
			RECT	100.313 17.708 100.345 17.772 ;
			RECT	100.481 17.708 100.513 17.772 ;
			RECT	100.649 17.708 100.681 17.772 ;
			RECT	100.817 17.708 100.849 17.772 ;
			RECT	100.985 17.708 101.017 17.772 ;
			RECT	101.153 17.708 101.185 17.772 ;
			RECT	101.321 17.708 101.353 17.772 ;
			RECT	101.489 17.708 101.521 17.772 ;
			RECT	101.657 17.708 101.689 17.772 ;
			RECT	101.825 17.708 101.857 17.772 ;
			RECT	101.993 17.708 102.025 17.772 ;
			RECT	102.123 17.724 102.155 17.756 ;
			RECT	102.245 17.729 102.277 17.761 ;
			RECT	102.375 17.708 102.407 17.772 ;
			RECT	103.795 17.708 103.827 17.772 ;
			RECT	103.925 17.729 103.957 17.761 ;
			RECT	104.047 17.724 104.079 17.756 ;
			RECT	104.177 17.708 104.209 17.772 ;
			RECT	104.345 17.708 104.377 17.772 ;
			RECT	104.513 17.708 104.545 17.772 ;
			RECT	104.681 17.708 104.713 17.772 ;
			RECT	104.849 17.708 104.881 17.772 ;
			RECT	105.017 17.708 105.049 17.772 ;
			RECT	105.185 17.708 105.217 17.772 ;
			RECT	105.353 17.708 105.385 17.772 ;
			RECT	105.521 17.708 105.553 17.772 ;
			RECT	105.689 17.708 105.721 17.772 ;
			RECT	105.857 17.708 105.889 17.772 ;
			RECT	106.025 17.708 106.057 17.772 ;
			RECT	106.193 17.708 106.225 17.772 ;
			RECT	106.361 17.708 106.393 17.772 ;
			RECT	106.529 17.708 106.561 17.772 ;
			RECT	106.697 17.708 106.729 17.772 ;
			RECT	106.865 17.708 106.897 17.772 ;
			RECT	107.033 17.708 107.065 17.772 ;
			RECT	107.201 17.708 107.233 17.772 ;
			RECT	107.369 17.708 107.401 17.772 ;
			RECT	107.537 17.708 107.569 17.772 ;
			RECT	107.705 17.708 107.737 17.772 ;
			RECT	107.873 17.708 107.905 17.772 ;
			RECT	108.041 17.708 108.073 17.772 ;
			RECT	108.209 17.708 108.241 17.772 ;
			RECT	108.377 17.708 108.409 17.772 ;
			RECT	108.545 17.708 108.577 17.772 ;
			RECT	108.713 17.708 108.745 17.772 ;
			RECT	108.881 17.708 108.913 17.772 ;
			RECT	109.049 17.708 109.081 17.772 ;
			RECT	109.217 17.708 109.249 17.772 ;
			RECT	109.385 17.708 109.417 17.772 ;
			RECT	109.553 17.708 109.585 17.772 ;
			RECT	109.721 17.708 109.753 17.772 ;
			RECT	109.889 17.708 109.921 17.772 ;
			RECT	110.057 17.708 110.089 17.772 ;
			RECT	110.225 17.708 110.257 17.772 ;
			RECT	110.393 17.708 110.425 17.772 ;
			RECT	110.561 17.708 110.593 17.772 ;
			RECT	110.729 17.708 110.761 17.772 ;
			RECT	110.897 17.708 110.929 17.772 ;
			RECT	111.065 17.708 111.097 17.772 ;
			RECT	111.233 17.708 111.265 17.772 ;
			RECT	111.401 17.708 111.433 17.772 ;
			RECT	111.569 17.708 111.601 17.772 ;
			RECT	111.737 17.708 111.769 17.772 ;
			RECT	111.905 17.708 111.937 17.772 ;
			RECT	112.073 17.708 112.105 17.772 ;
			RECT	112.241 17.708 112.273 17.772 ;
			RECT	112.409 17.708 112.441 17.772 ;
			RECT	112.577 17.708 112.609 17.772 ;
			RECT	112.745 17.708 112.777 17.772 ;
			RECT	112.913 17.708 112.945 17.772 ;
			RECT	113.081 17.708 113.113 17.772 ;
			RECT	113.249 17.708 113.281 17.772 ;
			RECT	113.417 17.708 113.449 17.772 ;
			RECT	113.585 17.708 113.617 17.772 ;
			RECT	113.753 17.708 113.785 17.772 ;
			RECT	113.921 17.708 113.953 17.772 ;
			RECT	114.089 17.708 114.121 17.772 ;
			RECT	114.257 17.708 114.289 17.772 ;
			RECT	114.425 17.708 114.457 17.772 ;
			RECT	114.593 17.708 114.625 17.772 ;
			RECT	114.761 17.708 114.793 17.772 ;
			RECT	114.929 17.708 114.961 17.772 ;
			RECT	115.097 17.708 115.129 17.772 ;
			RECT	115.265 17.708 115.297 17.772 ;
			RECT	115.433 17.708 115.465 17.772 ;
			RECT	115.601 17.708 115.633 17.772 ;
			RECT	115.769 17.708 115.801 17.772 ;
			RECT	115.937 17.708 115.969 17.772 ;
			RECT	116.105 17.708 116.137 17.772 ;
			RECT	116.273 17.708 116.305 17.772 ;
			RECT	116.441 17.708 116.473 17.772 ;
			RECT	116.609 17.708 116.641 17.772 ;
			RECT	116.777 17.708 116.809 17.772 ;
			RECT	116.945 17.708 116.977 17.772 ;
			RECT	117.113 17.708 117.145 17.772 ;
			RECT	117.281 17.708 117.313 17.772 ;
			RECT	117.449 17.708 117.481 17.772 ;
			RECT	117.617 17.708 117.649 17.772 ;
			RECT	117.785 17.708 117.817 17.772 ;
			RECT	117.953 17.708 117.985 17.772 ;
			RECT	118.121 17.708 118.153 17.772 ;
			RECT	118.289 17.708 118.321 17.772 ;
			RECT	118.457 17.708 118.489 17.772 ;
			RECT	118.625 17.708 118.657 17.772 ;
			RECT	118.793 17.708 118.825 17.772 ;
			RECT	118.961 17.708 118.993 17.772 ;
			RECT	119.129 17.708 119.161 17.772 ;
			RECT	119.297 17.708 119.329 17.772 ;
			RECT	119.465 17.708 119.497 17.772 ;
			RECT	119.633 17.708 119.665 17.772 ;
			RECT	119.801 17.708 119.833 17.772 ;
			RECT	119.969 17.708 120.001 17.772 ;
			RECT	120.137 17.708 120.169 17.772 ;
			RECT	120.305 17.708 120.337 17.772 ;
			RECT	120.473 17.708 120.505 17.772 ;
			RECT	120.641 17.708 120.673 17.772 ;
			RECT	120.809 17.708 120.841 17.772 ;
			RECT	120.977 17.708 121.009 17.772 ;
			RECT	121.145 17.708 121.177 17.772 ;
			RECT	121.313 17.708 121.345 17.772 ;
			RECT	121.481 17.708 121.513 17.772 ;
			RECT	121.649 17.708 121.681 17.772 ;
			RECT	121.817 17.708 121.849 17.772 ;
			RECT	121.985 17.708 122.017 17.772 ;
			RECT	122.153 17.708 122.185 17.772 ;
			RECT	122.321 17.708 122.353 17.772 ;
			RECT	122.489 17.708 122.521 17.772 ;
			RECT	122.657 17.708 122.689 17.772 ;
			RECT	122.825 17.708 122.857 17.772 ;
			RECT	122.993 17.708 123.025 17.772 ;
			RECT	123.161 17.708 123.193 17.772 ;
			RECT	123.329 17.708 123.361 17.772 ;
			RECT	123.497 17.708 123.529 17.772 ;
			RECT	123.665 17.708 123.697 17.772 ;
			RECT	123.833 17.708 123.865 17.772 ;
			RECT	124.001 17.708 124.033 17.772 ;
			RECT	124.169 17.708 124.201 17.772 ;
			RECT	124.337 17.708 124.369 17.772 ;
			RECT	124.505 17.708 124.537 17.772 ;
			RECT	124.673 17.708 124.705 17.772 ;
			RECT	124.841 17.708 124.873 17.772 ;
			RECT	125.009 17.708 125.041 17.772 ;
			RECT	125.177 17.708 125.209 17.772 ;
			RECT	125.345 17.708 125.377 17.772 ;
			RECT	125.513 17.708 125.545 17.772 ;
			RECT	125.681 17.708 125.713 17.772 ;
			RECT	125.849 17.708 125.881 17.772 ;
			RECT	126.017 17.708 126.049 17.772 ;
			RECT	126.185 17.708 126.217 17.772 ;
			RECT	126.353 17.708 126.385 17.772 ;
			RECT	126.521 17.708 126.553 17.772 ;
			RECT	126.689 17.708 126.721 17.772 ;
			RECT	126.857 17.708 126.889 17.772 ;
			RECT	127.025 17.708 127.057 17.772 ;
			RECT	127.193 17.708 127.225 17.772 ;
			RECT	127.361 17.708 127.393 17.772 ;
			RECT	127.529 17.708 127.561 17.772 ;
			RECT	127.697 17.708 127.729 17.772 ;
			RECT	127.865 17.708 127.897 17.772 ;
			RECT	128.033 17.708 128.065 17.772 ;
			RECT	128.201 17.708 128.233 17.772 ;
			RECT	128.369 17.708 128.401 17.772 ;
			RECT	128.537 17.708 128.569 17.772 ;
			RECT	128.705 17.708 128.737 17.772 ;
			RECT	128.873 17.708 128.905 17.772 ;
			RECT	129.041 17.708 129.073 17.772 ;
			RECT	129.209 17.708 129.241 17.772 ;
			RECT	129.377 17.708 129.409 17.772 ;
			RECT	129.545 17.708 129.577 17.772 ;
			RECT	129.713 17.708 129.745 17.772 ;
			RECT	129.881 17.708 129.913 17.772 ;
			RECT	130.049 17.708 130.081 17.772 ;
			RECT	130.217 17.708 130.249 17.772 ;
			RECT	130.385 17.708 130.417 17.772 ;
			RECT	130.553 17.708 130.585 17.772 ;
			RECT	130.721 17.708 130.753 17.772 ;
			RECT	130.889 17.708 130.921 17.772 ;
			RECT	131.057 17.708 131.089 17.772 ;
			RECT	131.225 17.708 131.257 17.772 ;
			RECT	131.393 17.708 131.425 17.772 ;
			RECT	131.561 17.708 131.593 17.772 ;
			RECT	131.729 17.708 131.761 17.772 ;
			RECT	131.897 17.708 131.929 17.772 ;
			RECT	132.065 17.708 132.097 17.772 ;
			RECT	132.233 17.708 132.265 17.772 ;
			RECT	132.401 17.708 132.433 17.772 ;
			RECT	132.569 17.708 132.601 17.772 ;
			RECT	132.737 17.708 132.769 17.772 ;
			RECT	132.905 17.708 132.937 17.772 ;
			RECT	133.073 17.708 133.105 17.772 ;
			RECT	133.241 17.708 133.273 17.772 ;
			RECT	133.409 17.708 133.441 17.772 ;
			RECT	133.577 17.708 133.609 17.772 ;
			RECT	133.745 17.708 133.777 17.772 ;
			RECT	133.913 17.708 133.945 17.772 ;
			RECT	134.081 17.708 134.113 17.772 ;
			RECT	134.249 17.708 134.281 17.772 ;
			RECT	134.417 17.708 134.449 17.772 ;
			RECT	134.585 17.708 134.617 17.772 ;
			RECT	134.753 17.708 134.785 17.772 ;
			RECT	134.921 17.708 134.953 17.772 ;
			RECT	135.089 17.708 135.121 17.772 ;
			RECT	135.257 17.708 135.289 17.772 ;
			RECT	135.425 17.708 135.457 17.772 ;
			RECT	135.593 17.708 135.625 17.772 ;
			RECT	135.761 17.708 135.793 17.772 ;
			RECT	135.929 17.708 135.961 17.772 ;
			RECT	136.097 17.708 136.129 17.772 ;
			RECT	136.265 17.708 136.297 17.772 ;
			RECT	136.433 17.708 136.465 17.772 ;
			RECT	136.601 17.708 136.633 17.772 ;
			RECT	136.769 17.708 136.801 17.772 ;
			RECT	136.937 17.708 136.969 17.772 ;
			RECT	137.105 17.708 137.137 17.772 ;
			RECT	137.273 17.708 137.305 17.772 ;
			RECT	137.441 17.708 137.473 17.772 ;
			RECT	137.609 17.708 137.641 17.772 ;
			RECT	137.777 17.708 137.809 17.772 ;
			RECT	137.945 17.708 137.977 17.772 ;
			RECT	138.113 17.708 138.145 17.772 ;
			RECT	138.281 17.708 138.313 17.772 ;
			RECT	138.449 17.708 138.481 17.772 ;
			RECT	138.617 17.708 138.649 17.772 ;
			RECT	138.785 17.708 138.817 17.772 ;
			RECT	138.953 17.708 138.985 17.772 ;
			RECT	139.121 17.708 139.153 17.772 ;
			RECT	139.289 17.708 139.321 17.772 ;
			RECT	139.457 17.708 139.489 17.772 ;
			RECT	139.625 17.708 139.657 17.772 ;
			RECT	139.793 17.708 139.825 17.772 ;
			RECT	139.961 17.708 139.993 17.772 ;
			RECT	140.129 17.708 140.161 17.772 ;
			RECT	140.297 17.708 140.329 17.772 ;
			RECT	140.465 17.708 140.497 17.772 ;
			RECT	140.633 17.708 140.665 17.772 ;
			RECT	140.801 17.708 140.833 17.772 ;
			RECT	140.969 17.708 141.001 17.772 ;
			RECT	141.137 17.708 141.169 17.772 ;
			RECT	141.305 17.708 141.337 17.772 ;
			RECT	141.473 17.708 141.505 17.772 ;
			RECT	141.641 17.708 141.673 17.772 ;
			RECT	141.809 17.708 141.841 17.772 ;
			RECT	141.977 17.708 142.009 17.772 ;
			RECT	142.145 17.708 142.177 17.772 ;
			RECT	142.313 17.708 142.345 17.772 ;
			RECT	142.481 17.708 142.513 17.772 ;
			RECT	142.649 17.708 142.681 17.772 ;
			RECT	142.817 17.708 142.849 17.772 ;
			RECT	142.985 17.708 143.017 17.772 ;
			RECT	143.153 17.708 143.185 17.772 ;
			RECT	143.321 17.708 143.353 17.772 ;
			RECT	143.489 17.708 143.521 17.772 ;
			RECT	143.657 17.708 143.689 17.772 ;
			RECT	143.825 17.708 143.857 17.772 ;
			RECT	143.993 17.708 144.025 17.772 ;
			RECT	144.161 17.708 144.193 17.772 ;
			RECT	144.329 17.708 144.361 17.772 ;
			RECT	144.497 17.708 144.529 17.772 ;
			RECT	144.665 17.708 144.697 17.772 ;
			RECT	144.833 17.708 144.865 17.772 ;
			RECT	145.001 17.708 145.033 17.772 ;
			RECT	145.169 17.708 145.201 17.772 ;
			RECT	145.337 17.708 145.369 17.772 ;
			RECT	145.505 17.708 145.537 17.772 ;
			RECT	145.673 17.708 145.705 17.772 ;
			RECT	145.841 17.708 145.873 17.772 ;
			RECT	146.009 17.708 146.041 17.772 ;
			RECT	146.177 17.708 146.209 17.772 ;
			RECT	146.345 17.708 146.377 17.772 ;
			RECT	146.513 17.708 146.545 17.772 ;
			RECT	146.681 17.708 146.713 17.772 ;
			RECT	146.849 17.708 146.881 17.772 ;
			RECT	147.017 17.708 147.049 17.772 ;
			RECT	147.185 17.708 147.217 17.772 ;
			RECT	147.316 17.724 147.348 17.756 ;
			RECT	147.437 17.724 147.469 17.756 ;
			RECT	147.567 17.708 147.599 17.772 ;
			RECT	149.879 17.708 149.911 17.772 ;
			RECT	151.13 17.708 151.194 17.772 ;
			RECT	151.81 17.708 151.842 17.772 ;
			RECT	152.249 17.708 152.281 17.772 ;
			RECT	153.56 17.708 153.624 17.772 ;
			RECT	156.601 17.708 156.633 17.772 ;
			RECT	156.731 17.724 156.763 17.756 ;
			RECT	156.852 17.724 156.884 17.756 ;
			RECT	156.983 17.708 157.015 17.772 ;
			RECT	157.151 17.708 157.183 17.772 ;
			RECT	157.319 17.708 157.351 17.772 ;
			RECT	157.487 17.708 157.519 17.772 ;
			RECT	157.655 17.708 157.687 17.772 ;
			RECT	157.823 17.708 157.855 17.772 ;
			RECT	157.991 17.708 158.023 17.772 ;
			RECT	158.159 17.708 158.191 17.772 ;
			RECT	158.327 17.708 158.359 17.772 ;
			RECT	158.495 17.708 158.527 17.772 ;
			RECT	158.663 17.708 158.695 17.772 ;
			RECT	158.831 17.708 158.863 17.772 ;
			RECT	158.999 17.708 159.031 17.772 ;
			RECT	159.167 17.708 159.199 17.772 ;
			RECT	159.335 17.708 159.367 17.772 ;
			RECT	159.503 17.708 159.535 17.772 ;
			RECT	159.671 17.708 159.703 17.772 ;
			RECT	159.839 17.708 159.871 17.772 ;
			RECT	160.007 17.708 160.039 17.772 ;
			RECT	160.175 17.708 160.207 17.772 ;
			RECT	160.343 17.708 160.375 17.772 ;
			RECT	160.511 17.708 160.543 17.772 ;
			RECT	160.679 17.708 160.711 17.772 ;
			RECT	160.847 17.708 160.879 17.772 ;
			RECT	161.015 17.708 161.047 17.772 ;
			RECT	161.183 17.708 161.215 17.772 ;
			RECT	161.351 17.708 161.383 17.772 ;
			RECT	161.519 17.708 161.551 17.772 ;
			RECT	161.687 17.708 161.719 17.772 ;
			RECT	161.855 17.708 161.887 17.772 ;
			RECT	162.023 17.708 162.055 17.772 ;
			RECT	162.191 17.708 162.223 17.772 ;
			RECT	162.359 17.708 162.391 17.772 ;
			RECT	162.527 17.708 162.559 17.772 ;
			RECT	162.695 17.708 162.727 17.772 ;
			RECT	162.863 17.708 162.895 17.772 ;
			RECT	163.031 17.708 163.063 17.772 ;
			RECT	163.199 17.708 163.231 17.772 ;
			RECT	163.367 17.708 163.399 17.772 ;
			RECT	163.535 17.708 163.567 17.772 ;
			RECT	163.703 17.708 163.735 17.772 ;
			RECT	163.871 17.708 163.903 17.772 ;
			RECT	164.039 17.708 164.071 17.772 ;
			RECT	164.207 17.708 164.239 17.772 ;
			RECT	164.375 17.708 164.407 17.772 ;
			RECT	164.543 17.708 164.575 17.772 ;
			RECT	164.711 17.708 164.743 17.772 ;
			RECT	164.879 17.708 164.911 17.772 ;
			RECT	165.047 17.708 165.079 17.772 ;
			RECT	165.215 17.708 165.247 17.772 ;
			RECT	165.383 17.708 165.415 17.772 ;
			RECT	165.551 17.708 165.583 17.772 ;
			RECT	165.719 17.708 165.751 17.772 ;
			RECT	165.887 17.708 165.919 17.772 ;
			RECT	166.055 17.708 166.087 17.772 ;
			RECT	166.223 17.708 166.255 17.772 ;
			RECT	166.391 17.708 166.423 17.772 ;
			RECT	166.559 17.708 166.591 17.772 ;
			RECT	166.727 17.708 166.759 17.772 ;
			RECT	166.895 17.708 166.927 17.772 ;
			RECT	167.063 17.708 167.095 17.772 ;
			RECT	167.231 17.708 167.263 17.772 ;
			RECT	167.399 17.708 167.431 17.772 ;
			RECT	167.567 17.708 167.599 17.772 ;
			RECT	167.735 17.708 167.767 17.772 ;
			RECT	167.903 17.708 167.935 17.772 ;
			RECT	168.071 17.708 168.103 17.772 ;
			RECT	168.239 17.708 168.271 17.772 ;
			RECT	168.407 17.708 168.439 17.772 ;
			RECT	168.575 17.708 168.607 17.772 ;
			RECT	168.743 17.708 168.775 17.772 ;
			RECT	168.911 17.708 168.943 17.772 ;
			RECT	169.079 17.708 169.111 17.772 ;
			RECT	169.247 17.708 169.279 17.772 ;
			RECT	169.415 17.708 169.447 17.772 ;
			RECT	169.583 17.708 169.615 17.772 ;
			RECT	169.751 17.708 169.783 17.772 ;
			RECT	169.919 17.708 169.951 17.772 ;
			RECT	170.087 17.708 170.119 17.772 ;
			RECT	170.255 17.708 170.287 17.772 ;
			RECT	170.423 17.708 170.455 17.772 ;
			RECT	170.591 17.708 170.623 17.772 ;
			RECT	170.759 17.708 170.791 17.772 ;
			RECT	170.927 17.708 170.959 17.772 ;
			RECT	171.095 17.708 171.127 17.772 ;
			RECT	171.263 17.708 171.295 17.772 ;
			RECT	171.431 17.708 171.463 17.772 ;
			RECT	171.599 17.708 171.631 17.772 ;
			RECT	171.767 17.708 171.799 17.772 ;
			RECT	171.935 17.708 171.967 17.772 ;
			RECT	172.103 17.708 172.135 17.772 ;
			RECT	172.271 17.708 172.303 17.772 ;
			RECT	172.439 17.708 172.471 17.772 ;
			RECT	172.607 17.708 172.639 17.772 ;
			RECT	172.775 17.708 172.807 17.772 ;
			RECT	172.943 17.708 172.975 17.772 ;
			RECT	173.111 17.708 173.143 17.772 ;
			RECT	173.279 17.708 173.311 17.772 ;
			RECT	173.447 17.708 173.479 17.772 ;
			RECT	173.615 17.708 173.647 17.772 ;
			RECT	173.783 17.708 173.815 17.772 ;
			RECT	173.951 17.708 173.983 17.772 ;
			RECT	174.119 17.708 174.151 17.772 ;
			RECT	174.287 17.708 174.319 17.772 ;
			RECT	174.455 17.708 174.487 17.772 ;
			RECT	174.623 17.708 174.655 17.772 ;
			RECT	174.791 17.708 174.823 17.772 ;
			RECT	174.959 17.708 174.991 17.772 ;
			RECT	175.127 17.708 175.159 17.772 ;
			RECT	175.295 17.708 175.327 17.772 ;
			RECT	175.463 17.708 175.495 17.772 ;
			RECT	175.631 17.708 175.663 17.772 ;
			RECT	175.799 17.708 175.831 17.772 ;
			RECT	175.967 17.708 175.999 17.772 ;
			RECT	176.135 17.708 176.167 17.772 ;
			RECT	176.303 17.708 176.335 17.772 ;
			RECT	176.471 17.708 176.503 17.772 ;
			RECT	176.639 17.708 176.671 17.772 ;
			RECT	176.807 17.708 176.839 17.772 ;
			RECT	176.975 17.708 177.007 17.772 ;
			RECT	177.143 17.708 177.175 17.772 ;
			RECT	177.311 17.708 177.343 17.772 ;
			RECT	177.479 17.708 177.511 17.772 ;
			RECT	177.647 17.708 177.679 17.772 ;
			RECT	177.815 17.708 177.847 17.772 ;
			RECT	177.983 17.708 178.015 17.772 ;
			RECT	178.151 17.708 178.183 17.772 ;
			RECT	178.319 17.708 178.351 17.772 ;
			RECT	178.487 17.708 178.519 17.772 ;
			RECT	178.655 17.708 178.687 17.772 ;
			RECT	178.823 17.708 178.855 17.772 ;
			RECT	178.991 17.708 179.023 17.772 ;
			RECT	179.159 17.708 179.191 17.772 ;
			RECT	179.327 17.708 179.359 17.772 ;
			RECT	179.495 17.708 179.527 17.772 ;
			RECT	179.663 17.708 179.695 17.772 ;
			RECT	179.831 17.708 179.863 17.772 ;
			RECT	179.999 17.708 180.031 17.772 ;
			RECT	180.167 17.708 180.199 17.772 ;
			RECT	180.335 17.708 180.367 17.772 ;
			RECT	180.503 17.708 180.535 17.772 ;
			RECT	180.671 17.708 180.703 17.772 ;
			RECT	180.839 17.708 180.871 17.772 ;
			RECT	181.007 17.708 181.039 17.772 ;
			RECT	181.175 17.708 181.207 17.772 ;
			RECT	181.343 17.708 181.375 17.772 ;
			RECT	181.511 17.708 181.543 17.772 ;
			RECT	181.679 17.708 181.711 17.772 ;
			RECT	181.847 17.708 181.879 17.772 ;
			RECT	182.015 17.708 182.047 17.772 ;
			RECT	182.183 17.708 182.215 17.772 ;
			RECT	182.351 17.708 182.383 17.772 ;
			RECT	182.519 17.708 182.551 17.772 ;
			RECT	182.687 17.708 182.719 17.772 ;
			RECT	182.855 17.708 182.887 17.772 ;
			RECT	183.023 17.708 183.055 17.772 ;
			RECT	183.191 17.708 183.223 17.772 ;
			RECT	183.359 17.708 183.391 17.772 ;
			RECT	183.527 17.708 183.559 17.772 ;
			RECT	183.695 17.708 183.727 17.772 ;
			RECT	183.863 17.708 183.895 17.772 ;
			RECT	184.031 17.708 184.063 17.772 ;
			RECT	184.199 17.708 184.231 17.772 ;
			RECT	184.367 17.708 184.399 17.772 ;
			RECT	184.535 17.708 184.567 17.772 ;
			RECT	184.703 17.708 184.735 17.772 ;
			RECT	184.871 17.708 184.903 17.772 ;
			RECT	185.039 17.708 185.071 17.772 ;
			RECT	185.207 17.708 185.239 17.772 ;
			RECT	185.375 17.708 185.407 17.772 ;
			RECT	185.543 17.708 185.575 17.772 ;
			RECT	185.711 17.708 185.743 17.772 ;
			RECT	185.879 17.708 185.911 17.772 ;
			RECT	186.047 17.708 186.079 17.772 ;
			RECT	186.215 17.708 186.247 17.772 ;
			RECT	186.383 17.708 186.415 17.772 ;
			RECT	186.551 17.708 186.583 17.772 ;
			RECT	186.719 17.708 186.751 17.772 ;
			RECT	186.887 17.708 186.919 17.772 ;
			RECT	187.055 17.708 187.087 17.772 ;
			RECT	187.223 17.708 187.255 17.772 ;
			RECT	187.391 17.708 187.423 17.772 ;
			RECT	187.559 17.708 187.591 17.772 ;
			RECT	187.727 17.708 187.759 17.772 ;
			RECT	187.895 17.708 187.927 17.772 ;
			RECT	188.063 17.708 188.095 17.772 ;
			RECT	188.231 17.708 188.263 17.772 ;
			RECT	188.399 17.708 188.431 17.772 ;
			RECT	188.567 17.708 188.599 17.772 ;
			RECT	188.735 17.708 188.767 17.772 ;
			RECT	188.903 17.708 188.935 17.772 ;
			RECT	189.071 17.708 189.103 17.772 ;
			RECT	189.239 17.708 189.271 17.772 ;
			RECT	189.407 17.708 189.439 17.772 ;
			RECT	189.575 17.708 189.607 17.772 ;
			RECT	189.743 17.708 189.775 17.772 ;
			RECT	189.911 17.708 189.943 17.772 ;
			RECT	190.079 17.708 190.111 17.772 ;
			RECT	190.247 17.708 190.279 17.772 ;
			RECT	190.415 17.708 190.447 17.772 ;
			RECT	190.583 17.708 190.615 17.772 ;
			RECT	190.751 17.708 190.783 17.772 ;
			RECT	190.919 17.708 190.951 17.772 ;
			RECT	191.087 17.708 191.119 17.772 ;
			RECT	191.255 17.708 191.287 17.772 ;
			RECT	191.423 17.708 191.455 17.772 ;
			RECT	191.591 17.708 191.623 17.772 ;
			RECT	191.759 17.708 191.791 17.772 ;
			RECT	191.927 17.708 191.959 17.772 ;
			RECT	192.095 17.708 192.127 17.772 ;
			RECT	192.263 17.708 192.295 17.772 ;
			RECT	192.431 17.708 192.463 17.772 ;
			RECT	192.599 17.708 192.631 17.772 ;
			RECT	192.767 17.708 192.799 17.772 ;
			RECT	192.935 17.708 192.967 17.772 ;
			RECT	193.103 17.708 193.135 17.772 ;
			RECT	193.271 17.708 193.303 17.772 ;
			RECT	193.439 17.708 193.471 17.772 ;
			RECT	193.607 17.708 193.639 17.772 ;
			RECT	193.775 17.708 193.807 17.772 ;
			RECT	193.943 17.708 193.975 17.772 ;
			RECT	194.111 17.708 194.143 17.772 ;
			RECT	194.279 17.708 194.311 17.772 ;
			RECT	194.447 17.708 194.479 17.772 ;
			RECT	194.615 17.708 194.647 17.772 ;
			RECT	194.783 17.708 194.815 17.772 ;
			RECT	194.951 17.708 194.983 17.772 ;
			RECT	195.119 17.708 195.151 17.772 ;
			RECT	195.287 17.708 195.319 17.772 ;
			RECT	195.455 17.708 195.487 17.772 ;
			RECT	195.623 17.708 195.655 17.772 ;
			RECT	195.791 17.708 195.823 17.772 ;
			RECT	195.959 17.708 195.991 17.772 ;
			RECT	196.127 17.708 196.159 17.772 ;
			RECT	196.295 17.708 196.327 17.772 ;
			RECT	196.463 17.708 196.495 17.772 ;
			RECT	196.631 17.708 196.663 17.772 ;
			RECT	196.799 17.708 196.831 17.772 ;
			RECT	196.967 17.708 196.999 17.772 ;
			RECT	197.135 17.708 197.167 17.772 ;
			RECT	197.303 17.708 197.335 17.772 ;
			RECT	197.471 17.708 197.503 17.772 ;
			RECT	197.639 17.708 197.671 17.772 ;
			RECT	197.807 17.708 197.839 17.772 ;
			RECT	197.975 17.708 198.007 17.772 ;
			RECT	198.143 17.708 198.175 17.772 ;
			RECT	198.311 17.708 198.343 17.772 ;
			RECT	198.479 17.708 198.511 17.772 ;
			RECT	198.647 17.708 198.679 17.772 ;
			RECT	198.815 17.708 198.847 17.772 ;
			RECT	198.983 17.708 199.015 17.772 ;
			RECT	199.151 17.708 199.183 17.772 ;
			RECT	199.319 17.708 199.351 17.772 ;
			RECT	199.487 17.708 199.519 17.772 ;
			RECT	199.655 17.708 199.687 17.772 ;
			RECT	199.823 17.708 199.855 17.772 ;
			RECT	199.991 17.708 200.023 17.772 ;
			RECT	200.121 17.724 200.153 17.756 ;
			RECT	200.243 17.729 200.275 17.761 ;
			RECT	200.373 17.708 200.405 17.772 ;
			RECT	200.9 17.708 200.932 17.772 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 15.76 201.665 15.88 ;
			LAYER	J3 ;
			RECT	0.755 15.788 0.787 15.852 ;
			RECT	1.645 15.788 1.709 15.852 ;
			RECT	2.323 15.788 2.387 15.852 ;
			RECT	3.438 15.788 3.47 15.852 ;
			RECT	3.585 15.788 3.617 15.852 ;
			RECT	4.195 15.788 4.227 15.852 ;
			RECT	4.72 15.788 4.752 15.852 ;
			RECT	4.944 15.788 5.008 15.852 ;
			RECT	5.267 15.788 5.299 15.852 ;
			RECT	5.797 15.788 5.829 15.852 ;
			RECT	5.927 15.809 5.959 15.841 ;
			RECT	6.049 15.804 6.081 15.836 ;
			RECT	6.179 15.788 6.211 15.852 ;
			RECT	6.347 15.788 6.379 15.852 ;
			RECT	6.515 15.788 6.547 15.852 ;
			RECT	6.683 15.788 6.715 15.852 ;
			RECT	6.851 15.788 6.883 15.852 ;
			RECT	7.019 15.788 7.051 15.852 ;
			RECT	7.187 15.788 7.219 15.852 ;
			RECT	7.355 15.788 7.387 15.852 ;
			RECT	7.523 15.788 7.555 15.852 ;
			RECT	7.691 15.788 7.723 15.852 ;
			RECT	7.859 15.788 7.891 15.852 ;
			RECT	8.027 15.788 8.059 15.852 ;
			RECT	8.195 15.788 8.227 15.852 ;
			RECT	8.363 15.788 8.395 15.852 ;
			RECT	8.531 15.788 8.563 15.852 ;
			RECT	8.699 15.788 8.731 15.852 ;
			RECT	8.867 15.788 8.899 15.852 ;
			RECT	9.035 15.788 9.067 15.852 ;
			RECT	9.203 15.788 9.235 15.852 ;
			RECT	9.371 15.788 9.403 15.852 ;
			RECT	9.539 15.788 9.571 15.852 ;
			RECT	9.707 15.788 9.739 15.852 ;
			RECT	9.875 15.788 9.907 15.852 ;
			RECT	10.043 15.788 10.075 15.852 ;
			RECT	10.211 15.788 10.243 15.852 ;
			RECT	10.379 15.788 10.411 15.852 ;
			RECT	10.547 15.788 10.579 15.852 ;
			RECT	10.715 15.788 10.747 15.852 ;
			RECT	10.883 15.788 10.915 15.852 ;
			RECT	11.051 15.788 11.083 15.852 ;
			RECT	11.219 15.788 11.251 15.852 ;
			RECT	11.387 15.788 11.419 15.852 ;
			RECT	11.555 15.788 11.587 15.852 ;
			RECT	11.723 15.788 11.755 15.852 ;
			RECT	11.891 15.788 11.923 15.852 ;
			RECT	12.059 15.788 12.091 15.852 ;
			RECT	12.227 15.788 12.259 15.852 ;
			RECT	12.395 15.788 12.427 15.852 ;
			RECT	12.563 15.788 12.595 15.852 ;
			RECT	12.731 15.788 12.763 15.852 ;
			RECT	12.899 15.788 12.931 15.852 ;
			RECT	13.067 15.788 13.099 15.852 ;
			RECT	13.235 15.788 13.267 15.852 ;
			RECT	13.403 15.788 13.435 15.852 ;
			RECT	13.571 15.788 13.603 15.852 ;
			RECT	13.739 15.788 13.771 15.852 ;
			RECT	13.907 15.788 13.939 15.852 ;
			RECT	14.075 15.788 14.107 15.852 ;
			RECT	14.243 15.788 14.275 15.852 ;
			RECT	14.411 15.788 14.443 15.852 ;
			RECT	14.579 15.788 14.611 15.852 ;
			RECT	14.747 15.788 14.779 15.852 ;
			RECT	14.915 15.788 14.947 15.852 ;
			RECT	15.083 15.788 15.115 15.852 ;
			RECT	15.251 15.788 15.283 15.852 ;
			RECT	15.419 15.788 15.451 15.852 ;
			RECT	15.587 15.788 15.619 15.852 ;
			RECT	15.755 15.788 15.787 15.852 ;
			RECT	15.923 15.788 15.955 15.852 ;
			RECT	16.091 15.788 16.123 15.852 ;
			RECT	16.259 15.788 16.291 15.852 ;
			RECT	16.427 15.788 16.459 15.852 ;
			RECT	16.595 15.788 16.627 15.852 ;
			RECT	16.763 15.788 16.795 15.852 ;
			RECT	16.931 15.788 16.963 15.852 ;
			RECT	17.099 15.788 17.131 15.852 ;
			RECT	17.267 15.788 17.299 15.852 ;
			RECT	17.435 15.788 17.467 15.852 ;
			RECT	17.603 15.788 17.635 15.852 ;
			RECT	17.771 15.788 17.803 15.852 ;
			RECT	17.939 15.788 17.971 15.852 ;
			RECT	18.107 15.788 18.139 15.852 ;
			RECT	18.275 15.788 18.307 15.852 ;
			RECT	18.443 15.788 18.475 15.852 ;
			RECT	18.611 15.788 18.643 15.852 ;
			RECT	18.779 15.788 18.811 15.852 ;
			RECT	18.947 15.788 18.979 15.852 ;
			RECT	19.115 15.788 19.147 15.852 ;
			RECT	19.283 15.788 19.315 15.852 ;
			RECT	19.451 15.788 19.483 15.852 ;
			RECT	19.619 15.788 19.651 15.852 ;
			RECT	19.787 15.788 19.819 15.852 ;
			RECT	19.955 15.788 19.987 15.852 ;
			RECT	20.123 15.788 20.155 15.852 ;
			RECT	20.291 15.788 20.323 15.852 ;
			RECT	20.459 15.788 20.491 15.852 ;
			RECT	20.627 15.788 20.659 15.852 ;
			RECT	20.795 15.788 20.827 15.852 ;
			RECT	20.963 15.788 20.995 15.852 ;
			RECT	21.131 15.788 21.163 15.852 ;
			RECT	21.299 15.788 21.331 15.852 ;
			RECT	21.467 15.788 21.499 15.852 ;
			RECT	21.635 15.788 21.667 15.852 ;
			RECT	21.803 15.788 21.835 15.852 ;
			RECT	21.971 15.788 22.003 15.852 ;
			RECT	22.139 15.788 22.171 15.852 ;
			RECT	22.307 15.788 22.339 15.852 ;
			RECT	22.475 15.788 22.507 15.852 ;
			RECT	22.643 15.788 22.675 15.852 ;
			RECT	22.811 15.788 22.843 15.852 ;
			RECT	22.979 15.788 23.011 15.852 ;
			RECT	23.147 15.788 23.179 15.852 ;
			RECT	23.315 15.788 23.347 15.852 ;
			RECT	23.483 15.788 23.515 15.852 ;
			RECT	23.651 15.788 23.683 15.852 ;
			RECT	23.819 15.788 23.851 15.852 ;
			RECT	23.987 15.788 24.019 15.852 ;
			RECT	24.155 15.788 24.187 15.852 ;
			RECT	24.323 15.788 24.355 15.852 ;
			RECT	24.491 15.788 24.523 15.852 ;
			RECT	24.659 15.788 24.691 15.852 ;
			RECT	24.827 15.788 24.859 15.852 ;
			RECT	24.995 15.788 25.027 15.852 ;
			RECT	25.163 15.788 25.195 15.852 ;
			RECT	25.331 15.788 25.363 15.852 ;
			RECT	25.499 15.788 25.531 15.852 ;
			RECT	25.667 15.788 25.699 15.852 ;
			RECT	25.835 15.788 25.867 15.852 ;
			RECT	26.003 15.788 26.035 15.852 ;
			RECT	26.171 15.788 26.203 15.852 ;
			RECT	26.339 15.788 26.371 15.852 ;
			RECT	26.507 15.788 26.539 15.852 ;
			RECT	26.675 15.788 26.707 15.852 ;
			RECT	26.843 15.788 26.875 15.852 ;
			RECT	27.011 15.788 27.043 15.852 ;
			RECT	27.179 15.788 27.211 15.852 ;
			RECT	27.347 15.788 27.379 15.852 ;
			RECT	27.515 15.788 27.547 15.852 ;
			RECT	27.683 15.788 27.715 15.852 ;
			RECT	27.851 15.788 27.883 15.852 ;
			RECT	28.019 15.788 28.051 15.852 ;
			RECT	28.187 15.788 28.219 15.852 ;
			RECT	28.355 15.788 28.387 15.852 ;
			RECT	28.523 15.788 28.555 15.852 ;
			RECT	28.691 15.788 28.723 15.852 ;
			RECT	28.859 15.788 28.891 15.852 ;
			RECT	29.027 15.788 29.059 15.852 ;
			RECT	29.195 15.788 29.227 15.852 ;
			RECT	29.363 15.788 29.395 15.852 ;
			RECT	29.531 15.788 29.563 15.852 ;
			RECT	29.699 15.788 29.731 15.852 ;
			RECT	29.867 15.788 29.899 15.852 ;
			RECT	30.035 15.788 30.067 15.852 ;
			RECT	30.203 15.788 30.235 15.852 ;
			RECT	30.371 15.788 30.403 15.852 ;
			RECT	30.539 15.788 30.571 15.852 ;
			RECT	30.707 15.788 30.739 15.852 ;
			RECT	30.875 15.788 30.907 15.852 ;
			RECT	31.043 15.788 31.075 15.852 ;
			RECT	31.211 15.788 31.243 15.852 ;
			RECT	31.379 15.788 31.411 15.852 ;
			RECT	31.547 15.788 31.579 15.852 ;
			RECT	31.715 15.788 31.747 15.852 ;
			RECT	31.883 15.788 31.915 15.852 ;
			RECT	32.051 15.788 32.083 15.852 ;
			RECT	32.219 15.788 32.251 15.852 ;
			RECT	32.387 15.788 32.419 15.852 ;
			RECT	32.555 15.788 32.587 15.852 ;
			RECT	32.723 15.788 32.755 15.852 ;
			RECT	32.891 15.788 32.923 15.852 ;
			RECT	33.059 15.788 33.091 15.852 ;
			RECT	33.227 15.788 33.259 15.852 ;
			RECT	33.395 15.788 33.427 15.852 ;
			RECT	33.563 15.788 33.595 15.852 ;
			RECT	33.731 15.788 33.763 15.852 ;
			RECT	33.899 15.788 33.931 15.852 ;
			RECT	34.067 15.788 34.099 15.852 ;
			RECT	34.235 15.788 34.267 15.852 ;
			RECT	34.403 15.788 34.435 15.852 ;
			RECT	34.571 15.788 34.603 15.852 ;
			RECT	34.739 15.788 34.771 15.852 ;
			RECT	34.907 15.788 34.939 15.852 ;
			RECT	35.075 15.788 35.107 15.852 ;
			RECT	35.243 15.788 35.275 15.852 ;
			RECT	35.411 15.788 35.443 15.852 ;
			RECT	35.579 15.788 35.611 15.852 ;
			RECT	35.747 15.788 35.779 15.852 ;
			RECT	35.915 15.788 35.947 15.852 ;
			RECT	36.083 15.788 36.115 15.852 ;
			RECT	36.251 15.788 36.283 15.852 ;
			RECT	36.419 15.788 36.451 15.852 ;
			RECT	36.587 15.788 36.619 15.852 ;
			RECT	36.755 15.788 36.787 15.852 ;
			RECT	36.923 15.788 36.955 15.852 ;
			RECT	37.091 15.788 37.123 15.852 ;
			RECT	37.259 15.788 37.291 15.852 ;
			RECT	37.427 15.788 37.459 15.852 ;
			RECT	37.595 15.788 37.627 15.852 ;
			RECT	37.763 15.788 37.795 15.852 ;
			RECT	37.931 15.788 37.963 15.852 ;
			RECT	38.099 15.788 38.131 15.852 ;
			RECT	38.267 15.788 38.299 15.852 ;
			RECT	38.435 15.788 38.467 15.852 ;
			RECT	38.603 15.788 38.635 15.852 ;
			RECT	38.771 15.788 38.803 15.852 ;
			RECT	38.939 15.788 38.971 15.852 ;
			RECT	39.107 15.788 39.139 15.852 ;
			RECT	39.275 15.788 39.307 15.852 ;
			RECT	39.443 15.788 39.475 15.852 ;
			RECT	39.611 15.788 39.643 15.852 ;
			RECT	39.779 15.788 39.811 15.852 ;
			RECT	39.947 15.788 39.979 15.852 ;
			RECT	40.115 15.788 40.147 15.852 ;
			RECT	40.283 15.788 40.315 15.852 ;
			RECT	40.451 15.788 40.483 15.852 ;
			RECT	40.619 15.788 40.651 15.852 ;
			RECT	40.787 15.788 40.819 15.852 ;
			RECT	40.955 15.788 40.987 15.852 ;
			RECT	41.123 15.788 41.155 15.852 ;
			RECT	41.291 15.788 41.323 15.852 ;
			RECT	41.459 15.788 41.491 15.852 ;
			RECT	41.627 15.788 41.659 15.852 ;
			RECT	41.795 15.788 41.827 15.852 ;
			RECT	41.963 15.788 41.995 15.852 ;
			RECT	42.131 15.788 42.163 15.852 ;
			RECT	42.299 15.788 42.331 15.852 ;
			RECT	42.467 15.788 42.499 15.852 ;
			RECT	42.635 15.788 42.667 15.852 ;
			RECT	42.803 15.788 42.835 15.852 ;
			RECT	42.971 15.788 43.003 15.852 ;
			RECT	43.139 15.788 43.171 15.852 ;
			RECT	43.307 15.788 43.339 15.852 ;
			RECT	43.475 15.788 43.507 15.852 ;
			RECT	43.643 15.788 43.675 15.852 ;
			RECT	43.811 15.788 43.843 15.852 ;
			RECT	43.979 15.788 44.011 15.852 ;
			RECT	44.147 15.788 44.179 15.852 ;
			RECT	44.315 15.788 44.347 15.852 ;
			RECT	44.483 15.788 44.515 15.852 ;
			RECT	44.651 15.788 44.683 15.852 ;
			RECT	44.819 15.788 44.851 15.852 ;
			RECT	44.987 15.788 45.019 15.852 ;
			RECT	45.155 15.788 45.187 15.852 ;
			RECT	45.323 15.788 45.355 15.852 ;
			RECT	45.491 15.788 45.523 15.852 ;
			RECT	45.659 15.788 45.691 15.852 ;
			RECT	45.827 15.788 45.859 15.852 ;
			RECT	45.995 15.788 46.027 15.852 ;
			RECT	46.163 15.788 46.195 15.852 ;
			RECT	46.331 15.788 46.363 15.852 ;
			RECT	46.499 15.788 46.531 15.852 ;
			RECT	46.667 15.788 46.699 15.852 ;
			RECT	46.835 15.788 46.867 15.852 ;
			RECT	47.003 15.788 47.035 15.852 ;
			RECT	47.171 15.788 47.203 15.852 ;
			RECT	47.339 15.788 47.371 15.852 ;
			RECT	47.507 15.788 47.539 15.852 ;
			RECT	47.675 15.788 47.707 15.852 ;
			RECT	47.843 15.788 47.875 15.852 ;
			RECT	48.011 15.788 48.043 15.852 ;
			RECT	48.179 15.788 48.211 15.852 ;
			RECT	48.347 15.788 48.379 15.852 ;
			RECT	48.515 15.788 48.547 15.852 ;
			RECT	48.683 15.788 48.715 15.852 ;
			RECT	48.851 15.788 48.883 15.852 ;
			RECT	49.019 15.788 49.051 15.852 ;
			RECT	49.187 15.788 49.219 15.852 ;
			RECT	49.318 15.804 49.35 15.836 ;
			RECT	49.439 15.804 49.471 15.836 ;
			RECT	49.569 15.788 49.601 15.852 ;
			RECT	51.881 15.788 51.913 15.852 ;
			RECT	53.132 15.788 53.196 15.852 ;
			RECT	53.812 15.788 53.844 15.852 ;
			RECT	54.251 15.788 54.283 15.852 ;
			RECT	55.562 15.788 55.626 15.852 ;
			RECT	58.603 15.788 58.635 15.852 ;
			RECT	58.733 15.804 58.765 15.836 ;
			RECT	58.854 15.804 58.886 15.836 ;
			RECT	58.985 15.788 59.017 15.852 ;
			RECT	59.153 15.788 59.185 15.852 ;
			RECT	59.321 15.788 59.353 15.852 ;
			RECT	59.489 15.788 59.521 15.852 ;
			RECT	59.657 15.788 59.689 15.852 ;
			RECT	59.825 15.788 59.857 15.852 ;
			RECT	59.993 15.788 60.025 15.852 ;
			RECT	60.161 15.788 60.193 15.852 ;
			RECT	60.329 15.788 60.361 15.852 ;
			RECT	60.497 15.788 60.529 15.852 ;
			RECT	60.665 15.788 60.697 15.852 ;
			RECT	60.833 15.788 60.865 15.852 ;
			RECT	61.001 15.788 61.033 15.852 ;
			RECT	61.169 15.788 61.201 15.852 ;
			RECT	61.337 15.788 61.369 15.852 ;
			RECT	61.505 15.788 61.537 15.852 ;
			RECT	61.673 15.788 61.705 15.852 ;
			RECT	61.841 15.788 61.873 15.852 ;
			RECT	62.009 15.788 62.041 15.852 ;
			RECT	62.177 15.788 62.209 15.852 ;
			RECT	62.345 15.788 62.377 15.852 ;
			RECT	62.513 15.788 62.545 15.852 ;
			RECT	62.681 15.788 62.713 15.852 ;
			RECT	62.849 15.788 62.881 15.852 ;
			RECT	63.017 15.788 63.049 15.852 ;
			RECT	63.185 15.788 63.217 15.852 ;
			RECT	63.353 15.788 63.385 15.852 ;
			RECT	63.521 15.788 63.553 15.852 ;
			RECT	63.689 15.788 63.721 15.852 ;
			RECT	63.857 15.788 63.889 15.852 ;
			RECT	64.025 15.788 64.057 15.852 ;
			RECT	64.193 15.788 64.225 15.852 ;
			RECT	64.361 15.788 64.393 15.852 ;
			RECT	64.529 15.788 64.561 15.852 ;
			RECT	64.697 15.788 64.729 15.852 ;
			RECT	64.865 15.788 64.897 15.852 ;
			RECT	65.033 15.788 65.065 15.852 ;
			RECT	65.201 15.788 65.233 15.852 ;
			RECT	65.369 15.788 65.401 15.852 ;
			RECT	65.537 15.788 65.569 15.852 ;
			RECT	65.705 15.788 65.737 15.852 ;
			RECT	65.873 15.788 65.905 15.852 ;
			RECT	66.041 15.788 66.073 15.852 ;
			RECT	66.209 15.788 66.241 15.852 ;
			RECT	66.377 15.788 66.409 15.852 ;
			RECT	66.545 15.788 66.577 15.852 ;
			RECT	66.713 15.788 66.745 15.852 ;
			RECT	66.881 15.788 66.913 15.852 ;
			RECT	67.049 15.788 67.081 15.852 ;
			RECT	67.217 15.788 67.249 15.852 ;
			RECT	67.385 15.788 67.417 15.852 ;
			RECT	67.553 15.788 67.585 15.852 ;
			RECT	67.721 15.788 67.753 15.852 ;
			RECT	67.889 15.788 67.921 15.852 ;
			RECT	68.057 15.788 68.089 15.852 ;
			RECT	68.225 15.788 68.257 15.852 ;
			RECT	68.393 15.788 68.425 15.852 ;
			RECT	68.561 15.788 68.593 15.852 ;
			RECT	68.729 15.788 68.761 15.852 ;
			RECT	68.897 15.788 68.929 15.852 ;
			RECT	69.065 15.788 69.097 15.852 ;
			RECT	69.233 15.788 69.265 15.852 ;
			RECT	69.401 15.788 69.433 15.852 ;
			RECT	69.569 15.788 69.601 15.852 ;
			RECT	69.737 15.788 69.769 15.852 ;
			RECT	69.905 15.788 69.937 15.852 ;
			RECT	70.073 15.788 70.105 15.852 ;
			RECT	70.241 15.788 70.273 15.852 ;
			RECT	70.409 15.788 70.441 15.852 ;
			RECT	70.577 15.788 70.609 15.852 ;
			RECT	70.745 15.788 70.777 15.852 ;
			RECT	70.913 15.788 70.945 15.852 ;
			RECT	71.081 15.788 71.113 15.852 ;
			RECT	71.249 15.788 71.281 15.852 ;
			RECT	71.417 15.788 71.449 15.852 ;
			RECT	71.585 15.788 71.617 15.852 ;
			RECT	71.753 15.788 71.785 15.852 ;
			RECT	71.921 15.788 71.953 15.852 ;
			RECT	72.089 15.788 72.121 15.852 ;
			RECT	72.257 15.788 72.289 15.852 ;
			RECT	72.425 15.788 72.457 15.852 ;
			RECT	72.593 15.788 72.625 15.852 ;
			RECT	72.761 15.788 72.793 15.852 ;
			RECT	72.929 15.788 72.961 15.852 ;
			RECT	73.097 15.788 73.129 15.852 ;
			RECT	73.265 15.788 73.297 15.852 ;
			RECT	73.433 15.788 73.465 15.852 ;
			RECT	73.601 15.788 73.633 15.852 ;
			RECT	73.769 15.788 73.801 15.852 ;
			RECT	73.937 15.788 73.969 15.852 ;
			RECT	74.105 15.788 74.137 15.852 ;
			RECT	74.273 15.788 74.305 15.852 ;
			RECT	74.441 15.788 74.473 15.852 ;
			RECT	74.609 15.788 74.641 15.852 ;
			RECT	74.777 15.788 74.809 15.852 ;
			RECT	74.945 15.788 74.977 15.852 ;
			RECT	75.113 15.788 75.145 15.852 ;
			RECT	75.281 15.788 75.313 15.852 ;
			RECT	75.449 15.788 75.481 15.852 ;
			RECT	75.617 15.788 75.649 15.852 ;
			RECT	75.785 15.788 75.817 15.852 ;
			RECT	75.953 15.788 75.985 15.852 ;
			RECT	76.121 15.788 76.153 15.852 ;
			RECT	76.289 15.788 76.321 15.852 ;
			RECT	76.457 15.788 76.489 15.852 ;
			RECT	76.625 15.788 76.657 15.852 ;
			RECT	76.793 15.788 76.825 15.852 ;
			RECT	76.961 15.788 76.993 15.852 ;
			RECT	77.129 15.788 77.161 15.852 ;
			RECT	77.297 15.788 77.329 15.852 ;
			RECT	77.465 15.788 77.497 15.852 ;
			RECT	77.633 15.788 77.665 15.852 ;
			RECT	77.801 15.788 77.833 15.852 ;
			RECT	77.969 15.788 78.001 15.852 ;
			RECT	78.137 15.788 78.169 15.852 ;
			RECT	78.305 15.788 78.337 15.852 ;
			RECT	78.473 15.788 78.505 15.852 ;
			RECT	78.641 15.788 78.673 15.852 ;
			RECT	78.809 15.788 78.841 15.852 ;
			RECT	78.977 15.788 79.009 15.852 ;
			RECT	79.145 15.788 79.177 15.852 ;
			RECT	79.313 15.788 79.345 15.852 ;
			RECT	79.481 15.788 79.513 15.852 ;
			RECT	79.649 15.788 79.681 15.852 ;
			RECT	79.817 15.788 79.849 15.852 ;
			RECT	79.985 15.788 80.017 15.852 ;
			RECT	80.153 15.788 80.185 15.852 ;
			RECT	80.321 15.788 80.353 15.852 ;
			RECT	80.489 15.788 80.521 15.852 ;
			RECT	80.657 15.788 80.689 15.852 ;
			RECT	80.825 15.788 80.857 15.852 ;
			RECT	80.993 15.788 81.025 15.852 ;
			RECT	81.161 15.788 81.193 15.852 ;
			RECT	81.329 15.788 81.361 15.852 ;
			RECT	81.497 15.788 81.529 15.852 ;
			RECT	81.665 15.788 81.697 15.852 ;
			RECT	81.833 15.788 81.865 15.852 ;
			RECT	82.001 15.788 82.033 15.852 ;
			RECT	82.169 15.788 82.201 15.852 ;
			RECT	82.337 15.788 82.369 15.852 ;
			RECT	82.505 15.788 82.537 15.852 ;
			RECT	82.673 15.788 82.705 15.852 ;
			RECT	82.841 15.788 82.873 15.852 ;
			RECT	83.009 15.788 83.041 15.852 ;
			RECT	83.177 15.788 83.209 15.852 ;
			RECT	83.345 15.788 83.377 15.852 ;
			RECT	83.513 15.788 83.545 15.852 ;
			RECT	83.681 15.788 83.713 15.852 ;
			RECT	83.849 15.788 83.881 15.852 ;
			RECT	84.017 15.788 84.049 15.852 ;
			RECT	84.185 15.788 84.217 15.852 ;
			RECT	84.353 15.788 84.385 15.852 ;
			RECT	84.521 15.788 84.553 15.852 ;
			RECT	84.689 15.788 84.721 15.852 ;
			RECT	84.857 15.788 84.889 15.852 ;
			RECT	85.025 15.788 85.057 15.852 ;
			RECT	85.193 15.788 85.225 15.852 ;
			RECT	85.361 15.788 85.393 15.852 ;
			RECT	85.529 15.788 85.561 15.852 ;
			RECT	85.697 15.788 85.729 15.852 ;
			RECT	85.865 15.788 85.897 15.852 ;
			RECT	86.033 15.788 86.065 15.852 ;
			RECT	86.201 15.788 86.233 15.852 ;
			RECT	86.369 15.788 86.401 15.852 ;
			RECT	86.537 15.788 86.569 15.852 ;
			RECT	86.705 15.788 86.737 15.852 ;
			RECT	86.873 15.788 86.905 15.852 ;
			RECT	87.041 15.788 87.073 15.852 ;
			RECT	87.209 15.788 87.241 15.852 ;
			RECT	87.377 15.788 87.409 15.852 ;
			RECT	87.545 15.788 87.577 15.852 ;
			RECT	87.713 15.788 87.745 15.852 ;
			RECT	87.881 15.788 87.913 15.852 ;
			RECT	88.049 15.788 88.081 15.852 ;
			RECT	88.217 15.788 88.249 15.852 ;
			RECT	88.385 15.788 88.417 15.852 ;
			RECT	88.553 15.788 88.585 15.852 ;
			RECT	88.721 15.788 88.753 15.852 ;
			RECT	88.889 15.788 88.921 15.852 ;
			RECT	89.057 15.788 89.089 15.852 ;
			RECT	89.225 15.788 89.257 15.852 ;
			RECT	89.393 15.788 89.425 15.852 ;
			RECT	89.561 15.788 89.593 15.852 ;
			RECT	89.729 15.788 89.761 15.852 ;
			RECT	89.897 15.788 89.929 15.852 ;
			RECT	90.065 15.788 90.097 15.852 ;
			RECT	90.233 15.788 90.265 15.852 ;
			RECT	90.401 15.788 90.433 15.852 ;
			RECT	90.569 15.788 90.601 15.852 ;
			RECT	90.737 15.788 90.769 15.852 ;
			RECT	90.905 15.788 90.937 15.852 ;
			RECT	91.073 15.788 91.105 15.852 ;
			RECT	91.241 15.788 91.273 15.852 ;
			RECT	91.409 15.788 91.441 15.852 ;
			RECT	91.577 15.788 91.609 15.852 ;
			RECT	91.745 15.788 91.777 15.852 ;
			RECT	91.913 15.788 91.945 15.852 ;
			RECT	92.081 15.788 92.113 15.852 ;
			RECT	92.249 15.788 92.281 15.852 ;
			RECT	92.417 15.788 92.449 15.852 ;
			RECT	92.585 15.788 92.617 15.852 ;
			RECT	92.753 15.788 92.785 15.852 ;
			RECT	92.921 15.788 92.953 15.852 ;
			RECT	93.089 15.788 93.121 15.852 ;
			RECT	93.257 15.788 93.289 15.852 ;
			RECT	93.425 15.788 93.457 15.852 ;
			RECT	93.593 15.788 93.625 15.852 ;
			RECT	93.761 15.788 93.793 15.852 ;
			RECT	93.929 15.788 93.961 15.852 ;
			RECT	94.097 15.788 94.129 15.852 ;
			RECT	94.265 15.788 94.297 15.852 ;
			RECT	94.433 15.788 94.465 15.852 ;
			RECT	94.601 15.788 94.633 15.852 ;
			RECT	94.769 15.788 94.801 15.852 ;
			RECT	94.937 15.788 94.969 15.852 ;
			RECT	95.105 15.788 95.137 15.852 ;
			RECT	95.273 15.788 95.305 15.852 ;
			RECT	95.441 15.788 95.473 15.852 ;
			RECT	95.609 15.788 95.641 15.852 ;
			RECT	95.777 15.788 95.809 15.852 ;
			RECT	95.945 15.788 95.977 15.852 ;
			RECT	96.113 15.788 96.145 15.852 ;
			RECT	96.281 15.788 96.313 15.852 ;
			RECT	96.449 15.788 96.481 15.852 ;
			RECT	96.617 15.788 96.649 15.852 ;
			RECT	96.785 15.788 96.817 15.852 ;
			RECT	96.953 15.788 96.985 15.852 ;
			RECT	97.121 15.788 97.153 15.852 ;
			RECT	97.289 15.788 97.321 15.852 ;
			RECT	97.457 15.788 97.489 15.852 ;
			RECT	97.625 15.788 97.657 15.852 ;
			RECT	97.793 15.788 97.825 15.852 ;
			RECT	97.961 15.788 97.993 15.852 ;
			RECT	98.129 15.788 98.161 15.852 ;
			RECT	98.297 15.788 98.329 15.852 ;
			RECT	98.465 15.788 98.497 15.852 ;
			RECT	98.633 15.788 98.665 15.852 ;
			RECT	98.801 15.788 98.833 15.852 ;
			RECT	98.969 15.788 99.001 15.852 ;
			RECT	99.137 15.788 99.169 15.852 ;
			RECT	99.305 15.788 99.337 15.852 ;
			RECT	99.473 15.788 99.505 15.852 ;
			RECT	99.641 15.788 99.673 15.852 ;
			RECT	99.809 15.788 99.841 15.852 ;
			RECT	99.977 15.788 100.009 15.852 ;
			RECT	100.145 15.788 100.177 15.852 ;
			RECT	100.313 15.788 100.345 15.852 ;
			RECT	100.481 15.788 100.513 15.852 ;
			RECT	100.649 15.788 100.681 15.852 ;
			RECT	100.817 15.788 100.849 15.852 ;
			RECT	100.985 15.788 101.017 15.852 ;
			RECT	101.153 15.788 101.185 15.852 ;
			RECT	101.321 15.788 101.353 15.852 ;
			RECT	101.489 15.788 101.521 15.852 ;
			RECT	101.657 15.788 101.689 15.852 ;
			RECT	101.825 15.788 101.857 15.852 ;
			RECT	101.993 15.788 102.025 15.852 ;
			RECT	102.123 15.804 102.155 15.836 ;
			RECT	102.245 15.809 102.277 15.841 ;
			RECT	102.375 15.788 102.407 15.852 ;
			RECT	103.795 15.788 103.827 15.852 ;
			RECT	103.925 15.809 103.957 15.841 ;
			RECT	104.047 15.804 104.079 15.836 ;
			RECT	104.177 15.788 104.209 15.852 ;
			RECT	104.345 15.788 104.377 15.852 ;
			RECT	104.513 15.788 104.545 15.852 ;
			RECT	104.681 15.788 104.713 15.852 ;
			RECT	104.849 15.788 104.881 15.852 ;
			RECT	105.017 15.788 105.049 15.852 ;
			RECT	105.185 15.788 105.217 15.852 ;
			RECT	105.353 15.788 105.385 15.852 ;
			RECT	105.521 15.788 105.553 15.852 ;
			RECT	105.689 15.788 105.721 15.852 ;
			RECT	105.857 15.788 105.889 15.852 ;
			RECT	106.025 15.788 106.057 15.852 ;
			RECT	106.193 15.788 106.225 15.852 ;
			RECT	106.361 15.788 106.393 15.852 ;
			RECT	106.529 15.788 106.561 15.852 ;
			RECT	106.697 15.788 106.729 15.852 ;
			RECT	106.865 15.788 106.897 15.852 ;
			RECT	107.033 15.788 107.065 15.852 ;
			RECT	107.201 15.788 107.233 15.852 ;
			RECT	107.369 15.788 107.401 15.852 ;
			RECT	107.537 15.788 107.569 15.852 ;
			RECT	107.705 15.788 107.737 15.852 ;
			RECT	107.873 15.788 107.905 15.852 ;
			RECT	108.041 15.788 108.073 15.852 ;
			RECT	108.209 15.788 108.241 15.852 ;
			RECT	108.377 15.788 108.409 15.852 ;
			RECT	108.545 15.788 108.577 15.852 ;
			RECT	108.713 15.788 108.745 15.852 ;
			RECT	108.881 15.788 108.913 15.852 ;
			RECT	109.049 15.788 109.081 15.852 ;
			RECT	109.217 15.788 109.249 15.852 ;
			RECT	109.385 15.788 109.417 15.852 ;
			RECT	109.553 15.788 109.585 15.852 ;
			RECT	109.721 15.788 109.753 15.852 ;
			RECT	109.889 15.788 109.921 15.852 ;
			RECT	110.057 15.788 110.089 15.852 ;
			RECT	110.225 15.788 110.257 15.852 ;
			RECT	110.393 15.788 110.425 15.852 ;
			RECT	110.561 15.788 110.593 15.852 ;
			RECT	110.729 15.788 110.761 15.852 ;
			RECT	110.897 15.788 110.929 15.852 ;
			RECT	111.065 15.788 111.097 15.852 ;
			RECT	111.233 15.788 111.265 15.852 ;
			RECT	111.401 15.788 111.433 15.852 ;
			RECT	111.569 15.788 111.601 15.852 ;
			RECT	111.737 15.788 111.769 15.852 ;
			RECT	111.905 15.788 111.937 15.852 ;
			RECT	112.073 15.788 112.105 15.852 ;
			RECT	112.241 15.788 112.273 15.852 ;
			RECT	112.409 15.788 112.441 15.852 ;
			RECT	112.577 15.788 112.609 15.852 ;
			RECT	112.745 15.788 112.777 15.852 ;
			RECT	112.913 15.788 112.945 15.852 ;
			RECT	113.081 15.788 113.113 15.852 ;
			RECT	113.249 15.788 113.281 15.852 ;
			RECT	113.417 15.788 113.449 15.852 ;
			RECT	113.585 15.788 113.617 15.852 ;
			RECT	113.753 15.788 113.785 15.852 ;
			RECT	113.921 15.788 113.953 15.852 ;
			RECT	114.089 15.788 114.121 15.852 ;
			RECT	114.257 15.788 114.289 15.852 ;
			RECT	114.425 15.788 114.457 15.852 ;
			RECT	114.593 15.788 114.625 15.852 ;
			RECT	114.761 15.788 114.793 15.852 ;
			RECT	114.929 15.788 114.961 15.852 ;
			RECT	115.097 15.788 115.129 15.852 ;
			RECT	115.265 15.788 115.297 15.852 ;
			RECT	115.433 15.788 115.465 15.852 ;
			RECT	115.601 15.788 115.633 15.852 ;
			RECT	115.769 15.788 115.801 15.852 ;
			RECT	115.937 15.788 115.969 15.852 ;
			RECT	116.105 15.788 116.137 15.852 ;
			RECT	116.273 15.788 116.305 15.852 ;
			RECT	116.441 15.788 116.473 15.852 ;
			RECT	116.609 15.788 116.641 15.852 ;
			RECT	116.777 15.788 116.809 15.852 ;
			RECT	116.945 15.788 116.977 15.852 ;
			RECT	117.113 15.788 117.145 15.852 ;
			RECT	117.281 15.788 117.313 15.852 ;
			RECT	117.449 15.788 117.481 15.852 ;
			RECT	117.617 15.788 117.649 15.852 ;
			RECT	117.785 15.788 117.817 15.852 ;
			RECT	117.953 15.788 117.985 15.852 ;
			RECT	118.121 15.788 118.153 15.852 ;
			RECT	118.289 15.788 118.321 15.852 ;
			RECT	118.457 15.788 118.489 15.852 ;
			RECT	118.625 15.788 118.657 15.852 ;
			RECT	118.793 15.788 118.825 15.852 ;
			RECT	118.961 15.788 118.993 15.852 ;
			RECT	119.129 15.788 119.161 15.852 ;
			RECT	119.297 15.788 119.329 15.852 ;
			RECT	119.465 15.788 119.497 15.852 ;
			RECT	119.633 15.788 119.665 15.852 ;
			RECT	119.801 15.788 119.833 15.852 ;
			RECT	119.969 15.788 120.001 15.852 ;
			RECT	120.137 15.788 120.169 15.852 ;
			RECT	120.305 15.788 120.337 15.852 ;
			RECT	120.473 15.788 120.505 15.852 ;
			RECT	120.641 15.788 120.673 15.852 ;
			RECT	120.809 15.788 120.841 15.852 ;
			RECT	120.977 15.788 121.009 15.852 ;
			RECT	121.145 15.788 121.177 15.852 ;
			RECT	121.313 15.788 121.345 15.852 ;
			RECT	121.481 15.788 121.513 15.852 ;
			RECT	121.649 15.788 121.681 15.852 ;
			RECT	121.817 15.788 121.849 15.852 ;
			RECT	121.985 15.788 122.017 15.852 ;
			RECT	122.153 15.788 122.185 15.852 ;
			RECT	122.321 15.788 122.353 15.852 ;
			RECT	122.489 15.788 122.521 15.852 ;
			RECT	122.657 15.788 122.689 15.852 ;
			RECT	122.825 15.788 122.857 15.852 ;
			RECT	122.993 15.788 123.025 15.852 ;
			RECT	123.161 15.788 123.193 15.852 ;
			RECT	123.329 15.788 123.361 15.852 ;
			RECT	123.497 15.788 123.529 15.852 ;
			RECT	123.665 15.788 123.697 15.852 ;
			RECT	123.833 15.788 123.865 15.852 ;
			RECT	124.001 15.788 124.033 15.852 ;
			RECT	124.169 15.788 124.201 15.852 ;
			RECT	124.337 15.788 124.369 15.852 ;
			RECT	124.505 15.788 124.537 15.852 ;
			RECT	124.673 15.788 124.705 15.852 ;
			RECT	124.841 15.788 124.873 15.852 ;
			RECT	125.009 15.788 125.041 15.852 ;
			RECT	125.177 15.788 125.209 15.852 ;
			RECT	125.345 15.788 125.377 15.852 ;
			RECT	125.513 15.788 125.545 15.852 ;
			RECT	125.681 15.788 125.713 15.852 ;
			RECT	125.849 15.788 125.881 15.852 ;
			RECT	126.017 15.788 126.049 15.852 ;
			RECT	126.185 15.788 126.217 15.852 ;
			RECT	126.353 15.788 126.385 15.852 ;
			RECT	126.521 15.788 126.553 15.852 ;
			RECT	126.689 15.788 126.721 15.852 ;
			RECT	126.857 15.788 126.889 15.852 ;
			RECT	127.025 15.788 127.057 15.852 ;
			RECT	127.193 15.788 127.225 15.852 ;
			RECT	127.361 15.788 127.393 15.852 ;
			RECT	127.529 15.788 127.561 15.852 ;
			RECT	127.697 15.788 127.729 15.852 ;
			RECT	127.865 15.788 127.897 15.852 ;
			RECT	128.033 15.788 128.065 15.852 ;
			RECT	128.201 15.788 128.233 15.852 ;
			RECT	128.369 15.788 128.401 15.852 ;
			RECT	128.537 15.788 128.569 15.852 ;
			RECT	128.705 15.788 128.737 15.852 ;
			RECT	128.873 15.788 128.905 15.852 ;
			RECT	129.041 15.788 129.073 15.852 ;
			RECT	129.209 15.788 129.241 15.852 ;
			RECT	129.377 15.788 129.409 15.852 ;
			RECT	129.545 15.788 129.577 15.852 ;
			RECT	129.713 15.788 129.745 15.852 ;
			RECT	129.881 15.788 129.913 15.852 ;
			RECT	130.049 15.788 130.081 15.852 ;
			RECT	130.217 15.788 130.249 15.852 ;
			RECT	130.385 15.788 130.417 15.852 ;
			RECT	130.553 15.788 130.585 15.852 ;
			RECT	130.721 15.788 130.753 15.852 ;
			RECT	130.889 15.788 130.921 15.852 ;
			RECT	131.057 15.788 131.089 15.852 ;
			RECT	131.225 15.788 131.257 15.852 ;
			RECT	131.393 15.788 131.425 15.852 ;
			RECT	131.561 15.788 131.593 15.852 ;
			RECT	131.729 15.788 131.761 15.852 ;
			RECT	131.897 15.788 131.929 15.852 ;
			RECT	132.065 15.788 132.097 15.852 ;
			RECT	132.233 15.788 132.265 15.852 ;
			RECT	132.401 15.788 132.433 15.852 ;
			RECT	132.569 15.788 132.601 15.852 ;
			RECT	132.737 15.788 132.769 15.852 ;
			RECT	132.905 15.788 132.937 15.852 ;
			RECT	133.073 15.788 133.105 15.852 ;
			RECT	133.241 15.788 133.273 15.852 ;
			RECT	133.409 15.788 133.441 15.852 ;
			RECT	133.577 15.788 133.609 15.852 ;
			RECT	133.745 15.788 133.777 15.852 ;
			RECT	133.913 15.788 133.945 15.852 ;
			RECT	134.081 15.788 134.113 15.852 ;
			RECT	134.249 15.788 134.281 15.852 ;
			RECT	134.417 15.788 134.449 15.852 ;
			RECT	134.585 15.788 134.617 15.852 ;
			RECT	134.753 15.788 134.785 15.852 ;
			RECT	134.921 15.788 134.953 15.852 ;
			RECT	135.089 15.788 135.121 15.852 ;
			RECT	135.257 15.788 135.289 15.852 ;
			RECT	135.425 15.788 135.457 15.852 ;
			RECT	135.593 15.788 135.625 15.852 ;
			RECT	135.761 15.788 135.793 15.852 ;
			RECT	135.929 15.788 135.961 15.852 ;
			RECT	136.097 15.788 136.129 15.852 ;
			RECT	136.265 15.788 136.297 15.852 ;
			RECT	136.433 15.788 136.465 15.852 ;
			RECT	136.601 15.788 136.633 15.852 ;
			RECT	136.769 15.788 136.801 15.852 ;
			RECT	136.937 15.788 136.969 15.852 ;
			RECT	137.105 15.788 137.137 15.852 ;
			RECT	137.273 15.788 137.305 15.852 ;
			RECT	137.441 15.788 137.473 15.852 ;
			RECT	137.609 15.788 137.641 15.852 ;
			RECT	137.777 15.788 137.809 15.852 ;
			RECT	137.945 15.788 137.977 15.852 ;
			RECT	138.113 15.788 138.145 15.852 ;
			RECT	138.281 15.788 138.313 15.852 ;
			RECT	138.449 15.788 138.481 15.852 ;
			RECT	138.617 15.788 138.649 15.852 ;
			RECT	138.785 15.788 138.817 15.852 ;
			RECT	138.953 15.788 138.985 15.852 ;
			RECT	139.121 15.788 139.153 15.852 ;
			RECT	139.289 15.788 139.321 15.852 ;
			RECT	139.457 15.788 139.489 15.852 ;
			RECT	139.625 15.788 139.657 15.852 ;
			RECT	139.793 15.788 139.825 15.852 ;
			RECT	139.961 15.788 139.993 15.852 ;
			RECT	140.129 15.788 140.161 15.852 ;
			RECT	140.297 15.788 140.329 15.852 ;
			RECT	140.465 15.788 140.497 15.852 ;
			RECT	140.633 15.788 140.665 15.852 ;
			RECT	140.801 15.788 140.833 15.852 ;
			RECT	140.969 15.788 141.001 15.852 ;
			RECT	141.137 15.788 141.169 15.852 ;
			RECT	141.305 15.788 141.337 15.852 ;
			RECT	141.473 15.788 141.505 15.852 ;
			RECT	141.641 15.788 141.673 15.852 ;
			RECT	141.809 15.788 141.841 15.852 ;
			RECT	141.977 15.788 142.009 15.852 ;
			RECT	142.145 15.788 142.177 15.852 ;
			RECT	142.313 15.788 142.345 15.852 ;
			RECT	142.481 15.788 142.513 15.852 ;
			RECT	142.649 15.788 142.681 15.852 ;
			RECT	142.817 15.788 142.849 15.852 ;
			RECT	142.985 15.788 143.017 15.852 ;
			RECT	143.153 15.788 143.185 15.852 ;
			RECT	143.321 15.788 143.353 15.852 ;
			RECT	143.489 15.788 143.521 15.852 ;
			RECT	143.657 15.788 143.689 15.852 ;
			RECT	143.825 15.788 143.857 15.852 ;
			RECT	143.993 15.788 144.025 15.852 ;
			RECT	144.161 15.788 144.193 15.852 ;
			RECT	144.329 15.788 144.361 15.852 ;
			RECT	144.497 15.788 144.529 15.852 ;
			RECT	144.665 15.788 144.697 15.852 ;
			RECT	144.833 15.788 144.865 15.852 ;
			RECT	145.001 15.788 145.033 15.852 ;
			RECT	145.169 15.788 145.201 15.852 ;
			RECT	145.337 15.788 145.369 15.852 ;
			RECT	145.505 15.788 145.537 15.852 ;
			RECT	145.673 15.788 145.705 15.852 ;
			RECT	145.841 15.788 145.873 15.852 ;
			RECT	146.009 15.788 146.041 15.852 ;
			RECT	146.177 15.788 146.209 15.852 ;
			RECT	146.345 15.788 146.377 15.852 ;
			RECT	146.513 15.788 146.545 15.852 ;
			RECT	146.681 15.788 146.713 15.852 ;
			RECT	146.849 15.788 146.881 15.852 ;
			RECT	147.017 15.788 147.049 15.852 ;
			RECT	147.185 15.788 147.217 15.852 ;
			RECT	147.316 15.804 147.348 15.836 ;
			RECT	147.437 15.804 147.469 15.836 ;
			RECT	147.567 15.788 147.599 15.852 ;
			RECT	149.879 15.788 149.911 15.852 ;
			RECT	151.13 15.788 151.194 15.852 ;
			RECT	151.81 15.788 151.842 15.852 ;
			RECT	152.249 15.788 152.281 15.852 ;
			RECT	153.56 15.788 153.624 15.852 ;
			RECT	156.601 15.788 156.633 15.852 ;
			RECT	156.731 15.804 156.763 15.836 ;
			RECT	156.852 15.804 156.884 15.836 ;
			RECT	156.983 15.788 157.015 15.852 ;
			RECT	157.151 15.788 157.183 15.852 ;
			RECT	157.319 15.788 157.351 15.852 ;
			RECT	157.487 15.788 157.519 15.852 ;
			RECT	157.655 15.788 157.687 15.852 ;
			RECT	157.823 15.788 157.855 15.852 ;
			RECT	157.991 15.788 158.023 15.852 ;
			RECT	158.159 15.788 158.191 15.852 ;
			RECT	158.327 15.788 158.359 15.852 ;
			RECT	158.495 15.788 158.527 15.852 ;
			RECT	158.663 15.788 158.695 15.852 ;
			RECT	158.831 15.788 158.863 15.852 ;
			RECT	158.999 15.788 159.031 15.852 ;
			RECT	159.167 15.788 159.199 15.852 ;
			RECT	159.335 15.788 159.367 15.852 ;
			RECT	159.503 15.788 159.535 15.852 ;
			RECT	159.671 15.788 159.703 15.852 ;
			RECT	159.839 15.788 159.871 15.852 ;
			RECT	160.007 15.788 160.039 15.852 ;
			RECT	160.175 15.788 160.207 15.852 ;
			RECT	160.343 15.788 160.375 15.852 ;
			RECT	160.511 15.788 160.543 15.852 ;
			RECT	160.679 15.788 160.711 15.852 ;
			RECT	160.847 15.788 160.879 15.852 ;
			RECT	161.015 15.788 161.047 15.852 ;
			RECT	161.183 15.788 161.215 15.852 ;
			RECT	161.351 15.788 161.383 15.852 ;
			RECT	161.519 15.788 161.551 15.852 ;
			RECT	161.687 15.788 161.719 15.852 ;
			RECT	161.855 15.788 161.887 15.852 ;
			RECT	162.023 15.788 162.055 15.852 ;
			RECT	162.191 15.788 162.223 15.852 ;
			RECT	162.359 15.788 162.391 15.852 ;
			RECT	162.527 15.788 162.559 15.852 ;
			RECT	162.695 15.788 162.727 15.852 ;
			RECT	162.863 15.788 162.895 15.852 ;
			RECT	163.031 15.788 163.063 15.852 ;
			RECT	163.199 15.788 163.231 15.852 ;
			RECT	163.367 15.788 163.399 15.852 ;
			RECT	163.535 15.788 163.567 15.852 ;
			RECT	163.703 15.788 163.735 15.852 ;
			RECT	163.871 15.788 163.903 15.852 ;
			RECT	164.039 15.788 164.071 15.852 ;
			RECT	164.207 15.788 164.239 15.852 ;
			RECT	164.375 15.788 164.407 15.852 ;
			RECT	164.543 15.788 164.575 15.852 ;
			RECT	164.711 15.788 164.743 15.852 ;
			RECT	164.879 15.788 164.911 15.852 ;
			RECT	165.047 15.788 165.079 15.852 ;
			RECT	165.215 15.788 165.247 15.852 ;
			RECT	165.383 15.788 165.415 15.852 ;
			RECT	165.551 15.788 165.583 15.852 ;
			RECT	165.719 15.788 165.751 15.852 ;
			RECT	165.887 15.788 165.919 15.852 ;
			RECT	166.055 15.788 166.087 15.852 ;
			RECT	166.223 15.788 166.255 15.852 ;
			RECT	166.391 15.788 166.423 15.852 ;
			RECT	166.559 15.788 166.591 15.852 ;
			RECT	166.727 15.788 166.759 15.852 ;
			RECT	166.895 15.788 166.927 15.852 ;
			RECT	167.063 15.788 167.095 15.852 ;
			RECT	167.231 15.788 167.263 15.852 ;
			RECT	167.399 15.788 167.431 15.852 ;
			RECT	167.567 15.788 167.599 15.852 ;
			RECT	167.735 15.788 167.767 15.852 ;
			RECT	167.903 15.788 167.935 15.852 ;
			RECT	168.071 15.788 168.103 15.852 ;
			RECT	168.239 15.788 168.271 15.852 ;
			RECT	168.407 15.788 168.439 15.852 ;
			RECT	168.575 15.788 168.607 15.852 ;
			RECT	168.743 15.788 168.775 15.852 ;
			RECT	168.911 15.788 168.943 15.852 ;
			RECT	169.079 15.788 169.111 15.852 ;
			RECT	169.247 15.788 169.279 15.852 ;
			RECT	169.415 15.788 169.447 15.852 ;
			RECT	169.583 15.788 169.615 15.852 ;
			RECT	169.751 15.788 169.783 15.852 ;
			RECT	169.919 15.788 169.951 15.852 ;
			RECT	170.087 15.788 170.119 15.852 ;
			RECT	170.255 15.788 170.287 15.852 ;
			RECT	170.423 15.788 170.455 15.852 ;
			RECT	170.591 15.788 170.623 15.852 ;
			RECT	170.759 15.788 170.791 15.852 ;
			RECT	170.927 15.788 170.959 15.852 ;
			RECT	171.095 15.788 171.127 15.852 ;
			RECT	171.263 15.788 171.295 15.852 ;
			RECT	171.431 15.788 171.463 15.852 ;
			RECT	171.599 15.788 171.631 15.852 ;
			RECT	171.767 15.788 171.799 15.852 ;
			RECT	171.935 15.788 171.967 15.852 ;
			RECT	172.103 15.788 172.135 15.852 ;
			RECT	172.271 15.788 172.303 15.852 ;
			RECT	172.439 15.788 172.471 15.852 ;
			RECT	172.607 15.788 172.639 15.852 ;
			RECT	172.775 15.788 172.807 15.852 ;
			RECT	172.943 15.788 172.975 15.852 ;
			RECT	173.111 15.788 173.143 15.852 ;
			RECT	173.279 15.788 173.311 15.852 ;
			RECT	173.447 15.788 173.479 15.852 ;
			RECT	173.615 15.788 173.647 15.852 ;
			RECT	173.783 15.788 173.815 15.852 ;
			RECT	173.951 15.788 173.983 15.852 ;
			RECT	174.119 15.788 174.151 15.852 ;
			RECT	174.287 15.788 174.319 15.852 ;
			RECT	174.455 15.788 174.487 15.852 ;
			RECT	174.623 15.788 174.655 15.852 ;
			RECT	174.791 15.788 174.823 15.852 ;
			RECT	174.959 15.788 174.991 15.852 ;
			RECT	175.127 15.788 175.159 15.852 ;
			RECT	175.295 15.788 175.327 15.852 ;
			RECT	175.463 15.788 175.495 15.852 ;
			RECT	175.631 15.788 175.663 15.852 ;
			RECT	175.799 15.788 175.831 15.852 ;
			RECT	175.967 15.788 175.999 15.852 ;
			RECT	176.135 15.788 176.167 15.852 ;
			RECT	176.303 15.788 176.335 15.852 ;
			RECT	176.471 15.788 176.503 15.852 ;
			RECT	176.639 15.788 176.671 15.852 ;
			RECT	176.807 15.788 176.839 15.852 ;
			RECT	176.975 15.788 177.007 15.852 ;
			RECT	177.143 15.788 177.175 15.852 ;
			RECT	177.311 15.788 177.343 15.852 ;
			RECT	177.479 15.788 177.511 15.852 ;
			RECT	177.647 15.788 177.679 15.852 ;
			RECT	177.815 15.788 177.847 15.852 ;
			RECT	177.983 15.788 178.015 15.852 ;
			RECT	178.151 15.788 178.183 15.852 ;
			RECT	178.319 15.788 178.351 15.852 ;
			RECT	178.487 15.788 178.519 15.852 ;
			RECT	178.655 15.788 178.687 15.852 ;
			RECT	178.823 15.788 178.855 15.852 ;
			RECT	178.991 15.788 179.023 15.852 ;
			RECT	179.159 15.788 179.191 15.852 ;
			RECT	179.327 15.788 179.359 15.852 ;
			RECT	179.495 15.788 179.527 15.852 ;
			RECT	179.663 15.788 179.695 15.852 ;
			RECT	179.831 15.788 179.863 15.852 ;
			RECT	179.999 15.788 180.031 15.852 ;
			RECT	180.167 15.788 180.199 15.852 ;
			RECT	180.335 15.788 180.367 15.852 ;
			RECT	180.503 15.788 180.535 15.852 ;
			RECT	180.671 15.788 180.703 15.852 ;
			RECT	180.839 15.788 180.871 15.852 ;
			RECT	181.007 15.788 181.039 15.852 ;
			RECT	181.175 15.788 181.207 15.852 ;
			RECT	181.343 15.788 181.375 15.852 ;
			RECT	181.511 15.788 181.543 15.852 ;
			RECT	181.679 15.788 181.711 15.852 ;
			RECT	181.847 15.788 181.879 15.852 ;
			RECT	182.015 15.788 182.047 15.852 ;
			RECT	182.183 15.788 182.215 15.852 ;
			RECT	182.351 15.788 182.383 15.852 ;
			RECT	182.519 15.788 182.551 15.852 ;
			RECT	182.687 15.788 182.719 15.852 ;
			RECT	182.855 15.788 182.887 15.852 ;
			RECT	183.023 15.788 183.055 15.852 ;
			RECT	183.191 15.788 183.223 15.852 ;
			RECT	183.359 15.788 183.391 15.852 ;
			RECT	183.527 15.788 183.559 15.852 ;
			RECT	183.695 15.788 183.727 15.852 ;
			RECT	183.863 15.788 183.895 15.852 ;
			RECT	184.031 15.788 184.063 15.852 ;
			RECT	184.199 15.788 184.231 15.852 ;
			RECT	184.367 15.788 184.399 15.852 ;
			RECT	184.535 15.788 184.567 15.852 ;
			RECT	184.703 15.788 184.735 15.852 ;
			RECT	184.871 15.788 184.903 15.852 ;
			RECT	185.039 15.788 185.071 15.852 ;
			RECT	185.207 15.788 185.239 15.852 ;
			RECT	185.375 15.788 185.407 15.852 ;
			RECT	185.543 15.788 185.575 15.852 ;
			RECT	185.711 15.788 185.743 15.852 ;
			RECT	185.879 15.788 185.911 15.852 ;
			RECT	186.047 15.788 186.079 15.852 ;
			RECT	186.215 15.788 186.247 15.852 ;
			RECT	186.383 15.788 186.415 15.852 ;
			RECT	186.551 15.788 186.583 15.852 ;
			RECT	186.719 15.788 186.751 15.852 ;
			RECT	186.887 15.788 186.919 15.852 ;
			RECT	187.055 15.788 187.087 15.852 ;
			RECT	187.223 15.788 187.255 15.852 ;
			RECT	187.391 15.788 187.423 15.852 ;
			RECT	187.559 15.788 187.591 15.852 ;
			RECT	187.727 15.788 187.759 15.852 ;
			RECT	187.895 15.788 187.927 15.852 ;
			RECT	188.063 15.788 188.095 15.852 ;
			RECT	188.231 15.788 188.263 15.852 ;
			RECT	188.399 15.788 188.431 15.852 ;
			RECT	188.567 15.788 188.599 15.852 ;
			RECT	188.735 15.788 188.767 15.852 ;
			RECT	188.903 15.788 188.935 15.852 ;
			RECT	189.071 15.788 189.103 15.852 ;
			RECT	189.239 15.788 189.271 15.852 ;
			RECT	189.407 15.788 189.439 15.852 ;
			RECT	189.575 15.788 189.607 15.852 ;
			RECT	189.743 15.788 189.775 15.852 ;
			RECT	189.911 15.788 189.943 15.852 ;
			RECT	190.079 15.788 190.111 15.852 ;
			RECT	190.247 15.788 190.279 15.852 ;
			RECT	190.415 15.788 190.447 15.852 ;
			RECT	190.583 15.788 190.615 15.852 ;
			RECT	190.751 15.788 190.783 15.852 ;
			RECT	190.919 15.788 190.951 15.852 ;
			RECT	191.087 15.788 191.119 15.852 ;
			RECT	191.255 15.788 191.287 15.852 ;
			RECT	191.423 15.788 191.455 15.852 ;
			RECT	191.591 15.788 191.623 15.852 ;
			RECT	191.759 15.788 191.791 15.852 ;
			RECT	191.927 15.788 191.959 15.852 ;
			RECT	192.095 15.788 192.127 15.852 ;
			RECT	192.263 15.788 192.295 15.852 ;
			RECT	192.431 15.788 192.463 15.852 ;
			RECT	192.599 15.788 192.631 15.852 ;
			RECT	192.767 15.788 192.799 15.852 ;
			RECT	192.935 15.788 192.967 15.852 ;
			RECT	193.103 15.788 193.135 15.852 ;
			RECT	193.271 15.788 193.303 15.852 ;
			RECT	193.439 15.788 193.471 15.852 ;
			RECT	193.607 15.788 193.639 15.852 ;
			RECT	193.775 15.788 193.807 15.852 ;
			RECT	193.943 15.788 193.975 15.852 ;
			RECT	194.111 15.788 194.143 15.852 ;
			RECT	194.279 15.788 194.311 15.852 ;
			RECT	194.447 15.788 194.479 15.852 ;
			RECT	194.615 15.788 194.647 15.852 ;
			RECT	194.783 15.788 194.815 15.852 ;
			RECT	194.951 15.788 194.983 15.852 ;
			RECT	195.119 15.788 195.151 15.852 ;
			RECT	195.287 15.788 195.319 15.852 ;
			RECT	195.455 15.788 195.487 15.852 ;
			RECT	195.623 15.788 195.655 15.852 ;
			RECT	195.791 15.788 195.823 15.852 ;
			RECT	195.959 15.788 195.991 15.852 ;
			RECT	196.127 15.788 196.159 15.852 ;
			RECT	196.295 15.788 196.327 15.852 ;
			RECT	196.463 15.788 196.495 15.852 ;
			RECT	196.631 15.788 196.663 15.852 ;
			RECT	196.799 15.788 196.831 15.852 ;
			RECT	196.967 15.788 196.999 15.852 ;
			RECT	197.135 15.788 197.167 15.852 ;
			RECT	197.303 15.788 197.335 15.852 ;
			RECT	197.471 15.788 197.503 15.852 ;
			RECT	197.639 15.788 197.671 15.852 ;
			RECT	197.807 15.788 197.839 15.852 ;
			RECT	197.975 15.788 198.007 15.852 ;
			RECT	198.143 15.788 198.175 15.852 ;
			RECT	198.311 15.788 198.343 15.852 ;
			RECT	198.479 15.788 198.511 15.852 ;
			RECT	198.647 15.788 198.679 15.852 ;
			RECT	198.815 15.788 198.847 15.852 ;
			RECT	198.983 15.788 199.015 15.852 ;
			RECT	199.151 15.788 199.183 15.852 ;
			RECT	199.319 15.788 199.351 15.852 ;
			RECT	199.487 15.788 199.519 15.852 ;
			RECT	199.655 15.788 199.687 15.852 ;
			RECT	199.823 15.788 199.855 15.852 ;
			RECT	199.991 15.788 200.023 15.852 ;
			RECT	200.121 15.804 200.153 15.836 ;
			RECT	200.243 15.809 200.275 15.841 ;
			RECT	200.373 15.788 200.405 15.852 ;
			RECT	200.9 15.788 200.932 15.852 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 13.84 201.665 13.96 ;
			LAYER	J3 ;
			RECT	0.755 13.868 0.787 13.932 ;
			RECT	1.645 13.868 1.709 13.932 ;
			RECT	2.323 13.868 2.387 13.932 ;
			RECT	3.438 13.868 3.47 13.932 ;
			RECT	3.585 13.868 3.617 13.932 ;
			RECT	4.195 13.868 4.227 13.932 ;
			RECT	4.72 13.868 4.752 13.932 ;
			RECT	4.944 13.868 5.008 13.932 ;
			RECT	5.267 13.868 5.299 13.932 ;
			RECT	5.797 13.868 5.829 13.932 ;
			RECT	5.927 13.889 5.959 13.921 ;
			RECT	6.049 13.884 6.081 13.916 ;
			RECT	6.179 13.868 6.211 13.932 ;
			RECT	6.347 13.868 6.379 13.932 ;
			RECT	6.515 13.868 6.547 13.932 ;
			RECT	6.683 13.868 6.715 13.932 ;
			RECT	6.851 13.868 6.883 13.932 ;
			RECT	7.019 13.868 7.051 13.932 ;
			RECT	7.187 13.868 7.219 13.932 ;
			RECT	7.355 13.868 7.387 13.932 ;
			RECT	7.523 13.868 7.555 13.932 ;
			RECT	7.691 13.868 7.723 13.932 ;
			RECT	7.859 13.868 7.891 13.932 ;
			RECT	8.027 13.868 8.059 13.932 ;
			RECT	8.195 13.868 8.227 13.932 ;
			RECT	8.363 13.868 8.395 13.932 ;
			RECT	8.531 13.868 8.563 13.932 ;
			RECT	8.699 13.868 8.731 13.932 ;
			RECT	8.867 13.868 8.899 13.932 ;
			RECT	9.035 13.868 9.067 13.932 ;
			RECT	9.203 13.868 9.235 13.932 ;
			RECT	9.371 13.868 9.403 13.932 ;
			RECT	9.539 13.868 9.571 13.932 ;
			RECT	9.707 13.868 9.739 13.932 ;
			RECT	9.875 13.868 9.907 13.932 ;
			RECT	10.043 13.868 10.075 13.932 ;
			RECT	10.211 13.868 10.243 13.932 ;
			RECT	10.379 13.868 10.411 13.932 ;
			RECT	10.547 13.868 10.579 13.932 ;
			RECT	10.715 13.868 10.747 13.932 ;
			RECT	10.883 13.868 10.915 13.932 ;
			RECT	11.051 13.868 11.083 13.932 ;
			RECT	11.219 13.868 11.251 13.932 ;
			RECT	11.387 13.868 11.419 13.932 ;
			RECT	11.555 13.868 11.587 13.932 ;
			RECT	11.723 13.868 11.755 13.932 ;
			RECT	11.891 13.868 11.923 13.932 ;
			RECT	12.059 13.868 12.091 13.932 ;
			RECT	12.227 13.868 12.259 13.932 ;
			RECT	12.395 13.868 12.427 13.932 ;
			RECT	12.563 13.868 12.595 13.932 ;
			RECT	12.731 13.868 12.763 13.932 ;
			RECT	12.899 13.868 12.931 13.932 ;
			RECT	13.067 13.868 13.099 13.932 ;
			RECT	13.235 13.868 13.267 13.932 ;
			RECT	13.403 13.868 13.435 13.932 ;
			RECT	13.571 13.868 13.603 13.932 ;
			RECT	13.739 13.868 13.771 13.932 ;
			RECT	13.907 13.868 13.939 13.932 ;
			RECT	14.075 13.868 14.107 13.932 ;
			RECT	14.243 13.868 14.275 13.932 ;
			RECT	14.411 13.868 14.443 13.932 ;
			RECT	14.579 13.868 14.611 13.932 ;
			RECT	14.747 13.868 14.779 13.932 ;
			RECT	14.915 13.868 14.947 13.932 ;
			RECT	15.083 13.868 15.115 13.932 ;
			RECT	15.251 13.868 15.283 13.932 ;
			RECT	15.419 13.868 15.451 13.932 ;
			RECT	15.587 13.868 15.619 13.932 ;
			RECT	15.755 13.868 15.787 13.932 ;
			RECT	15.923 13.868 15.955 13.932 ;
			RECT	16.091 13.868 16.123 13.932 ;
			RECT	16.259 13.868 16.291 13.932 ;
			RECT	16.427 13.868 16.459 13.932 ;
			RECT	16.595 13.868 16.627 13.932 ;
			RECT	16.763 13.868 16.795 13.932 ;
			RECT	16.931 13.868 16.963 13.932 ;
			RECT	17.099 13.868 17.131 13.932 ;
			RECT	17.267 13.868 17.299 13.932 ;
			RECT	17.435 13.868 17.467 13.932 ;
			RECT	17.603 13.868 17.635 13.932 ;
			RECT	17.771 13.868 17.803 13.932 ;
			RECT	17.939 13.868 17.971 13.932 ;
			RECT	18.107 13.868 18.139 13.932 ;
			RECT	18.275 13.868 18.307 13.932 ;
			RECT	18.443 13.868 18.475 13.932 ;
			RECT	18.611 13.868 18.643 13.932 ;
			RECT	18.779 13.868 18.811 13.932 ;
			RECT	18.947 13.868 18.979 13.932 ;
			RECT	19.115 13.868 19.147 13.932 ;
			RECT	19.283 13.868 19.315 13.932 ;
			RECT	19.451 13.868 19.483 13.932 ;
			RECT	19.619 13.868 19.651 13.932 ;
			RECT	19.787 13.868 19.819 13.932 ;
			RECT	19.955 13.868 19.987 13.932 ;
			RECT	20.123 13.868 20.155 13.932 ;
			RECT	20.291 13.868 20.323 13.932 ;
			RECT	20.459 13.868 20.491 13.932 ;
			RECT	20.627 13.868 20.659 13.932 ;
			RECT	20.795 13.868 20.827 13.932 ;
			RECT	20.963 13.868 20.995 13.932 ;
			RECT	21.131 13.868 21.163 13.932 ;
			RECT	21.299 13.868 21.331 13.932 ;
			RECT	21.467 13.868 21.499 13.932 ;
			RECT	21.635 13.868 21.667 13.932 ;
			RECT	21.803 13.868 21.835 13.932 ;
			RECT	21.971 13.868 22.003 13.932 ;
			RECT	22.139 13.868 22.171 13.932 ;
			RECT	22.307 13.868 22.339 13.932 ;
			RECT	22.475 13.868 22.507 13.932 ;
			RECT	22.643 13.868 22.675 13.932 ;
			RECT	22.811 13.868 22.843 13.932 ;
			RECT	22.979 13.868 23.011 13.932 ;
			RECT	23.147 13.868 23.179 13.932 ;
			RECT	23.315 13.868 23.347 13.932 ;
			RECT	23.483 13.868 23.515 13.932 ;
			RECT	23.651 13.868 23.683 13.932 ;
			RECT	23.819 13.868 23.851 13.932 ;
			RECT	23.987 13.868 24.019 13.932 ;
			RECT	24.155 13.868 24.187 13.932 ;
			RECT	24.323 13.868 24.355 13.932 ;
			RECT	24.491 13.868 24.523 13.932 ;
			RECT	24.659 13.868 24.691 13.932 ;
			RECT	24.827 13.868 24.859 13.932 ;
			RECT	24.995 13.868 25.027 13.932 ;
			RECT	25.163 13.868 25.195 13.932 ;
			RECT	25.331 13.868 25.363 13.932 ;
			RECT	25.499 13.868 25.531 13.932 ;
			RECT	25.667 13.868 25.699 13.932 ;
			RECT	25.835 13.868 25.867 13.932 ;
			RECT	26.003 13.868 26.035 13.932 ;
			RECT	26.171 13.868 26.203 13.932 ;
			RECT	26.339 13.868 26.371 13.932 ;
			RECT	26.507 13.868 26.539 13.932 ;
			RECT	26.675 13.868 26.707 13.932 ;
			RECT	26.843 13.868 26.875 13.932 ;
			RECT	27.011 13.868 27.043 13.932 ;
			RECT	27.179 13.868 27.211 13.932 ;
			RECT	27.347 13.868 27.379 13.932 ;
			RECT	27.515 13.868 27.547 13.932 ;
			RECT	27.683 13.868 27.715 13.932 ;
			RECT	27.851 13.868 27.883 13.932 ;
			RECT	28.019 13.868 28.051 13.932 ;
			RECT	28.187 13.868 28.219 13.932 ;
			RECT	28.355 13.868 28.387 13.932 ;
			RECT	28.523 13.868 28.555 13.932 ;
			RECT	28.691 13.868 28.723 13.932 ;
			RECT	28.859 13.868 28.891 13.932 ;
			RECT	29.027 13.868 29.059 13.932 ;
			RECT	29.195 13.868 29.227 13.932 ;
			RECT	29.363 13.868 29.395 13.932 ;
			RECT	29.531 13.868 29.563 13.932 ;
			RECT	29.699 13.868 29.731 13.932 ;
			RECT	29.867 13.868 29.899 13.932 ;
			RECT	30.035 13.868 30.067 13.932 ;
			RECT	30.203 13.868 30.235 13.932 ;
			RECT	30.371 13.868 30.403 13.932 ;
			RECT	30.539 13.868 30.571 13.932 ;
			RECT	30.707 13.868 30.739 13.932 ;
			RECT	30.875 13.868 30.907 13.932 ;
			RECT	31.043 13.868 31.075 13.932 ;
			RECT	31.211 13.868 31.243 13.932 ;
			RECT	31.379 13.868 31.411 13.932 ;
			RECT	31.547 13.868 31.579 13.932 ;
			RECT	31.715 13.868 31.747 13.932 ;
			RECT	31.883 13.868 31.915 13.932 ;
			RECT	32.051 13.868 32.083 13.932 ;
			RECT	32.219 13.868 32.251 13.932 ;
			RECT	32.387 13.868 32.419 13.932 ;
			RECT	32.555 13.868 32.587 13.932 ;
			RECT	32.723 13.868 32.755 13.932 ;
			RECT	32.891 13.868 32.923 13.932 ;
			RECT	33.059 13.868 33.091 13.932 ;
			RECT	33.227 13.868 33.259 13.932 ;
			RECT	33.395 13.868 33.427 13.932 ;
			RECT	33.563 13.868 33.595 13.932 ;
			RECT	33.731 13.868 33.763 13.932 ;
			RECT	33.899 13.868 33.931 13.932 ;
			RECT	34.067 13.868 34.099 13.932 ;
			RECT	34.235 13.868 34.267 13.932 ;
			RECT	34.403 13.868 34.435 13.932 ;
			RECT	34.571 13.868 34.603 13.932 ;
			RECT	34.739 13.868 34.771 13.932 ;
			RECT	34.907 13.868 34.939 13.932 ;
			RECT	35.075 13.868 35.107 13.932 ;
			RECT	35.243 13.868 35.275 13.932 ;
			RECT	35.411 13.868 35.443 13.932 ;
			RECT	35.579 13.868 35.611 13.932 ;
			RECT	35.747 13.868 35.779 13.932 ;
			RECT	35.915 13.868 35.947 13.932 ;
			RECT	36.083 13.868 36.115 13.932 ;
			RECT	36.251 13.868 36.283 13.932 ;
			RECT	36.419 13.868 36.451 13.932 ;
			RECT	36.587 13.868 36.619 13.932 ;
			RECT	36.755 13.868 36.787 13.932 ;
			RECT	36.923 13.868 36.955 13.932 ;
			RECT	37.091 13.868 37.123 13.932 ;
			RECT	37.259 13.868 37.291 13.932 ;
			RECT	37.427 13.868 37.459 13.932 ;
			RECT	37.595 13.868 37.627 13.932 ;
			RECT	37.763 13.868 37.795 13.932 ;
			RECT	37.931 13.868 37.963 13.932 ;
			RECT	38.099 13.868 38.131 13.932 ;
			RECT	38.267 13.868 38.299 13.932 ;
			RECT	38.435 13.868 38.467 13.932 ;
			RECT	38.603 13.868 38.635 13.932 ;
			RECT	38.771 13.868 38.803 13.932 ;
			RECT	38.939 13.868 38.971 13.932 ;
			RECT	39.107 13.868 39.139 13.932 ;
			RECT	39.275 13.868 39.307 13.932 ;
			RECT	39.443 13.868 39.475 13.932 ;
			RECT	39.611 13.868 39.643 13.932 ;
			RECT	39.779 13.868 39.811 13.932 ;
			RECT	39.947 13.868 39.979 13.932 ;
			RECT	40.115 13.868 40.147 13.932 ;
			RECT	40.283 13.868 40.315 13.932 ;
			RECT	40.451 13.868 40.483 13.932 ;
			RECT	40.619 13.868 40.651 13.932 ;
			RECT	40.787 13.868 40.819 13.932 ;
			RECT	40.955 13.868 40.987 13.932 ;
			RECT	41.123 13.868 41.155 13.932 ;
			RECT	41.291 13.868 41.323 13.932 ;
			RECT	41.459 13.868 41.491 13.932 ;
			RECT	41.627 13.868 41.659 13.932 ;
			RECT	41.795 13.868 41.827 13.932 ;
			RECT	41.963 13.868 41.995 13.932 ;
			RECT	42.131 13.868 42.163 13.932 ;
			RECT	42.299 13.868 42.331 13.932 ;
			RECT	42.467 13.868 42.499 13.932 ;
			RECT	42.635 13.868 42.667 13.932 ;
			RECT	42.803 13.868 42.835 13.932 ;
			RECT	42.971 13.868 43.003 13.932 ;
			RECT	43.139 13.868 43.171 13.932 ;
			RECT	43.307 13.868 43.339 13.932 ;
			RECT	43.475 13.868 43.507 13.932 ;
			RECT	43.643 13.868 43.675 13.932 ;
			RECT	43.811 13.868 43.843 13.932 ;
			RECT	43.979 13.868 44.011 13.932 ;
			RECT	44.147 13.868 44.179 13.932 ;
			RECT	44.315 13.868 44.347 13.932 ;
			RECT	44.483 13.868 44.515 13.932 ;
			RECT	44.651 13.868 44.683 13.932 ;
			RECT	44.819 13.868 44.851 13.932 ;
			RECT	44.987 13.868 45.019 13.932 ;
			RECT	45.155 13.868 45.187 13.932 ;
			RECT	45.323 13.868 45.355 13.932 ;
			RECT	45.491 13.868 45.523 13.932 ;
			RECT	45.659 13.868 45.691 13.932 ;
			RECT	45.827 13.868 45.859 13.932 ;
			RECT	45.995 13.868 46.027 13.932 ;
			RECT	46.163 13.868 46.195 13.932 ;
			RECT	46.331 13.868 46.363 13.932 ;
			RECT	46.499 13.868 46.531 13.932 ;
			RECT	46.667 13.868 46.699 13.932 ;
			RECT	46.835 13.868 46.867 13.932 ;
			RECT	47.003 13.868 47.035 13.932 ;
			RECT	47.171 13.868 47.203 13.932 ;
			RECT	47.339 13.868 47.371 13.932 ;
			RECT	47.507 13.868 47.539 13.932 ;
			RECT	47.675 13.868 47.707 13.932 ;
			RECT	47.843 13.868 47.875 13.932 ;
			RECT	48.011 13.868 48.043 13.932 ;
			RECT	48.179 13.868 48.211 13.932 ;
			RECT	48.347 13.868 48.379 13.932 ;
			RECT	48.515 13.868 48.547 13.932 ;
			RECT	48.683 13.868 48.715 13.932 ;
			RECT	48.851 13.868 48.883 13.932 ;
			RECT	49.019 13.868 49.051 13.932 ;
			RECT	49.187 13.868 49.219 13.932 ;
			RECT	49.318 13.884 49.35 13.916 ;
			RECT	49.439 13.884 49.471 13.916 ;
			RECT	49.569 13.868 49.601 13.932 ;
			RECT	51.881 13.868 51.913 13.932 ;
			RECT	53.132 13.868 53.196 13.932 ;
			RECT	53.812 13.868 53.844 13.932 ;
			RECT	54.251 13.868 54.283 13.932 ;
			RECT	55.562 13.868 55.626 13.932 ;
			RECT	58.603 13.868 58.635 13.932 ;
			RECT	58.733 13.884 58.765 13.916 ;
			RECT	58.854 13.884 58.886 13.916 ;
			RECT	58.985 13.868 59.017 13.932 ;
			RECT	59.153 13.868 59.185 13.932 ;
			RECT	59.321 13.868 59.353 13.932 ;
			RECT	59.489 13.868 59.521 13.932 ;
			RECT	59.657 13.868 59.689 13.932 ;
			RECT	59.825 13.868 59.857 13.932 ;
			RECT	59.993 13.868 60.025 13.932 ;
			RECT	60.161 13.868 60.193 13.932 ;
			RECT	60.329 13.868 60.361 13.932 ;
			RECT	60.497 13.868 60.529 13.932 ;
			RECT	60.665 13.868 60.697 13.932 ;
			RECT	60.833 13.868 60.865 13.932 ;
			RECT	61.001 13.868 61.033 13.932 ;
			RECT	61.169 13.868 61.201 13.932 ;
			RECT	61.337 13.868 61.369 13.932 ;
			RECT	61.505 13.868 61.537 13.932 ;
			RECT	61.673 13.868 61.705 13.932 ;
			RECT	61.841 13.868 61.873 13.932 ;
			RECT	62.009 13.868 62.041 13.932 ;
			RECT	62.177 13.868 62.209 13.932 ;
			RECT	62.345 13.868 62.377 13.932 ;
			RECT	62.513 13.868 62.545 13.932 ;
			RECT	62.681 13.868 62.713 13.932 ;
			RECT	62.849 13.868 62.881 13.932 ;
			RECT	63.017 13.868 63.049 13.932 ;
			RECT	63.185 13.868 63.217 13.932 ;
			RECT	63.353 13.868 63.385 13.932 ;
			RECT	63.521 13.868 63.553 13.932 ;
			RECT	63.689 13.868 63.721 13.932 ;
			RECT	63.857 13.868 63.889 13.932 ;
			RECT	64.025 13.868 64.057 13.932 ;
			RECT	64.193 13.868 64.225 13.932 ;
			RECT	64.361 13.868 64.393 13.932 ;
			RECT	64.529 13.868 64.561 13.932 ;
			RECT	64.697 13.868 64.729 13.932 ;
			RECT	64.865 13.868 64.897 13.932 ;
			RECT	65.033 13.868 65.065 13.932 ;
			RECT	65.201 13.868 65.233 13.932 ;
			RECT	65.369 13.868 65.401 13.932 ;
			RECT	65.537 13.868 65.569 13.932 ;
			RECT	65.705 13.868 65.737 13.932 ;
			RECT	65.873 13.868 65.905 13.932 ;
			RECT	66.041 13.868 66.073 13.932 ;
			RECT	66.209 13.868 66.241 13.932 ;
			RECT	66.377 13.868 66.409 13.932 ;
			RECT	66.545 13.868 66.577 13.932 ;
			RECT	66.713 13.868 66.745 13.932 ;
			RECT	66.881 13.868 66.913 13.932 ;
			RECT	67.049 13.868 67.081 13.932 ;
			RECT	67.217 13.868 67.249 13.932 ;
			RECT	67.385 13.868 67.417 13.932 ;
			RECT	67.553 13.868 67.585 13.932 ;
			RECT	67.721 13.868 67.753 13.932 ;
			RECT	67.889 13.868 67.921 13.932 ;
			RECT	68.057 13.868 68.089 13.932 ;
			RECT	68.225 13.868 68.257 13.932 ;
			RECT	68.393 13.868 68.425 13.932 ;
			RECT	68.561 13.868 68.593 13.932 ;
			RECT	68.729 13.868 68.761 13.932 ;
			RECT	68.897 13.868 68.929 13.932 ;
			RECT	69.065 13.868 69.097 13.932 ;
			RECT	69.233 13.868 69.265 13.932 ;
			RECT	69.401 13.868 69.433 13.932 ;
			RECT	69.569 13.868 69.601 13.932 ;
			RECT	69.737 13.868 69.769 13.932 ;
			RECT	69.905 13.868 69.937 13.932 ;
			RECT	70.073 13.868 70.105 13.932 ;
			RECT	70.241 13.868 70.273 13.932 ;
			RECT	70.409 13.868 70.441 13.932 ;
			RECT	70.577 13.868 70.609 13.932 ;
			RECT	70.745 13.868 70.777 13.932 ;
			RECT	70.913 13.868 70.945 13.932 ;
			RECT	71.081 13.868 71.113 13.932 ;
			RECT	71.249 13.868 71.281 13.932 ;
			RECT	71.417 13.868 71.449 13.932 ;
			RECT	71.585 13.868 71.617 13.932 ;
			RECT	71.753 13.868 71.785 13.932 ;
			RECT	71.921 13.868 71.953 13.932 ;
			RECT	72.089 13.868 72.121 13.932 ;
			RECT	72.257 13.868 72.289 13.932 ;
			RECT	72.425 13.868 72.457 13.932 ;
			RECT	72.593 13.868 72.625 13.932 ;
			RECT	72.761 13.868 72.793 13.932 ;
			RECT	72.929 13.868 72.961 13.932 ;
			RECT	73.097 13.868 73.129 13.932 ;
			RECT	73.265 13.868 73.297 13.932 ;
			RECT	73.433 13.868 73.465 13.932 ;
			RECT	73.601 13.868 73.633 13.932 ;
			RECT	73.769 13.868 73.801 13.932 ;
			RECT	73.937 13.868 73.969 13.932 ;
			RECT	74.105 13.868 74.137 13.932 ;
			RECT	74.273 13.868 74.305 13.932 ;
			RECT	74.441 13.868 74.473 13.932 ;
			RECT	74.609 13.868 74.641 13.932 ;
			RECT	74.777 13.868 74.809 13.932 ;
			RECT	74.945 13.868 74.977 13.932 ;
			RECT	75.113 13.868 75.145 13.932 ;
			RECT	75.281 13.868 75.313 13.932 ;
			RECT	75.449 13.868 75.481 13.932 ;
			RECT	75.617 13.868 75.649 13.932 ;
			RECT	75.785 13.868 75.817 13.932 ;
			RECT	75.953 13.868 75.985 13.932 ;
			RECT	76.121 13.868 76.153 13.932 ;
			RECT	76.289 13.868 76.321 13.932 ;
			RECT	76.457 13.868 76.489 13.932 ;
			RECT	76.625 13.868 76.657 13.932 ;
			RECT	76.793 13.868 76.825 13.932 ;
			RECT	76.961 13.868 76.993 13.932 ;
			RECT	77.129 13.868 77.161 13.932 ;
			RECT	77.297 13.868 77.329 13.932 ;
			RECT	77.465 13.868 77.497 13.932 ;
			RECT	77.633 13.868 77.665 13.932 ;
			RECT	77.801 13.868 77.833 13.932 ;
			RECT	77.969 13.868 78.001 13.932 ;
			RECT	78.137 13.868 78.169 13.932 ;
			RECT	78.305 13.868 78.337 13.932 ;
			RECT	78.473 13.868 78.505 13.932 ;
			RECT	78.641 13.868 78.673 13.932 ;
			RECT	78.809 13.868 78.841 13.932 ;
			RECT	78.977 13.868 79.009 13.932 ;
			RECT	79.145 13.868 79.177 13.932 ;
			RECT	79.313 13.868 79.345 13.932 ;
			RECT	79.481 13.868 79.513 13.932 ;
			RECT	79.649 13.868 79.681 13.932 ;
			RECT	79.817 13.868 79.849 13.932 ;
			RECT	79.985 13.868 80.017 13.932 ;
			RECT	80.153 13.868 80.185 13.932 ;
			RECT	80.321 13.868 80.353 13.932 ;
			RECT	80.489 13.868 80.521 13.932 ;
			RECT	80.657 13.868 80.689 13.932 ;
			RECT	80.825 13.868 80.857 13.932 ;
			RECT	80.993 13.868 81.025 13.932 ;
			RECT	81.161 13.868 81.193 13.932 ;
			RECT	81.329 13.868 81.361 13.932 ;
			RECT	81.497 13.868 81.529 13.932 ;
			RECT	81.665 13.868 81.697 13.932 ;
			RECT	81.833 13.868 81.865 13.932 ;
			RECT	82.001 13.868 82.033 13.932 ;
			RECT	82.169 13.868 82.201 13.932 ;
			RECT	82.337 13.868 82.369 13.932 ;
			RECT	82.505 13.868 82.537 13.932 ;
			RECT	82.673 13.868 82.705 13.932 ;
			RECT	82.841 13.868 82.873 13.932 ;
			RECT	83.009 13.868 83.041 13.932 ;
			RECT	83.177 13.868 83.209 13.932 ;
			RECT	83.345 13.868 83.377 13.932 ;
			RECT	83.513 13.868 83.545 13.932 ;
			RECT	83.681 13.868 83.713 13.932 ;
			RECT	83.849 13.868 83.881 13.932 ;
			RECT	84.017 13.868 84.049 13.932 ;
			RECT	84.185 13.868 84.217 13.932 ;
			RECT	84.353 13.868 84.385 13.932 ;
			RECT	84.521 13.868 84.553 13.932 ;
			RECT	84.689 13.868 84.721 13.932 ;
			RECT	84.857 13.868 84.889 13.932 ;
			RECT	85.025 13.868 85.057 13.932 ;
			RECT	85.193 13.868 85.225 13.932 ;
			RECT	85.361 13.868 85.393 13.932 ;
			RECT	85.529 13.868 85.561 13.932 ;
			RECT	85.697 13.868 85.729 13.932 ;
			RECT	85.865 13.868 85.897 13.932 ;
			RECT	86.033 13.868 86.065 13.932 ;
			RECT	86.201 13.868 86.233 13.932 ;
			RECT	86.369 13.868 86.401 13.932 ;
			RECT	86.537 13.868 86.569 13.932 ;
			RECT	86.705 13.868 86.737 13.932 ;
			RECT	86.873 13.868 86.905 13.932 ;
			RECT	87.041 13.868 87.073 13.932 ;
			RECT	87.209 13.868 87.241 13.932 ;
			RECT	87.377 13.868 87.409 13.932 ;
			RECT	87.545 13.868 87.577 13.932 ;
			RECT	87.713 13.868 87.745 13.932 ;
			RECT	87.881 13.868 87.913 13.932 ;
			RECT	88.049 13.868 88.081 13.932 ;
			RECT	88.217 13.868 88.249 13.932 ;
			RECT	88.385 13.868 88.417 13.932 ;
			RECT	88.553 13.868 88.585 13.932 ;
			RECT	88.721 13.868 88.753 13.932 ;
			RECT	88.889 13.868 88.921 13.932 ;
			RECT	89.057 13.868 89.089 13.932 ;
			RECT	89.225 13.868 89.257 13.932 ;
			RECT	89.393 13.868 89.425 13.932 ;
			RECT	89.561 13.868 89.593 13.932 ;
			RECT	89.729 13.868 89.761 13.932 ;
			RECT	89.897 13.868 89.929 13.932 ;
			RECT	90.065 13.868 90.097 13.932 ;
			RECT	90.233 13.868 90.265 13.932 ;
			RECT	90.401 13.868 90.433 13.932 ;
			RECT	90.569 13.868 90.601 13.932 ;
			RECT	90.737 13.868 90.769 13.932 ;
			RECT	90.905 13.868 90.937 13.932 ;
			RECT	91.073 13.868 91.105 13.932 ;
			RECT	91.241 13.868 91.273 13.932 ;
			RECT	91.409 13.868 91.441 13.932 ;
			RECT	91.577 13.868 91.609 13.932 ;
			RECT	91.745 13.868 91.777 13.932 ;
			RECT	91.913 13.868 91.945 13.932 ;
			RECT	92.081 13.868 92.113 13.932 ;
			RECT	92.249 13.868 92.281 13.932 ;
			RECT	92.417 13.868 92.449 13.932 ;
			RECT	92.585 13.868 92.617 13.932 ;
			RECT	92.753 13.868 92.785 13.932 ;
			RECT	92.921 13.868 92.953 13.932 ;
			RECT	93.089 13.868 93.121 13.932 ;
			RECT	93.257 13.868 93.289 13.932 ;
			RECT	93.425 13.868 93.457 13.932 ;
			RECT	93.593 13.868 93.625 13.932 ;
			RECT	93.761 13.868 93.793 13.932 ;
			RECT	93.929 13.868 93.961 13.932 ;
			RECT	94.097 13.868 94.129 13.932 ;
			RECT	94.265 13.868 94.297 13.932 ;
			RECT	94.433 13.868 94.465 13.932 ;
			RECT	94.601 13.868 94.633 13.932 ;
			RECT	94.769 13.868 94.801 13.932 ;
			RECT	94.937 13.868 94.969 13.932 ;
			RECT	95.105 13.868 95.137 13.932 ;
			RECT	95.273 13.868 95.305 13.932 ;
			RECT	95.441 13.868 95.473 13.932 ;
			RECT	95.609 13.868 95.641 13.932 ;
			RECT	95.777 13.868 95.809 13.932 ;
			RECT	95.945 13.868 95.977 13.932 ;
			RECT	96.113 13.868 96.145 13.932 ;
			RECT	96.281 13.868 96.313 13.932 ;
			RECT	96.449 13.868 96.481 13.932 ;
			RECT	96.617 13.868 96.649 13.932 ;
			RECT	96.785 13.868 96.817 13.932 ;
			RECT	96.953 13.868 96.985 13.932 ;
			RECT	97.121 13.868 97.153 13.932 ;
			RECT	97.289 13.868 97.321 13.932 ;
			RECT	97.457 13.868 97.489 13.932 ;
			RECT	97.625 13.868 97.657 13.932 ;
			RECT	97.793 13.868 97.825 13.932 ;
			RECT	97.961 13.868 97.993 13.932 ;
			RECT	98.129 13.868 98.161 13.932 ;
			RECT	98.297 13.868 98.329 13.932 ;
			RECT	98.465 13.868 98.497 13.932 ;
			RECT	98.633 13.868 98.665 13.932 ;
			RECT	98.801 13.868 98.833 13.932 ;
			RECT	98.969 13.868 99.001 13.932 ;
			RECT	99.137 13.868 99.169 13.932 ;
			RECT	99.305 13.868 99.337 13.932 ;
			RECT	99.473 13.868 99.505 13.932 ;
			RECT	99.641 13.868 99.673 13.932 ;
			RECT	99.809 13.868 99.841 13.932 ;
			RECT	99.977 13.868 100.009 13.932 ;
			RECT	100.145 13.868 100.177 13.932 ;
			RECT	100.313 13.868 100.345 13.932 ;
			RECT	100.481 13.868 100.513 13.932 ;
			RECT	100.649 13.868 100.681 13.932 ;
			RECT	100.817 13.868 100.849 13.932 ;
			RECT	100.985 13.868 101.017 13.932 ;
			RECT	101.153 13.868 101.185 13.932 ;
			RECT	101.321 13.868 101.353 13.932 ;
			RECT	101.489 13.868 101.521 13.932 ;
			RECT	101.657 13.868 101.689 13.932 ;
			RECT	101.825 13.868 101.857 13.932 ;
			RECT	101.993 13.868 102.025 13.932 ;
			RECT	102.123 13.884 102.155 13.916 ;
			RECT	102.245 13.889 102.277 13.921 ;
			RECT	102.375 13.868 102.407 13.932 ;
			RECT	103.795 13.868 103.827 13.932 ;
			RECT	103.925 13.889 103.957 13.921 ;
			RECT	104.047 13.884 104.079 13.916 ;
			RECT	104.177 13.868 104.209 13.932 ;
			RECT	104.345 13.868 104.377 13.932 ;
			RECT	104.513 13.868 104.545 13.932 ;
			RECT	104.681 13.868 104.713 13.932 ;
			RECT	104.849 13.868 104.881 13.932 ;
			RECT	105.017 13.868 105.049 13.932 ;
			RECT	105.185 13.868 105.217 13.932 ;
			RECT	105.353 13.868 105.385 13.932 ;
			RECT	105.521 13.868 105.553 13.932 ;
			RECT	105.689 13.868 105.721 13.932 ;
			RECT	105.857 13.868 105.889 13.932 ;
			RECT	106.025 13.868 106.057 13.932 ;
			RECT	106.193 13.868 106.225 13.932 ;
			RECT	106.361 13.868 106.393 13.932 ;
			RECT	106.529 13.868 106.561 13.932 ;
			RECT	106.697 13.868 106.729 13.932 ;
			RECT	106.865 13.868 106.897 13.932 ;
			RECT	107.033 13.868 107.065 13.932 ;
			RECT	107.201 13.868 107.233 13.932 ;
			RECT	107.369 13.868 107.401 13.932 ;
			RECT	107.537 13.868 107.569 13.932 ;
			RECT	107.705 13.868 107.737 13.932 ;
			RECT	107.873 13.868 107.905 13.932 ;
			RECT	108.041 13.868 108.073 13.932 ;
			RECT	108.209 13.868 108.241 13.932 ;
			RECT	108.377 13.868 108.409 13.932 ;
			RECT	108.545 13.868 108.577 13.932 ;
			RECT	108.713 13.868 108.745 13.932 ;
			RECT	108.881 13.868 108.913 13.932 ;
			RECT	109.049 13.868 109.081 13.932 ;
			RECT	109.217 13.868 109.249 13.932 ;
			RECT	109.385 13.868 109.417 13.932 ;
			RECT	109.553 13.868 109.585 13.932 ;
			RECT	109.721 13.868 109.753 13.932 ;
			RECT	109.889 13.868 109.921 13.932 ;
			RECT	110.057 13.868 110.089 13.932 ;
			RECT	110.225 13.868 110.257 13.932 ;
			RECT	110.393 13.868 110.425 13.932 ;
			RECT	110.561 13.868 110.593 13.932 ;
			RECT	110.729 13.868 110.761 13.932 ;
			RECT	110.897 13.868 110.929 13.932 ;
			RECT	111.065 13.868 111.097 13.932 ;
			RECT	111.233 13.868 111.265 13.932 ;
			RECT	111.401 13.868 111.433 13.932 ;
			RECT	111.569 13.868 111.601 13.932 ;
			RECT	111.737 13.868 111.769 13.932 ;
			RECT	111.905 13.868 111.937 13.932 ;
			RECT	112.073 13.868 112.105 13.932 ;
			RECT	112.241 13.868 112.273 13.932 ;
			RECT	112.409 13.868 112.441 13.932 ;
			RECT	112.577 13.868 112.609 13.932 ;
			RECT	112.745 13.868 112.777 13.932 ;
			RECT	112.913 13.868 112.945 13.932 ;
			RECT	113.081 13.868 113.113 13.932 ;
			RECT	113.249 13.868 113.281 13.932 ;
			RECT	113.417 13.868 113.449 13.932 ;
			RECT	113.585 13.868 113.617 13.932 ;
			RECT	113.753 13.868 113.785 13.932 ;
			RECT	113.921 13.868 113.953 13.932 ;
			RECT	114.089 13.868 114.121 13.932 ;
			RECT	114.257 13.868 114.289 13.932 ;
			RECT	114.425 13.868 114.457 13.932 ;
			RECT	114.593 13.868 114.625 13.932 ;
			RECT	114.761 13.868 114.793 13.932 ;
			RECT	114.929 13.868 114.961 13.932 ;
			RECT	115.097 13.868 115.129 13.932 ;
			RECT	115.265 13.868 115.297 13.932 ;
			RECT	115.433 13.868 115.465 13.932 ;
			RECT	115.601 13.868 115.633 13.932 ;
			RECT	115.769 13.868 115.801 13.932 ;
			RECT	115.937 13.868 115.969 13.932 ;
			RECT	116.105 13.868 116.137 13.932 ;
			RECT	116.273 13.868 116.305 13.932 ;
			RECT	116.441 13.868 116.473 13.932 ;
			RECT	116.609 13.868 116.641 13.932 ;
			RECT	116.777 13.868 116.809 13.932 ;
			RECT	116.945 13.868 116.977 13.932 ;
			RECT	117.113 13.868 117.145 13.932 ;
			RECT	117.281 13.868 117.313 13.932 ;
			RECT	117.449 13.868 117.481 13.932 ;
			RECT	117.617 13.868 117.649 13.932 ;
			RECT	117.785 13.868 117.817 13.932 ;
			RECT	117.953 13.868 117.985 13.932 ;
			RECT	118.121 13.868 118.153 13.932 ;
			RECT	118.289 13.868 118.321 13.932 ;
			RECT	118.457 13.868 118.489 13.932 ;
			RECT	118.625 13.868 118.657 13.932 ;
			RECT	118.793 13.868 118.825 13.932 ;
			RECT	118.961 13.868 118.993 13.932 ;
			RECT	119.129 13.868 119.161 13.932 ;
			RECT	119.297 13.868 119.329 13.932 ;
			RECT	119.465 13.868 119.497 13.932 ;
			RECT	119.633 13.868 119.665 13.932 ;
			RECT	119.801 13.868 119.833 13.932 ;
			RECT	119.969 13.868 120.001 13.932 ;
			RECT	120.137 13.868 120.169 13.932 ;
			RECT	120.305 13.868 120.337 13.932 ;
			RECT	120.473 13.868 120.505 13.932 ;
			RECT	120.641 13.868 120.673 13.932 ;
			RECT	120.809 13.868 120.841 13.932 ;
			RECT	120.977 13.868 121.009 13.932 ;
			RECT	121.145 13.868 121.177 13.932 ;
			RECT	121.313 13.868 121.345 13.932 ;
			RECT	121.481 13.868 121.513 13.932 ;
			RECT	121.649 13.868 121.681 13.932 ;
			RECT	121.817 13.868 121.849 13.932 ;
			RECT	121.985 13.868 122.017 13.932 ;
			RECT	122.153 13.868 122.185 13.932 ;
			RECT	122.321 13.868 122.353 13.932 ;
			RECT	122.489 13.868 122.521 13.932 ;
			RECT	122.657 13.868 122.689 13.932 ;
			RECT	122.825 13.868 122.857 13.932 ;
			RECT	122.993 13.868 123.025 13.932 ;
			RECT	123.161 13.868 123.193 13.932 ;
			RECT	123.329 13.868 123.361 13.932 ;
			RECT	123.497 13.868 123.529 13.932 ;
			RECT	123.665 13.868 123.697 13.932 ;
			RECT	123.833 13.868 123.865 13.932 ;
			RECT	124.001 13.868 124.033 13.932 ;
			RECT	124.169 13.868 124.201 13.932 ;
			RECT	124.337 13.868 124.369 13.932 ;
			RECT	124.505 13.868 124.537 13.932 ;
			RECT	124.673 13.868 124.705 13.932 ;
			RECT	124.841 13.868 124.873 13.932 ;
			RECT	125.009 13.868 125.041 13.932 ;
			RECT	125.177 13.868 125.209 13.932 ;
			RECT	125.345 13.868 125.377 13.932 ;
			RECT	125.513 13.868 125.545 13.932 ;
			RECT	125.681 13.868 125.713 13.932 ;
			RECT	125.849 13.868 125.881 13.932 ;
			RECT	126.017 13.868 126.049 13.932 ;
			RECT	126.185 13.868 126.217 13.932 ;
			RECT	126.353 13.868 126.385 13.932 ;
			RECT	126.521 13.868 126.553 13.932 ;
			RECT	126.689 13.868 126.721 13.932 ;
			RECT	126.857 13.868 126.889 13.932 ;
			RECT	127.025 13.868 127.057 13.932 ;
			RECT	127.193 13.868 127.225 13.932 ;
			RECT	127.361 13.868 127.393 13.932 ;
			RECT	127.529 13.868 127.561 13.932 ;
			RECT	127.697 13.868 127.729 13.932 ;
			RECT	127.865 13.868 127.897 13.932 ;
			RECT	128.033 13.868 128.065 13.932 ;
			RECT	128.201 13.868 128.233 13.932 ;
			RECT	128.369 13.868 128.401 13.932 ;
			RECT	128.537 13.868 128.569 13.932 ;
			RECT	128.705 13.868 128.737 13.932 ;
			RECT	128.873 13.868 128.905 13.932 ;
			RECT	129.041 13.868 129.073 13.932 ;
			RECT	129.209 13.868 129.241 13.932 ;
			RECT	129.377 13.868 129.409 13.932 ;
			RECT	129.545 13.868 129.577 13.932 ;
			RECT	129.713 13.868 129.745 13.932 ;
			RECT	129.881 13.868 129.913 13.932 ;
			RECT	130.049 13.868 130.081 13.932 ;
			RECT	130.217 13.868 130.249 13.932 ;
			RECT	130.385 13.868 130.417 13.932 ;
			RECT	130.553 13.868 130.585 13.932 ;
			RECT	130.721 13.868 130.753 13.932 ;
			RECT	130.889 13.868 130.921 13.932 ;
			RECT	131.057 13.868 131.089 13.932 ;
			RECT	131.225 13.868 131.257 13.932 ;
			RECT	131.393 13.868 131.425 13.932 ;
			RECT	131.561 13.868 131.593 13.932 ;
			RECT	131.729 13.868 131.761 13.932 ;
			RECT	131.897 13.868 131.929 13.932 ;
			RECT	132.065 13.868 132.097 13.932 ;
			RECT	132.233 13.868 132.265 13.932 ;
			RECT	132.401 13.868 132.433 13.932 ;
			RECT	132.569 13.868 132.601 13.932 ;
			RECT	132.737 13.868 132.769 13.932 ;
			RECT	132.905 13.868 132.937 13.932 ;
			RECT	133.073 13.868 133.105 13.932 ;
			RECT	133.241 13.868 133.273 13.932 ;
			RECT	133.409 13.868 133.441 13.932 ;
			RECT	133.577 13.868 133.609 13.932 ;
			RECT	133.745 13.868 133.777 13.932 ;
			RECT	133.913 13.868 133.945 13.932 ;
			RECT	134.081 13.868 134.113 13.932 ;
			RECT	134.249 13.868 134.281 13.932 ;
			RECT	134.417 13.868 134.449 13.932 ;
			RECT	134.585 13.868 134.617 13.932 ;
			RECT	134.753 13.868 134.785 13.932 ;
			RECT	134.921 13.868 134.953 13.932 ;
			RECT	135.089 13.868 135.121 13.932 ;
			RECT	135.257 13.868 135.289 13.932 ;
			RECT	135.425 13.868 135.457 13.932 ;
			RECT	135.593 13.868 135.625 13.932 ;
			RECT	135.761 13.868 135.793 13.932 ;
			RECT	135.929 13.868 135.961 13.932 ;
			RECT	136.097 13.868 136.129 13.932 ;
			RECT	136.265 13.868 136.297 13.932 ;
			RECT	136.433 13.868 136.465 13.932 ;
			RECT	136.601 13.868 136.633 13.932 ;
			RECT	136.769 13.868 136.801 13.932 ;
			RECT	136.937 13.868 136.969 13.932 ;
			RECT	137.105 13.868 137.137 13.932 ;
			RECT	137.273 13.868 137.305 13.932 ;
			RECT	137.441 13.868 137.473 13.932 ;
			RECT	137.609 13.868 137.641 13.932 ;
			RECT	137.777 13.868 137.809 13.932 ;
			RECT	137.945 13.868 137.977 13.932 ;
			RECT	138.113 13.868 138.145 13.932 ;
			RECT	138.281 13.868 138.313 13.932 ;
			RECT	138.449 13.868 138.481 13.932 ;
			RECT	138.617 13.868 138.649 13.932 ;
			RECT	138.785 13.868 138.817 13.932 ;
			RECT	138.953 13.868 138.985 13.932 ;
			RECT	139.121 13.868 139.153 13.932 ;
			RECT	139.289 13.868 139.321 13.932 ;
			RECT	139.457 13.868 139.489 13.932 ;
			RECT	139.625 13.868 139.657 13.932 ;
			RECT	139.793 13.868 139.825 13.932 ;
			RECT	139.961 13.868 139.993 13.932 ;
			RECT	140.129 13.868 140.161 13.932 ;
			RECT	140.297 13.868 140.329 13.932 ;
			RECT	140.465 13.868 140.497 13.932 ;
			RECT	140.633 13.868 140.665 13.932 ;
			RECT	140.801 13.868 140.833 13.932 ;
			RECT	140.969 13.868 141.001 13.932 ;
			RECT	141.137 13.868 141.169 13.932 ;
			RECT	141.305 13.868 141.337 13.932 ;
			RECT	141.473 13.868 141.505 13.932 ;
			RECT	141.641 13.868 141.673 13.932 ;
			RECT	141.809 13.868 141.841 13.932 ;
			RECT	141.977 13.868 142.009 13.932 ;
			RECT	142.145 13.868 142.177 13.932 ;
			RECT	142.313 13.868 142.345 13.932 ;
			RECT	142.481 13.868 142.513 13.932 ;
			RECT	142.649 13.868 142.681 13.932 ;
			RECT	142.817 13.868 142.849 13.932 ;
			RECT	142.985 13.868 143.017 13.932 ;
			RECT	143.153 13.868 143.185 13.932 ;
			RECT	143.321 13.868 143.353 13.932 ;
			RECT	143.489 13.868 143.521 13.932 ;
			RECT	143.657 13.868 143.689 13.932 ;
			RECT	143.825 13.868 143.857 13.932 ;
			RECT	143.993 13.868 144.025 13.932 ;
			RECT	144.161 13.868 144.193 13.932 ;
			RECT	144.329 13.868 144.361 13.932 ;
			RECT	144.497 13.868 144.529 13.932 ;
			RECT	144.665 13.868 144.697 13.932 ;
			RECT	144.833 13.868 144.865 13.932 ;
			RECT	145.001 13.868 145.033 13.932 ;
			RECT	145.169 13.868 145.201 13.932 ;
			RECT	145.337 13.868 145.369 13.932 ;
			RECT	145.505 13.868 145.537 13.932 ;
			RECT	145.673 13.868 145.705 13.932 ;
			RECT	145.841 13.868 145.873 13.932 ;
			RECT	146.009 13.868 146.041 13.932 ;
			RECT	146.177 13.868 146.209 13.932 ;
			RECT	146.345 13.868 146.377 13.932 ;
			RECT	146.513 13.868 146.545 13.932 ;
			RECT	146.681 13.868 146.713 13.932 ;
			RECT	146.849 13.868 146.881 13.932 ;
			RECT	147.017 13.868 147.049 13.932 ;
			RECT	147.185 13.868 147.217 13.932 ;
			RECT	147.316 13.884 147.348 13.916 ;
			RECT	147.437 13.884 147.469 13.916 ;
			RECT	147.567 13.868 147.599 13.932 ;
			RECT	149.879 13.868 149.911 13.932 ;
			RECT	151.13 13.868 151.194 13.932 ;
			RECT	151.81 13.868 151.842 13.932 ;
			RECT	152.249 13.868 152.281 13.932 ;
			RECT	153.56 13.868 153.624 13.932 ;
			RECT	156.601 13.868 156.633 13.932 ;
			RECT	156.731 13.884 156.763 13.916 ;
			RECT	156.852 13.884 156.884 13.916 ;
			RECT	156.983 13.868 157.015 13.932 ;
			RECT	157.151 13.868 157.183 13.932 ;
			RECT	157.319 13.868 157.351 13.932 ;
			RECT	157.487 13.868 157.519 13.932 ;
			RECT	157.655 13.868 157.687 13.932 ;
			RECT	157.823 13.868 157.855 13.932 ;
			RECT	157.991 13.868 158.023 13.932 ;
			RECT	158.159 13.868 158.191 13.932 ;
			RECT	158.327 13.868 158.359 13.932 ;
			RECT	158.495 13.868 158.527 13.932 ;
			RECT	158.663 13.868 158.695 13.932 ;
			RECT	158.831 13.868 158.863 13.932 ;
			RECT	158.999 13.868 159.031 13.932 ;
			RECT	159.167 13.868 159.199 13.932 ;
			RECT	159.335 13.868 159.367 13.932 ;
			RECT	159.503 13.868 159.535 13.932 ;
			RECT	159.671 13.868 159.703 13.932 ;
			RECT	159.839 13.868 159.871 13.932 ;
			RECT	160.007 13.868 160.039 13.932 ;
			RECT	160.175 13.868 160.207 13.932 ;
			RECT	160.343 13.868 160.375 13.932 ;
			RECT	160.511 13.868 160.543 13.932 ;
			RECT	160.679 13.868 160.711 13.932 ;
			RECT	160.847 13.868 160.879 13.932 ;
			RECT	161.015 13.868 161.047 13.932 ;
			RECT	161.183 13.868 161.215 13.932 ;
			RECT	161.351 13.868 161.383 13.932 ;
			RECT	161.519 13.868 161.551 13.932 ;
			RECT	161.687 13.868 161.719 13.932 ;
			RECT	161.855 13.868 161.887 13.932 ;
			RECT	162.023 13.868 162.055 13.932 ;
			RECT	162.191 13.868 162.223 13.932 ;
			RECT	162.359 13.868 162.391 13.932 ;
			RECT	162.527 13.868 162.559 13.932 ;
			RECT	162.695 13.868 162.727 13.932 ;
			RECT	162.863 13.868 162.895 13.932 ;
			RECT	163.031 13.868 163.063 13.932 ;
			RECT	163.199 13.868 163.231 13.932 ;
			RECT	163.367 13.868 163.399 13.932 ;
			RECT	163.535 13.868 163.567 13.932 ;
			RECT	163.703 13.868 163.735 13.932 ;
			RECT	163.871 13.868 163.903 13.932 ;
			RECT	164.039 13.868 164.071 13.932 ;
			RECT	164.207 13.868 164.239 13.932 ;
			RECT	164.375 13.868 164.407 13.932 ;
			RECT	164.543 13.868 164.575 13.932 ;
			RECT	164.711 13.868 164.743 13.932 ;
			RECT	164.879 13.868 164.911 13.932 ;
			RECT	165.047 13.868 165.079 13.932 ;
			RECT	165.215 13.868 165.247 13.932 ;
			RECT	165.383 13.868 165.415 13.932 ;
			RECT	165.551 13.868 165.583 13.932 ;
			RECT	165.719 13.868 165.751 13.932 ;
			RECT	165.887 13.868 165.919 13.932 ;
			RECT	166.055 13.868 166.087 13.932 ;
			RECT	166.223 13.868 166.255 13.932 ;
			RECT	166.391 13.868 166.423 13.932 ;
			RECT	166.559 13.868 166.591 13.932 ;
			RECT	166.727 13.868 166.759 13.932 ;
			RECT	166.895 13.868 166.927 13.932 ;
			RECT	167.063 13.868 167.095 13.932 ;
			RECT	167.231 13.868 167.263 13.932 ;
			RECT	167.399 13.868 167.431 13.932 ;
			RECT	167.567 13.868 167.599 13.932 ;
			RECT	167.735 13.868 167.767 13.932 ;
			RECT	167.903 13.868 167.935 13.932 ;
			RECT	168.071 13.868 168.103 13.932 ;
			RECT	168.239 13.868 168.271 13.932 ;
			RECT	168.407 13.868 168.439 13.932 ;
			RECT	168.575 13.868 168.607 13.932 ;
			RECT	168.743 13.868 168.775 13.932 ;
			RECT	168.911 13.868 168.943 13.932 ;
			RECT	169.079 13.868 169.111 13.932 ;
			RECT	169.247 13.868 169.279 13.932 ;
			RECT	169.415 13.868 169.447 13.932 ;
			RECT	169.583 13.868 169.615 13.932 ;
			RECT	169.751 13.868 169.783 13.932 ;
			RECT	169.919 13.868 169.951 13.932 ;
			RECT	170.087 13.868 170.119 13.932 ;
			RECT	170.255 13.868 170.287 13.932 ;
			RECT	170.423 13.868 170.455 13.932 ;
			RECT	170.591 13.868 170.623 13.932 ;
			RECT	170.759 13.868 170.791 13.932 ;
			RECT	170.927 13.868 170.959 13.932 ;
			RECT	171.095 13.868 171.127 13.932 ;
			RECT	171.263 13.868 171.295 13.932 ;
			RECT	171.431 13.868 171.463 13.932 ;
			RECT	171.599 13.868 171.631 13.932 ;
			RECT	171.767 13.868 171.799 13.932 ;
			RECT	171.935 13.868 171.967 13.932 ;
			RECT	172.103 13.868 172.135 13.932 ;
			RECT	172.271 13.868 172.303 13.932 ;
			RECT	172.439 13.868 172.471 13.932 ;
			RECT	172.607 13.868 172.639 13.932 ;
			RECT	172.775 13.868 172.807 13.932 ;
			RECT	172.943 13.868 172.975 13.932 ;
			RECT	173.111 13.868 173.143 13.932 ;
			RECT	173.279 13.868 173.311 13.932 ;
			RECT	173.447 13.868 173.479 13.932 ;
			RECT	173.615 13.868 173.647 13.932 ;
			RECT	173.783 13.868 173.815 13.932 ;
			RECT	173.951 13.868 173.983 13.932 ;
			RECT	174.119 13.868 174.151 13.932 ;
			RECT	174.287 13.868 174.319 13.932 ;
			RECT	174.455 13.868 174.487 13.932 ;
			RECT	174.623 13.868 174.655 13.932 ;
			RECT	174.791 13.868 174.823 13.932 ;
			RECT	174.959 13.868 174.991 13.932 ;
			RECT	175.127 13.868 175.159 13.932 ;
			RECT	175.295 13.868 175.327 13.932 ;
			RECT	175.463 13.868 175.495 13.932 ;
			RECT	175.631 13.868 175.663 13.932 ;
			RECT	175.799 13.868 175.831 13.932 ;
			RECT	175.967 13.868 175.999 13.932 ;
			RECT	176.135 13.868 176.167 13.932 ;
			RECT	176.303 13.868 176.335 13.932 ;
			RECT	176.471 13.868 176.503 13.932 ;
			RECT	176.639 13.868 176.671 13.932 ;
			RECT	176.807 13.868 176.839 13.932 ;
			RECT	176.975 13.868 177.007 13.932 ;
			RECT	177.143 13.868 177.175 13.932 ;
			RECT	177.311 13.868 177.343 13.932 ;
			RECT	177.479 13.868 177.511 13.932 ;
			RECT	177.647 13.868 177.679 13.932 ;
			RECT	177.815 13.868 177.847 13.932 ;
			RECT	177.983 13.868 178.015 13.932 ;
			RECT	178.151 13.868 178.183 13.932 ;
			RECT	178.319 13.868 178.351 13.932 ;
			RECT	178.487 13.868 178.519 13.932 ;
			RECT	178.655 13.868 178.687 13.932 ;
			RECT	178.823 13.868 178.855 13.932 ;
			RECT	178.991 13.868 179.023 13.932 ;
			RECT	179.159 13.868 179.191 13.932 ;
			RECT	179.327 13.868 179.359 13.932 ;
			RECT	179.495 13.868 179.527 13.932 ;
			RECT	179.663 13.868 179.695 13.932 ;
			RECT	179.831 13.868 179.863 13.932 ;
			RECT	179.999 13.868 180.031 13.932 ;
			RECT	180.167 13.868 180.199 13.932 ;
			RECT	180.335 13.868 180.367 13.932 ;
			RECT	180.503 13.868 180.535 13.932 ;
			RECT	180.671 13.868 180.703 13.932 ;
			RECT	180.839 13.868 180.871 13.932 ;
			RECT	181.007 13.868 181.039 13.932 ;
			RECT	181.175 13.868 181.207 13.932 ;
			RECT	181.343 13.868 181.375 13.932 ;
			RECT	181.511 13.868 181.543 13.932 ;
			RECT	181.679 13.868 181.711 13.932 ;
			RECT	181.847 13.868 181.879 13.932 ;
			RECT	182.015 13.868 182.047 13.932 ;
			RECT	182.183 13.868 182.215 13.932 ;
			RECT	182.351 13.868 182.383 13.932 ;
			RECT	182.519 13.868 182.551 13.932 ;
			RECT	182.687 13.868 182.719 13.932 ;
			RECT	182.855 13.868 182.887 13.932 ;
			RECT	183.023 13.868 183.055 13.932 ;
			RECT	183.191 13.868 183.223 13.932 ;
			RECT	183.359 13.868 183.391 13.932 ;
			RECT	183.527 13.868 183.559 13.932 ;
			RECT	183.695 13.868 183.727 13.932 ;
			RECT	183.863 13.868 183.895 13.932 ;
			RECT	184.031 13.868 184.063 13.932 ;
			RECT	184.199 13.868 184.231 13.932 ;
			RECT	184.367 13.868 184.399 13.932 ;
			RECT	184.535 13.868 184.567 13.932 ;
			RECT	184.703 13.868 184.735 13.932 ;
			RECT	184.871 13.868 184.903 13.932 ;
			RECT	185.039 13.868 185.071 13.932 ;
			RECT	185.207 13.868 185.239 13.932 ;
			RECT	185.375 13.868 185.407 13.932 ;
			RECT	185.543 13.868 185.575 13.932 ;
			RECT	185.711 13.868 185.743 13.932 ;
			RECT	185.879 13.868 185.911 13.932 ;
			RECT	186.047 13.868 186.079 13.932 ;
			RECT	186.215 13.868 186.247 13.932 ;
			RECT	186.383 13.868 186.415 13.932 ;
			RECT	186.551 13.868 186.583 13.932 ;
			RECT	186.719 13.868 186.751 13.932 ;
			RECT	186.887 13.868 186.919 13.932 ;
			RECT	187.055 13.868 187.087 13.932 ;
			RECT	187.223 13.868 187.255 13.932 ;
			RECT	187.391 13.868 187.423 13.932 ;
			RECT	187.559 13.868 187.591 13.932 ;
			RECT	187.727 13.868 187.759 13.932 ;
			RECT	187.895 13.868 187.927 13.932 ;
			RECT	188.063 13.868 188.095 13.932 ;
			RECT	188.231 13.868 188.263 13.932 ;
			RECT	188.399 13.868 188.431 13.932 ;
			RECT	188.567 13.868 188.599 13.932 ;
			RECT	188.735 13.868 188.767 13.932 ;
			RECT	188.903 13.868 188.935 13.932 ;
			RECT	189.071 13.868 189.103 13.932 ;
			RECT	189.239 13.868 189.271 13.932 ;
			RECT	189.407 13.868 189.439 13.932 ;
			RECT	189.575 13.868 189.607 13.932 ;
			RECT	189.743 13.868 189.775 13.932 ;
			RECT	189.911 13.868 189.943 13.932 ;
			RECT	190.079 13.868 190.111 13.932 ;
			RECT	190.247 13.868 190.279 13.932 ;
			RECT	190.415 13.868 190.447 13.932 ;
			RECT	190.583 13.868 190.615 13.932 ;
			RECT	190.751 13.868 190.783 13.932 ;
			RECT	190.919 13.868 190.951 13.932 ;
			RECT	191.087 13.868 191.119 13.932 ;
			RECT	191.255 13.868 191.287 13.932 ;
			RECT	191.423 13.868 191.455 13.932 ;
			RECT	191.591 13.868 191.623 13.932 ;
			RECT	191.759 13.868 191.791 13.932 ;
			RECT	191.927 13.868 191.959 13.932 ;
			RECT	192.095 13.868 192.127 13.932 ;
			RECT	192.263 13.868 192.295 13.932 ;
			RECT	192.431 13.868 192.463 13.932 ;
			RECT	192.599 13.868 192.631 13.932 ;
			RECT	192.767 13.868 192.799 13.932 ;
			RECT	192.935 13.868 192.967 13.932 ;
			RECT	193.103 13.868 193.135 13.932 ;
			RECT	193.271 13.868 193.303 13.932 ;
			RECT	193.439 13.868 193.471 13.932 ;
			RECT	193.607 13.868 193.639 13.932 ;
			RECT	193.775 13.868 193.807 13.932 ;
			RECT	193.943 13.868 193.975 13.932 ;
			RECT	194.111 13.868 194.143 13.932 ;
			RECT	194.279 13.868 194.311 13.932 ;
			RECT	194.447 13.868 194.479 13.932 ;
			RECT	194.615 13.868 194.647 13.932 ;
			RECT	194.783 13.868 194.815 13.932 ;
			RECT	194.951 13.868 194.983 13.932 ;
			RECT	195.119 13.868 195.151 13.932 ;
			RECT	195.287 13.868 195.319 13.932 ;
			RECT	195.455 13.868 195.487 13.932 ;
			RECT	195.623 13.868 195.655 13.932 ;
			RECT	195.791 13.868 195.823 13.932 ;
			RECT	195.959 13.868 195.991 13.932 ;
			RECT	196.127 13.868 196.159 13.932 ;
			RECT	196.295 13.868 196.327 13.932 ;
			RECT	196.463 13.868 196.495 13.932 ;
			RECT	196.631 13.868 196.663 13.932 ;
			RECT	196.799 13.868 196.831 13.932 ;
			RECT	196.967 13.868 196.999 13.932 ;
			RECT	197.135 13.868 197.167 13.932 ;
			RECT	197.303 13.868 197.335 13.932 ;
			RECT	197.471 13.868 197.503 13.932 ;
			RECT	197.639 13.868 197.671 13.932 ;
			RECT	197.807 13.868 197.839 13.932 ;
			RECT	197.975 13.868 198.007 13.932 ;
			RECT	198.143 13.868 198.175 13.932 ;
			RECT	198.311 13.868 198.343 13.932 ;
			RECT	198.479 13.868 198.511 13.932 ;
			RECT	198.647 13.868 198.679 13.932 ;
			RECT	198.815 13.868 198.847 13.932 ;
			RECT	198.983 13.868 199.015 13.932 ;
			RECT	199.151 13.868 199.183 13.932 ;
			RECT	199.319 13.868 199.351 13.932 ;
			RECT	199.487 13.868 199.519 13.932 ;
			RECT	199.655 13.868 199.687 13.932 ;
			RECT	199.823 13.868 199.855 13.932 ;
			RECT	199.991 13.868 200.023 13.932 ;
			RECT	200.121 13.884 200.153 13.916 ;
			RECT	200.243 13.889 200.275 13.921 ;
			RECT	200.373 13.868 200.405 13.932 ;
			RECT	200.9 13.868 200.932 13.932 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 11.92 201.665 12.04 ;
			LAYER	J3 ;
			RECT	0.755 11.948 0.787 12.012 ;
			RECT	1.645 11.948 1.709 12.012 ;
			RECT	2.323 11.948 2.387 12.012 ;
			RECT	3.438 11.948 3.47 12.012 ;
			RECT	3.585 11.948 3.617 12.012 ;
			RECT	4.195 11.948 4.227 12.012 ;
			RECT	4.72 11.948 4.752 12.012 ;
			RECT	4.944 11.948 5.008 12.012 ;
			RECT	5.267 11.948 5.299 12.012 ;
			RECT	5.797 11.948 5.829 12.012 ;
			RECT	5.927 11.969 5.959 12.001 ;
			RECT	6.049 11.964 6.081 11.996 ;
			RECT	6.179 11.948 6.211 12.012 ;
			RECT	6.347 11.948 6.379 12.012 ;
			RECT	6.515 11.948 6.547 12.012 ;
			RECT	6.683 11.948 6.715 12.012 ;
			RECT	6.851 11.948 6.883 12.012 ;
			RECT	7.019 11.948 7.051 12.012 ;
			RECT	7.187 11.948 7.219 12.012 ;
			RECT	7.355 11.948 7.387 12.012 ;
			RECT	7.523 11.948 7.555 12.012 ;
			RECT	7.691 11.948 7.723 12.012 ;
			RECT	7.859 11.948 7.891 12.012 ;
			RECT	8.027 11.948 8.059 12.012 ;
			RECT	8.195 11.948 8.227 12.012 ;
			RECT	8.363 11.948 8.395 12.012 ;
			RECT	8.531 11.948 8.563 12.012 ;
			RECT	8.699 11.948 8.731 12.012 ;
			RECT	8.867 11.948 8.899 12.012 ;
			RECT	9.035 11.948 9.067 12.012 ;
			RECT	9.203 11.948 9.235 12.012 ;
			RECT	9.371 11.948 9.403 12.012 ;
			RECT	9.539 11.948 9.571 12.012 ;
			RECT	9.707 11.948 9.739 12.012 ;
			RECT	9.875 11.948 9.907 12.012 ;
			RECT	10.043 11.948 10.075 12.012 ;
			RECT	10.211 11.948 10.243 12.012 ;
			RECT	10.379 11.948 10.411 12.012 ;
			RECT	10.547 11.948 10.579 12.012 ;
			RECT	10.715 11.948 10.747 12.012 ;
			RECT	10.883 11.948 10.915 12.012 ;
			RECT	11.051 11.948 11.083 12.012 ;
			RECT	11.219 11.948 11.251 12.012 ;
			RECT	11.387 11.948 11.419 12.012 ;
			RECT	11.555 11.948 11.587 12.012 ;
			RECT	11.723 11.948 11.755 12.012 ;
			RECT	11.891 11.948 11.923 12.012 ;
			RECT	12.059 11.948 12.091 12.012 ;
			RECT	12.227 11.948 12.259 12.012 ;
			RECT	12.395 11.948 12.427 12.012 ;
			RECT	12.563 11.948 12.595 12.012 ;
			RECT	12.731 11.948 12.763 12.012 ;
			RECT	12.899 11.948 12.931 12.012 ;
			RECT	13.067 11.948 13.099 12.012 ;
			RECT	13.235 11.948 13.267 12.012 ;
			RECT	13.403 11.948 13.435 12.012 ;
			RECT	13.571 11.948 13.603 12.012 ;
			RECT	13.739 11.948 13.771 12.012 ;
			RECT	13.907 11.948 13.939 12.012 ;
			RECT	14.075 11.948 14.107 12.012 ;
			RECT	14.243 11.948 14.275 12.012 ;
			RECT	14.411 11.948 14.443 12.012 ;
			RECT	14.579 11.948 14.611 12.012 ;
			RECT	14.747 11.948 14.779 12.012 ;
			RECT	14.915 11.948 14.947 12.012 ;
			RECT	15.083 11.948 15.115 12.012 ;
			RECT	15.251 11.948 15.283 12.012 ;
			RECT	15.419 11.948 15.451 12.012 ;
			RECT	15.587 11.948 15.619 12.012 ;
			RECT	15.755 11.948 15.787 12.012 ;
			RECT	15.923 11.948 15.955 12.012 ;
			RECT	16.091 11.948 16.123 12.012 ;
			RECT	16.259 11.948 16.291 12.012 ;
			RECT	16.427 11.948 16.459 12.012 ;
			RECT	16.595 11.948 16.627 12.012 ;
			RECT	16.763 11.948 16.795 12.012 ;
			RECT	16.931 11.948 16.963 12.012 ;
			RECT	17.099 11.948 17.131 12.012 ;
			RECT	17.267 11.948 17.299 12.012 ;
			RECT	17.435 11.948 17.467 12.012 ;
			RECT	17.603 11.948 17.635 12.012 ;
			RECT	17.771 11.948 17.803 12.012 ;
			RECT	17.939 11.948 17.971 12.012 ;
			RECT	18.107 11.948 18.139 12.012 ;
			RECT	18.275 11.948 18.307 12.012 ;
			RECT	18.443 11.948 18.475 12.012 ;
			RECT	18.611 11.948 18.643 12.012 ;
			RECT	18.779 11.948 18.811 12.012 ;
			RECT	18.947 11.948 18.979 12.012 ;
			RECT	19.115 11.948 19.147 12.012 ;
			RECT	19.283 11.948 19.315 12.012 ;
			RECT	19.451 11.948 19.483 12.012 ;
			RECT	19.619 11.948 19.651 12.012 ;
			RECT	19.787 11.948 19.819 12.012 ;
			RECT	19.955 11.948 19.987 12.012 ;
			RECT	20.123 11.948 20.155 12.012 ;
			RECT	20.291 11.948 20.323 12.012 ;
			RECT	20.459 11.948 20.491 12.012 ;
			RECT	20.627 11.948 20.659 12.012 ;
			RECT	20.795 11.948 20.827 12.012 ;
			RECT	20.963 11.948 20.995 12.012 ;
			RECT	21.131 11.948 21.163 12.012 ;
			RECT	21.299 11.948 21.331 12.012 ;
			RECT	21.467 11.948 21.499 12.012 ;
			RECT	21.635 11.948 21.667 12.012 ;
			RECT	21.803 11.948 21.835 12.012 ;
			RECT	21.971 11.948 22.003 12.012 ;
			RECT	22.139 11.948 22.171 12.012 ;
			RECT	22.307 11.948 22.339 12.012 ;
			RECT	22.475 11.948 22.507 12.012 ;
			RECT	22.643 11.948 22.675 12.012 ;
			RECT	22.811 11.948 22.843 12.012 ;
			RECT	22.979 11.948 23.011 12.012 ;
			RECT	23.147 11.948 23.179 12.012 ;
			RECT	23.315 11.948 23.347 12.012 ;
			RECT	23.483 11.948 23.515 12.012 ;
			RECT	23.651 11.948 23.683 12.012 ;
			RECT	23.819 11.948 23.851 12.012 ;
			RECT	23.987 11.948 24.019 12.012 ;
			RECT	24.155 11.948 24.187 12.012 ;
			RECT	24.323 11.948 24.355 12.012 ;
			RECT	24.491 11.948 24.523 12.012 ;
			RECT	24.659 11.948 24.691 12.012 ;
			RECT	24.827 11.948 24.859 12.012 ;
			RECT	24.995 11.948 25.027 12.012 ;
			RECT	25.163 11.948 25.195 12.012 ;
			RECT	25.331 11.948 25.363 12.012 ;
			RECT	25.499 11.948 25.531 12.012 ;
			RECT	25.667 11.948 25.699 12.012 ;
			RECT	25.835 11.948 25.867 12.012 ;
			RECT	26.003 11.948 26.035 12.012 ;
			RECT	26.171 11.948 26.203 12.012 ;
			RECT	26.339 11.948 26.371 12.012 ;
			RECT	26.507 11.948 26.539 12.012 ;
			RECT	26.675 11.948 26.707 12.012 ;
			RECT	26.843 11.948 26.875 12.012 ;
			RECT	27.011 11.948 27.043 12.012 ;
			RECT	27.179 11.948 27.211 12.012 ;
			RECT	27.347 11.948 27.379 12.012 ;
			RECT	27.515 11.948 27.547 12.012 ;
			RECT	27.683 11.948 27.715 12.012 ;
			RECT	27.851 11.948 27.883 12.012 ;
			RECT	28.019 11.948 28.051 12.012 ;
			RECT	28.187 11.948 28.219 12.012 ;
			RECT	28.355 11.948 28.387 12.012 ;
			RECT	28.523 11.948 28.555 12.012 ;
			RECT	28.691 11.948 28.723 12.012 ;
			RECT	28.859 11.948 28.891 12.012 ;
			RECT	29.027 11.948 29.059 12.012 ;
			RECT	29.195 11.948 29.227 12.012 ;
			RECT	29.363 11.948 29.395 12.012 ;
			RECT	29.531 11.948 29.563 12.012 ;
			RECT	29.699 11.948 29.731 12.012 ;
			RECT	29.867 11.948 29.899 12.012 ;
			RECT	30.035 11.948 30.067 12.012 ;
			RECT	30.203 11.948 30.235 12.012 ;
			RECT	30.371 11.948 30.403 12.012 ;
			RECT	30.539 11.948 30.571 12.012 ;
			RECT	30.707 11.948 30.739 12.012 ;
			RECT	30.875 11.948 30.907 12.012 ;
			RECT	31.043 11.948 31.075 12.012 ;
			RECT	31.211 11.948 31.243 12.012 ;
			RECT	31.379 11.948 31.411 12.012 ;
			RECT	31.547 11.948 31.579 12.012 ;
			RECT	31.715 11.948 31.747 12.012 ;
			RECT	31.883 11.948 31.915 12.012 ;
			RECT	32.051 11.948 32.083 12.012 ;
			RECT	32.219 11.948 32.251 12.012 ;
			RECT	32.387 11.948 32.419 12.012 ;
			RECT	32.555 11.948 32.587 12.012 ;
			RECT	32.723 11.948 32.755 12.012 ;
			RECT	32.891 11.948 32.923 12.012 ;
			RECT	33.059 11.948 33.091 12.012 ;
			RECT	33.227 11.948 33.259 12.012 ;
			RECT	33.395 11.948 33.427 12.012 ;
			RECT	33.563 11.948 33.595 12.012 ;
			RECT	33.731 11.948 33.763 12.012 ;
			RECT	33.899 11.948 33.931 12.012 ;
			RECT	34.067 11.948 34.099 12.012 ;
			RECT	34.235 11.948 34.267 12.012 ;
			RECT	34.403 11.948 34.435 12.012 ;
			RECT	34.571 11.948 34.603 12.012 ;
			RECT	34.739 11.948 34.771 12.012 ;
			RECT	34.907 11.948 34.939 12.012 ;
			RECT	35.075 11.948 35.107 12.012 ;
			RECT	35.243 11.948 35.275 12.012 ;
			RECT	35.411 11.948 35.443 12.012 ;
			RECT	35.579 11.948 35.611 12.012 ;
			RECT	35.747 11.948 35.779 12.012 ;
			RECT	35.915 11.948 35.947 12.012 ;
			RECT	36.083 11.948 36.115 12.012 ;
			RECT	36.251 11.948 36.283 12.012 ;
			RECT	36.419 11.948 36.451 12.012 ;
			RECT	36.587 11.948 36.619 12.012 ;
			RECT	36.755 11.948 36.787 12.012 ;
			RECT	36.923 11.948 36.955 12.012 ;
			RECT	37.091 11.948 37.123 12.012 ;
			RECT	37.259 11.948 37.291 12.012 ;
			RECT	37.427 11.948 37.459 12.012 ;
			RECT	37.595 11.948 37.627 12.012 ;
			RECT	37.763 11.948 37.795 12.012 ;
			RECT	37.931 11.948 37.963 12.012 ;
			RECT	38.099 11.948 38.131 12.012 ;
			RECT	38.267 11.948 38.299 12.012 ;
			RECT	38.435 11.948 38.467 12.012 ;
			RECT	38.603 11.948 38.635 12.012 ;
			RECT	38.771 11.948 38.803 12.012 ;
			RECT	38.939 11.948 38.971 12.012 ;
			RECT	39.107 11.948 39.139 12.012 ;
			RECT	39.275 11.948 39.307 12.012 ;
			RECT	39.443 11.948 39.475 12.012 ;
			RECT	39.611 11.948 39.643 12.012 ;
			RECT	39.779 11.948 39.811 12.012 ;
			RECT	39.947 11.948 39.979 12.012 ;
			RECT	40.115 11.948 40.147 12.012 ;
			RECT	40.283 11.948 40.315 12.012 ;
			RECT	40.451 11.948 40.483 12.012 ;
			RECT	40.619 11.948 40.651 12.012 ;
			RECT	40.787 11.948 40.819 12.012 ;
			RECT	40.955 11.948 40.987 12.012 ;
			RECT	41.123 11.948 41.155 12.012 ;
			RECT	41.291 11.948 41.323 12.012 ;
			RECT	41.459 11.948 41.491 12.012 ;
			RECT	41.627 11.948 41.659 12.012 ;
			RECT	41.795 11.948 41.827 12.012 ;
			RECT	41.963 11.948 41.995 12.012 ;
			RECT	42.131 11.948 42.163 12.012 ;
			RECT	42.299 11.948 42.331 12.012 ;
			RECT	42.467 11.948 42.499 12.012 ;
			RECT	42.635 11.948 42.667 12.012 ;
			RECT	42.803 11.948 42.835 12.012 ;
			RECT	42.971 11.948 43.003 12.012 ;
			RECT	43.139 11.948 43.171 12.012 ;
			RECT	43.307 11.948 43.339 12.012 ;
			RECT	43.475 11.948 43.507 12.012 ;
			RECT	43.643 11.948 43.675 12.012 ;
			RECT	43.811 11.948 43.843 12.012 ;
			RECT	43.979 11.948 44.011 12.012 ;
			RECT	44.147 11.948 44.179 12.012 ;
			RECT	44.315 11.948 44.347 12.012 ;
			RECT	44.483 11.948 44.515 12.012 ;
			RECT	44.651 11.948 44.683 12.012 ;
			RECT	44.819 11.948 44.851 12.012 ;
			RECT	44.987 11.948 45.019 12.012 ;
			RECT	45.155 11.948 45.187 12.012 ;
			RECT	45.323 11.948 45.355 12.012 ;
			RECT	45.491 11.948 45.523 12.012 ;
			RECT	45.659 11.948 45.691 12.012 ;
			RECT	45.827 11.948 45.859 12.012 ;
			RECT	45.995 11.948 46.027 12.012 ;
			RECT	46.163 11.948 46.195 12.012 ;
			RECT	46.331 11.948 46.363 12.012 ;
			RECT	46.499 11.948 46.531 12.012 ;
			RECT	46.667 11.948 46.699 12.012 ;
			RECT	46.835 11.948 46.867 12.012 ;
			RECT	47.003 11.948 47.035 12.012 ;
			RECT	47.171 11.948 47.203 12.012 ;
			RECT	47.339 11.948 47.371 12.012 ;
			RECT	47.507 11.948 47.539 12.012 ;
			RECT	47.675 11.948 47.707 12.012 ;
			RECT	47.843 11.948 47.875 12.012 ;
			RECT	48.011 11.948 48.043 12.012 ;
			RECT	48.179 11.948 48.211 12.012 ;
			RECT	48.347 11.948 48.379 12.012 ;
			RECT	48.515 11.948 48.547 12.012 ;
			RECT	48.683 11.948 48.715 12.012 ;
			RECT	48.851 11.948 48.883 12.012 ;
			RECT	49.019 11.948 49.051 12.012 ;
			RECT	49.187 11.948 49.219 12.012 ;
			RECT	49.318 11.964 49.35 11.996 ;
			RECT	49.439 11.964 49.471 11.996 ;
			RECT	49.569 11.948 49.601 12.012 ;
			RECT	51.881 11.948 51.913 12.012 ;
			RECT	53.132 11.948 53.196 12.012 ;
			RECT	53.812 11.948 53.844 12.012 ;
			RECT	54.251 11.948 54.283 12.012 ;
			RECT	55.562 11.948 55.626 12.012 ;
			RECT	58.603 11.948 58.635 12.012 ;
			RECT	58.733 11.964 58.765 11.996 ;
			RECT	58.854 11.964 58.886 11.996 ;
			RECT	58.985 11.948 59.017 12.012 ;
			RECT	59.153 11.948 59.185 12.012 ;
			RECT	59.321 11.948 59.353 12.012 ;
			RECT	59.489 11.948 59.521 12.012 ;
			RECT	59.657 11.948 59.689 12.012 ;
			RECT	59.825 11.948 59.857 12.012 ;
			RECT	59.993 11.948 60.025 12.012 ;
			RECT	60.161 11.948 60.193 12.012 ;
			RECT	60.329 11.948 60.361 12.012 ;
			RECT	60.497 11.948 60.529 12.012 ;
			RECT	60.665 11.948 60.697 12.012 ;
			RECT	60.833 11.948 60.865 12.012 ;
			RECT	61.001 11.948 61.033 12.012 ;
			RECT	61.169 11.948 61.201 12.012 ;
			RECT	61.337 11.948 61.369 12.012 ;
			RECT	61.505 11.948 61.537 12.012 ;
			RECT	61.673 11.948 61.705 12.012 ;
			RECT	61.841 11.948 61.873 12.012 ;
			RECT	62.009 11.948 62.041 12.012 ;
			RECT	62.177 11.948 62.209 12.012 ;
			RECT	62.345 11.948 62.377 12.012 ;
			RECT	62.513 11.948 62.545 12.012 ;
			RECT	62.681 11.948 62.713 12.012 ;
			RECT	62.849 11.948 62.881 12.012 ;
			RECT	63.017 11.948 63.049 12.012 ;
			RECT	63.185 11.948 63.217 12.012 ;
			RECT	63.353 11.948 63.385 12.012 ;
			RECT	63.521 11.948 63.553 12.012 ;
			RECT	63.689 11.948 63.721 12.012 ;
			RECT	63.857 11.948 63.889 12.012 ;
			RECT	64.025 11.948 64.057 12.012 ;
			RECT	64.193 11.948 64.225 12.012 ;
			RECT	64.361 11.948 64.393 12.012 ;
			RECT	64.529 11.948 64.561 12.012 ;
			RECT	64.697 11.948 64.729 12.012 ;
			RECT	64.865 11.948 64.897 12.012 ;
			RECT	65.033 11.948 65.065 12.012 ;
			RECT	65.201 11.948 65.233 12.012 ;
			RECT	65.369 11.948 65.401 12.012 ;
			RECT	65.537 11.948 65.569 12.012 ;
			RECT	65.705 11.948 65.737 12.012 ;
			RECT	65.873 11.948 65.905 12.012 ;
			RECT	66.041 11.948 66.073 12.012 ;
			RECT	66.209 11.948 66.241 12.012 ;
			RECT	66.377 11.948 66.409 12.012 ;
			RECT	66.545 11.948 66.577 12.012 ;
			RECT	66.713 11.948 66.745 12.012 ;
			RECT	66.881 11.948 66.913 12.012 ;
			RECT	67.049 11.948 67.081 12.012 ;
			RECT	67.217 11.948 67.249 12.012 ;
			RECT	67.385 11.948 67.417 12.012 ;
			RECT	67.553 11.948 67.585 12.012 ;
			RECT	67.721 11.948 67.753 12.012 ;
			RECT	67.889 11.948 67.921 12.012 ;
			RECT	68.057 11.948 68.089 12.012 ;
			RECT	68.225 11.948 68.257 12.012 ;
			RECT	68.393 11.948 68.425 12.012 ;
			RECT	68.561 11.948 68.593 12.012 ;
			RECT	68.729 11.948 68.761 12.012 ;
			RECT	68.897 11.948 68.929 12.012 ;
			RECT	69.065 11.948 69.097 12.012 ;
			RECT	69.233 11.948 69.265 12.012 ;
			RECT	69.401 11.948 69.433 12.012 ;
			RECT	69.569 11.948 69.601 12.012 ;
			RECT	69.737 11.948 69.769 12.012 ;
			RECT	69.905 11.948 69.937 12.012 ;
			RECT	70.073 11.948 70.105 12.012 ;
			RECT	70.241 11.948 70.273 12.012 ;
			RECT	70.409 11.948 70.441 12.012 ;
			RECT	70.577 11.948 70.609 12.012 ;
			RECT	70.745 11.948 70.777 12.012 ;
			RECT	70.913 11.948 70.945 12.012 ;
			RECT	71.081 11.948 71.113 12.012 ;
			RECT	71.249 11.948 71.281 12.012 ;
			RECT	71.417 11.948 71.449 12.012 ;
			RECT	71.585 11.948 71.617 12.012 ;
			RECT	71.753 11.948 71.785 12.012 ;
			RECT	71.921 11.948 71.953 12.012 ;
			RECT	72.089 11.948 72.121 12.012 ;
			RECT	72.257 11.948 72.289 12.012 ;
			RECT	72.425 11.948 72.457 12.012 ;
			RECT	72.593 11.948 72.625 12.012 ;
			RECT	72.761 11.948 72.793 12.012 ;
			RECT	72.929 11.948 72.961 12.012 ;
			RECT	73.097 11.948 73.129 12.012 ;
			RECT	73.265 11.948 73.297 12.012 ;
			RECT	73.433 11.948 73.465 12.012 ;
			RECT	73.601 11.948 73.633 12.012 ;
			RECT	73.769 11.948 73.801 12.012 ;
			RECT	73.937 11.948 73.969 12.012 ;
			RECT	74.105 11.948 74.137 12.012 ;
			RECT	74.273 11.948 74.305 12.012 ;
			RECT	74.441 11.948 74.473 12.012 ;
			RECT	74.609 11.948 74.641 12.012 ;
			RECT	74.777 11.948 74.809 12.012 ;
			RECT	74.945 11.948 74.977 12.012 ;
			RECT	75.113 11.948 75.145 12.012 ;
			RECT	75.281 11.948 75.313 12.012 ;
			RECT	75.449 11.948 75.481 12.012 ;
			RECT	75.617 11.948 75.649 12.012 ;
			RECT	75.785 11.948 75.817 12.012 ;
			RECT	75.953 11.948 75.985 12.012 ;
			RECT	76.121 11.948 76.153 12.012 ;
			RECT	76.289 11.948 76.321 12.012 ;
			RECT	76.457 11.948 76.489 12.012 ;
			RECT	76.625 11.948 76.657 12.012 ;
			RECT	76.793 11.948 76.825 12.012 ;
			RECT	76.961 11.948 76.993 12.012 ;
			RECT	77.129 11.948 77.161 12.012 ;
			RECT	77.297 11.948 77.329 12.012 ;
			RECT	77.465 11.948 77.497 12.012 ;
			RECT	77.633 11.948 77.665 12.012 ;
			RECT	77.801 11.948 77.833 12.012 ;
			RECT	77.969 11.948 78.001 12.012 ;
			RECT	78.137 11.948 78.169 12.012 ;
			RECT	78.305 11.948 78.337 12.012 ;
			RECT	78.473 11.948 78.505 12.012 ;
			RECT	78.641 11.948 78.673 12.012 ;
			RECT	78.809 11.948 78.841 12.012 ;
			RECT	78.977 11.948 79.009 12.012 ;
			RECT	79.145 11.948 79.177 12.012 ;
			RECT	79.313 11.948 79.345 12.012 ;
			RECT	79.481 11.948 79.513 12.012 ;
			RECT	79.649 11.948 79.681 12.012 ;
			RECT	79.817 11.948 79.849 12.012 ;
			RECT	79.985 11.948 80.017 12.012 ;
			RECT	80.153 11.948 80.185 12.012 ;
			RECT	80.321 11.948 80.353 12.012 ;
			RECT	80.489 11.948 80.521 12.012 ;
			RECT	80.657 11.948 80.689 12.012 ;
			RECT	80.825 11.948 80.857 12.012 ;
			RECT	80.993 11.948 81.025 12.012 ;
			RECT	81.161 11.948 81.193 12.012 ;
			RECT	81.329 11.948 81.361 12.012 ;
			RECT	81.497 11.948 81.529 12.012 ;
			RECT	81.665 11.948 81.697 12.012 ;
			RECT	81.833 11.948 81.865 12.012 ;
			RECT	82.001 11.948 82.033 12.012 ;
			RECT	82.169 11.948 82.201 12.012 ;
			RECT	82.337 11.948 82.369 12.012 ;
			RECT	82.505 11.948 82.537 12.012 ;
			RECT	82.673 11.948 82.705 12.012 ;
			RECT	82.841 11.948 82.873 12.012 ;
			RECT	83.009 11.948 83.041 12.012 ;
			RECT	83.177 11.948 83.209 12.012 ;
			RECT	83.345 11.948 83.377 12.012 ;
			RECT	83.513 11.948 83.545 12.012 ;
			RECT	83.681 11.948 83.713 12.012 ;
			RECT	83.849 11.948 83.881 12.012 ;
			RECT	84.017 11.948 84.049 12.012 ;
			RECT	84.185 11.948 84.217 12.012 ;
			RECT	84.353 11.948 84.385 12.012 ;
			RECT	84.521 11.948 84.553 12.012 ;
			RECT	84.689 11.948 84.721 12.012 ;
			RECT	84.857 11.948 84.889 12.012 ;
			RECT	85.025 11.948 85.057 12.012 ;
			RECT	85.193 11.948 85.225 12.012 ;
			RECT	85.361 11.948 85.393 12.012 ;
			RECT	85.529 11.948 85.561 12.012 ;
			RECT	85.697 11.948 85.729 12.012 ;
			RECT	85.865 11.948 85.897 12.012 ;
			RECT	86.033 11.948 86.065 12.012 ;
			RECT	86.201 11.948 86.233 12.012 ;
			RECT	86.369 11.948 86.401 12.012 ;
			RECT	86.537 11.948 86.569 12.012 ;
			RECT	86.705 11.948 86.737 12.012 ;
			RECT	86.873 11.948 86.905 12.012 ;
			RECT	87.041 11.948 87.073 12.012 ;
			RECT	87.209 11.948 87.241 12.012 ;
			RECT	87.377 11.948 87.409 12.012 ;
			RECT	87.545 11.948 87.577 12.012 ;
			RECT	87.713 11.948 87.745 12.012 ;
			RECT	87.881 11.948 87.913 12.012 ;
			RECT	88.049 11.948 88.081 12.012 ;
			RECT	88.217 11.948 88.249 12.012 ;
			RECT	88.385 11.948 88.417 12.012 ;
			RECT	88.553 11.948 88.585 12.012 ;
			RECT	88.721 11.948 88.753 12.012 ;
			RECT	88.889 11.948 88.921 12.012 ;
			RECT	89.057 11.948 89.089 12.012 ;
			RECT	89.225 11.948 89.257 12.012 ;
			RECT	89.393 11.948 89.425 12.012 ;
			RECT	89.561 11.948 89.593 12.012 ;
			RECT	89.729 11.948 89.761 12.012 ;
			RECT	89.897 11.948 89.929 12.012 ;
			RECT	90.065 11.948 90.097 12.012 ;
			RECT	90.233 11.948 90.265 12.012 ;
			RECT	90.401 11.948 90.433 12.012 ;
			RECT	90.569 11.948 90.601 12.012 ;
			RECT	90.737 11.948 90.769 12.012 ;
			RECT	90.905 11.948 90.937 12.012 ;
			RECT	91.073 11.948 91.105 12.012 ;
			RECT	91.241 11.948 91.273 12.012 ;
			RECT	91.409 11.948 91.441 12.012 ;
			RECT	91.577 11.948 91.609 12.012 ;
			RECT	91.745 11.948 91.777 12.012 ;
			RECT	91.913 11.948 91.945 12.012 ;
			RECT	92.081 11.948 92.113 12.012 ;
			RECT	92.249 11.948 92.281 12.012 ;
			RECT	92.417 11.948 92.449 12.012 ;
			RECT	92.585 11.948 92.617 12.012 ;
			RECT	92.753 11.948 92.785 12.012 ;
			RECT	92.921 11.948 92.953 12.012 ;
			RECT	93.089 11.948 93.121 12.012 ;
			RECT	93.257 11.948 93.289 12.012 ;
			RECT	93.425 11.948 93.457 12.012 ;
			RECT	93.593 11.948 93.625 12.012 ;
			RECT	93.761 11.948 93.793 12.012 ;
			RECT	93.929 11.948 93.961 12.012 ;
			RECT	94.097 11.948 94.129 12.012 ;
			RECT	94.265 11.948 94.297 12.012 ;
			RECT	94.433 11.948 94.465 12.012 ;
			RECT	94.601 11.948 94.633 12.012 ;
			RECT	94.769 11.948 94.801 12.012 ;
			RECT	94.937 11.948 94.969 12.012 ;
			RECT	95.105 11.948 95.137 12.012 ;
			RECT	95.273 11.948 95.305 12.012 ;
			RECT	95.441 11.948 95.473 12.012 ;
			RECT	95.609 11.948 95.641 12.012 ;
			RECT	95.777 11.948 95.809 12.012 ;
			RECT	95.945 11.948 95.977 12.012 ;
			RECT	96.113 11.948 96.145 12.012 ;
			RECT	96.281 11.948 96.313 12.012 ;
			RECT	96.449 11.948 96.481 12.012 ;
			RECT	96.617 11.948 96.649 12.012 ;
			RECT	96.785 11.948 96.817 12.012 ;
			RECT	96.953 11.948 96.985 12.012 ;
			RECT	97.121 11.948 97.153 12.012 ;
			RECT	97.289 11.948 97.321 12.012 ;
			RECT	97.457 11.948 97.489 12.012 ;
			RECT	97.625 11.948 97.657 12.012 ;
			RECT	97.793 11.948 97.825 12.012 ;
			RECT	97.961 11.948 97.993 12.012 ;
			RECT	98.129 11.948 98.161 12.012 ;
			RECT	98.297 11.948 98.329 12.012 ;
			RECT	98.465 11.948 98.497 12.012 ;
			RECT	98.633 11.948 98.665 12.012 ;
			RECT	98.801 11.948 98.833 12.012 ;
			RECT	98.969 11.948 99.001 12.012 ;
			RECT	99.137 11.948 99.169 12.012 ;
			RECT	99.305 11.948 99.337 12.012 ;
			RECT	99.473 11.948 99.505 12.012 ;
			RECT	99.641 11.948 99.673 12.012 ;
			RECT	99.809 11.948 99.841 12.012 ;
			RECT	99.977 11.948 100.009 12.012 ;
			RECT	100.145 11.948 100.177 12.012 ;
			RECT	100.313 11.948 100.345 12.012 ;
			RECT	100.481 11.948 100.513 12.012 ;
			RECT	100.649 11.948 100.681 12.012 ;
			RECT	100.817 11.948 100.849 12.012 ;
			RECT	100.985 11.948 101.017 12.012 ;
			RECT	101.153 11.948 101.185 12.012 ;
			RECT	101.321 11.948 101.353 12.012 ;
			RECT	101.489 11.948 101.521 12.012 ;
			RECT	101.657 11.948 101.689 12.012 ;
			RECT	101.825 11.948 101.857 12.012 ;
			RECT	101.993 11.948 102.025 12.012 ;
			RECT	102.123 11.964 102.155 11.996 ;
			RECT	102.245 11.969 102.277 12.001 ;
			RECT	102.375 11.948 102.407 12.012 ;
			RECT	103.795 11.948 103.827 12.012 ;
			RECT	103.925 11.969 103.957 12.001 ;
			RECT	104.047 11.964 104.079 11.996 ;
			RECT	104.177 11.948 104.209 12.012 ;
			RECT	104.345 11.948 104.377 12.012 ;
			RECT	104.513 11.948 104.545 12.012 ;
			RECT	104.681 11.948 104.713 12.012 ;
			RECT	104.849 11.948 104.881 12.012 ;
			RECT	105.017 11.948 105.049 12.012 ;
			RECT	105.185 11.948 105.217 12.012 ;
			RECT	105.353 11.948 105.385 12.012 ;
			RECT	105.521 11.948 105.553 12.012 ;
			RECT	105.689 11.948 105.721 12.012 ;
			RECT	105.857 11.948 105.889 12.012 ;
			RECT	106.025 11.948 106.057 12.012 ;
			RECT	106.193 11.948 106.225 12.012 ;
			RECT	106.361 11.948 106.393 12.012 ;
			RECT	106.529 11.948 106.561 12.012 ;
			RECT	106.697 11.948 106.729 12.012 ;
			RECT	106.865 11.948 106.897 12.012 ;
			RECT	107.033 11.948 107.065 12.012 ;
			RECT	107.201 11.948 107.233 12.012 ;
			RECT	107.369 11.948 107.401 12.012 ;
			RECT	107.537 11.948 107.569 12.012 ;
			RECT	107.705 11.948 107.737 12.012 ;
			RECT	107.873 11.948 107.905 12.012 ;
			RECT	108.041 11.948 108.073 12.012 ;
			RECT	108.209 11.948 108.241 12.012 ;
			RECT	108.377 11.948 108.409 12.012 ;
			RECT	108.545 11.948 108.577 12.012 ;
			RECT	108.713 11.948 108.745 12.012 ;
			RECT	108.881 11.948 108.913 12.012 ;
			RECT	109.049 11.948 109.081 12.012 ;
			RECT	109.217 11.948 109.249 12.012 ;
			RECT	109.385 11.948 109.417 12.012 ;
			RECT	109.553 11.948 109.585 12.012 ;
			RECT	109.721 11.948 109.753 12.012 ;
			RECT	109.889 11.948 109.921 12.012 ;
			RECT	110.057 11.948 110.089 12.012 ;
			RECT	110.225 11.948 110.257 12.012 ;
			RECT	110.393 11.948 110.425 12.012 ;
			RECT	110.561 11.948 110.593 12.012 ;
			RECT	110.729 11.948 110.761 12.012 ;
			RECT	110.897 11.948 110.929 12.012 ;
			RECT	111.065 11.948 111.097 12.012 ;
			RECT	111.233 11.948 111.265 12.012 ;
			RECT	111.401 11.948 111.433 12.012 ;
			RECT	111.569 11.948 111.601 12.012 ;
			RECT	111.737 11.948 111.769 12.012 ;
			RECT	111.905 11.948 111.937 12.012 ;
			RECT	112.073 11.948 112.105 12.012 ;
			RECT	112.241 11.948 112.273 12.012 ;
			RECT	112.409 11.948 112.441 12.012 ;
			RECT	112.577 11.948 112.609 12.012 ;
			RECT	112.745 11.948 112.777 12.012 ;
			RECT	112.913 11.948 112.945 12.012 ;
			RECT	113.081 11.948 113.113 12.012 ;
			RECT	113.249 11.948 113.281 12.012 ;
			RECT	113.417 11.948 113.449 12.012 ;
			RECT	113.585 11.948 113.617 12.012 ;
			RECT	113.753 11.948 113.785 12.012 ;
			RECT	113.921 11.948 113.953 12.012 ;
			RECT	114.089 11.948 114.121 12.012 ;
			RECT	114.257 11.948 114.289 12.012 ;
			RECT	114.425 11.948 114.457 12.012 ;
			RECT	114.593 11.948 114.625 12.012 ;
			RECT	114.761 11.948 114.793 12.012 ;
			RECT	114.929 11.948 114.961 12.012 ;
			RECT	115.097 11.948 115.129 12.012 ;
			RECT	115.265 11.948 115.297 12.012 ;
			RECT	115.433 11.948 115.465 12.012 ;
			RECT	115.601 11.948 115.633 12.012 ;
			RECT	115.769 11.948 115.801 12.012 ;
			RECT	115.937 11.948 115.969 12.012 ;
			RECT	116.105 11.948 116.137 12.012 ;
			RECT	116.273 11.948 116.305 12.012 ;
			RECT	116.441 11.948 116.473 12.012 ;
			RECT	116.609 11.948 116.641 12.012 ;
			RECT	116.777 11.948 116.809 12.012 ;
			RECT	116.945 11.948 116.977 12.012 ;
			RECT	117.113 11.948 117.145 12.012 ;
			RECT	117.281 11.948 117.313 12.012 ;
			RECT	117.449 11.948 117.481 12.012 ;
			RECT	117.617 11.948 117.649 12.012 ;
			RECT	117.785 11.948 117.817 12.012 ;
			RECT	117.953 11.948 117.985 12.012 ;
			RECT	118.121 11.948 118.153 12.012 ;
			RECT	118.289 11.948 118.321 12.012 ;
			RECT	118.457 11.948 118.489 12.012 ;
			RECT	118.625 11.948 118.657 12.012 ;
			RECT	118.793 11.948 118.825 12.012 ;
			RECT	118.961 11.948 118.993 12.012 ;
			RECT	119.129 11.948 119.161 12.012 ;
			RECT	119.297 11.948 119.329 12.012 ;
			RECT	119.465 11.948 119.497 12.012 ;
			RECT	119.633 11.948 119.665 12.012 ;
			RECT	119.801 11.948 119.833 12.012 ;
			RECT	119.969 11.948 120.001 12.012 ;
			RECT	120.137 11.948 120.169 12.012 ;
			RECT	120.305 11.948 120.337 12.012 ;
			RECT	120.473 11.948 120.505 12.012 ;
			RECT	120.641 11.948 120.673 12.012 ;
			RECT	120.809 11.948 120.841 12.012 ;
			RECT	120.977 11.948 121.009 12.012 ;
			RECT	121.145 11.948 121.177 12.012 ;
			RECT	121.313 11.948 121.345 12.012 ;
			RECT	121.481 11.948 121.513 12.012 ;
			RECT	121.649 11.948 121.681 12.012 ;
			RECT	121.817 11.948 121.849 12.012 ;
			RECT	121.985 11.948 122.017 12.012 ;
			RECT	122.153 11.948 122.185 12.012 ;
			RECT	122.321 11.948 122.353 12.012 ;
			RECT	122.489 11.948 122.521 12.012 ;
			RECT	122.657 11.948 122.689 12.012 ;
			RECT	122.825 11.948 122.857 12.012 ;
			RECT	122.993 11.948 123.025 12.012 ;
			RECT	123.161 11.948 123.193 12.012 ;
			RECT	123.329 11.948 123.361 12.012 ;
			RECT	123.497 11.948 123.529 12.012 ;
			RECT	123.665 11.948 123.697 12.012 ;
			RECT	123.833 11.948 123.865 12.012 ;
			RECT	124.001 11.948 124.033 12.012 ;
			RECT	124.169 11.948 124.201 12.012 ;
			RECT	124.337 11.948 124.369 12.012 ;
			RECT	124.505 11.948 124.537 12.012 ;
			RECT	124.673 11.948 124.705 12.012 ;
			RECT	124.841 11.948 124.873 12.012 ;
			RECT	125.009 11.948 125.041 12.012 ;
			RECT	125.177 11.948 125.209 12.012 ;
			RECT	125.345 11.948 125.377 12.012 ;
			RECT	125.513 11.948 125.545 12.012 ;
			RECT	125.681 11.948 125.713 12.012 ;
			RECT	125.849 11.948 125.881 12.012 ;
			RECT	126.017 11.948 126.049 12.012 ;
			RECT	126.185 11.948 126.217 12.012 ;
			RECT	126.353 11.948 126.385 12.012 ;
			RECT	126.521 11.948 126.553 12.012 ;
			RECT	126.689 11.948 126.721 12.012 ;
			RECT	126.857 11.948 126.889 12.012 ;
			RECT	127.025 11.948 127.057 12.012 ;
			RECT	127.193 11.948 127.225 12.012 ;
			RECT	127.361 11.948 127.393 12.012 ;
			RECT	127.529 11.948 127.561 12.012 ;
			RECT	127.697 11.948 127.729 12.012 ;
			RECT	127.865 11.948 127.897 12.012 ;
			RECT	128.033 11.948 128.065 12.012 ;
			RECT	128.201 11.948 128.233 12.012 ;
			RECT	128.369 11.948 128.401 12.012 ;
			RECT	128.537 11.948 128.569 12.012 ;
			RECT	128.705 11.948 128.737 12.012 ;
			RECT	128.873 11.948 128.905 12.012 ;
			RECT	129.041 11.948 129.073 12.012 ;
			RECT	129.209 11.948 129.241 12.012 ;
			RECT	129.377 11.948 129.409 12.012 ;
			RECT	129.545 11.948 129.577 12.012 ;
			RECT	129.713 11.948 129.745 12.012 ;
			RECT	129.881 11.948 129.913 12.012 ;
			RECT	130.049 11.948 130.081 12.012 ;
			RECT	130.217 11.948 130.249 12.012 ;
			RECT	130.385 11.948 130.417 12.012 ;
			RECT	130.553 11.948 130.585 12.012 ;
			RECT	130.721 11.948 130.753 12.012 ;
			RECT	130.889 11.948 130.921 12.012 ;
			RECT	131.057 11.948 131.089 12.012 ;
			RECT	131.225 11.948 131.257 12.012 ;
			RECT	131.393 11.948 131.425 12.012 ;
			RECT	131.561 11.948 131.593 12.012 ;
			RECT	131.729 11.948 131.761 12.012 ;
			RECT	131.897 11.948 131.929 12.012 ;
			RECT	132.065 11.948 132.097 12.012 ;
			RECT	132.233 11.948 132.265 12.012 ;
			RECT	132.401 11.948 132.433 12.012 ;
			RECT	132.569 11.948 132.601 12.012 ;
			RECT	132.737 11.948 132.769 12.012 ;
			RECT	132.905 11.948 132.937 12.012 ;
			RECT	133.073 11.948 133.105 12.012 ;
			RECT	133.241 11.948 133.273 12.012 ;
			RECT	133.409 11.948 133.441 12.012 ;
			RECT	133.577 11.948 133.609 12.012 ;
			RECT	133.745 11.948 133.777 12.012 ;
			RECT	133.913 11.948 133.945 12.012 ;
			RECT	134.081 11.948 134.113 12.012 ;
			RECT	134.249 11.948 134.281 12.012 ;
			RECT	134.417 11.948 134.449 12.012 ;
			RECT	134.585 11.948 134.617 12.012 ;
			RECT	134.753 11.948 134.785 12.012 ;
			RECT	134.921 11.948 134.953 12.012 ;
			RECT	135.089 11.948 135.121 12.012 ;
			RECT	135.257 11.948 135.289 12.012 ;
			RECT	135.425 11.948 135.457 12.012 ;
			RECT	135.593 11.948 135.625 12.012 ;
			RECT	135.761 11.948 135.793 12.012 ;
			RECT	135.929 11.948 135.961 12.012 ;
			RECT	136.097 11.948 136.129 12.012 ;
			RECT	136.265 11.948 136.297 12.012 ;
			RECT	136.433 11.948 136.465 12.012 ;
			RECT	136.601 11.948 136.633 12.012 ;
			RECT	136.769 11.948 136.801 12.012 ;
			RECT	136.937 11.948 136.969 12.012 ;
			RECT	137.105 11.948 137.137 12.012 ;
			RECT	137.273 11.948 137.305 12.012 ;
			RECT	137.441 11.948 137.473 12.012 ;
			RECT	137.609 11.948 137.641 12.012 ;
			RECT	137.777 11.948 137.809 12.012 ;
			RECT	137.945 11.948 137.977 12.012 ;
			RECT	138.113 11.948 138.145 12.012 ;
			RECT	138.281 11.948 138.313 12.012 ;
			RECT	138.449 11.948 138.481 12.012 ;
			RECT	138.617 11.948 138.649 12.012 ;
			RECT	138.785 11.948 138.817 12.012 ;
			RECT	138.953 11.948 138.985 12.012 ;
			RECT	139.121 11.948 139.153 12.012 ;
			RECT	139.289 11.948 139.321 12.012 ;
			RECT	139.457 11.948 139.489 12.012 ;
			RECT	139.625 11.948 139.657 12.012 ;
			RECT	139.793 11.948 139.825 12.012 ;
			RECT	139.961 11.948 139.993 12.012 ;
			RECT	140.129 11.948 140.161 12.012 ;
			RECT	140.297 11.948 140.329 12.012 ;
			RECT	140.465 11.948 140.497 12.012 ;
			RECT	140.633 11.948 140.665 12.012 ;
			RECT	140.801 11.948 140.833 12.012 ;
			RECT	140.969 11.948 141.001 12.012 ;
			RECT	141.137 11.948 141.169 12.012 ;
			RECT	141.305 11.948 141.337 12.012 ;
			RECT	141.473 11.948 141.505 12.012 ;
			RECT	141.641 11.948 141.673 12.012 ;
			RECT	141.809 11.948 141.841 12.012 ;
			RECT	141.977 11.948 142.009 12.012 ;
			RECT	142.145 11.948 142.177 12.012 ;
			RECT	142.313 11.948 142.345 12.012 ;
			RECT	142.481 11.948 142.513 12.012 ;
			RECT	142.649 11.948 142.681 12.012 ;
			RECT	142.817 11.948 142.849 12.012 ;
			RECT	142.985 11.948 143.017 12.012 ;
			RECT	143.153 11.948 143.185 12.012 ;
			RECT	143.321 11.948 143.353 12.012 ;
			RECT	143.489 11.948 143.521 12.012 ;
			RECT	143.657 11.948 143.689 12.012 ;
			RECT	143.825 11.948 143.857 12.012 ;
			RECT	143.993 11.948 144.025 12.012 ;
			RECT	144.161 11.948 144.193 12.012 ;
			RECT	144.329 11.948 144.361 12.012 ;
			RECT	144.497 11.948 144.529 12.012 ;
			RECT	144.665 11.948 144.697 12.012 ;
			RECT	144.833 11.948 144.865 12.012 ;
			RECT	145.001 11.948 145.033 12.012 ;
			RECT	145.169 11.948 145.201 12.012 ;
			RECT	145.337 11.948 145.369 12.012 ;
			RECT	145.505 11.948 145.537 12.012 ;
			RECT	145.673 11.948 145.705 12.012 ;
			RECT	145.841 11.948 145.873 12.012 ;
			RECT	146.009 11.948 146.041 12.012 ;
			RECT	146.177 11.948 146.209 12.012 ;
			RECT	146.345 11.948 146.377 12.012 ;
			RECT	146.513 11.948 146.545 12.012 ;
			RECT	146.681 11.948 146.713 12.012 ;
			RECT	146.849 11.948 146.881 12.012 ;
			RECT	147.017 11.948 147.049 12.012 ;
			RECT	147.185 11.948 147.217 12.012 ;
			RECT	147.316 11.964 147.348 11.996 ;
			RECT	147.437 11.964 147.469 11.996 ;
			RECT	147.567 11.948 147.599 12.012 ;
			RECT	149.879 11.948 149.911 12.012 ;
			RECT	151.13 11.948 151.194 12.012 ;
			RECT	151.81 11.948 151.842 12.012 ;
			RECT	152.249 11.948 152.281 12.012 ;
			RECT	153.56 11.948 153.624 12.012 ;
			RECT	156.601 11.948 156.633 12.012 ;
			RECT	156.731 11.964 156.763 11.996 ;
			RECT	156.852 11.964 156.884 11.996 ;
			RECT	156.983 11.948 157.015 12.012 ;
			RECT	157.151 11.948 157.183 12.012 ;
			RECT	157.319 11.948 157.351 12.012 ;
			RECT	157.487 11.948 157.519 12.012 ;
			RECT	157.655 11.948 157.687 12.012 ;
			RECT	157.823 11.948 157.855 12.012 ;
			RECT	157.991 11.948 158.023 12.012 ;
			RECT	158.159 11.948 158.191 12.012 ;
			RECT	158.327 11.948 158.359 12.012 ;
			RECT	158.495 11.948 158.527 12.012 ;
			RECT	158.663 11.948 158.695 12.012 ;
			RECT	158.831 11.948 158.863 12.012 ;
			RECT	158.999 11.948 159.031 12.012 ;
			RECT	159.167 11.948 159.199 12.012 ;
			RECT	159.335 11.948 159.367 12.012 ;
			RECT	159.503 11.948 159.535 12.012 ;
			RECT	159.671 11.948 159.703 12.012 ;
			RECT	159.839 11.948 159.871 12.012 ;
			RECT	160.007 11.948 160.039 12.012 ;
			RECT	160.175 11.948 160.207 12.012 ;
			RECT	160.343 11.948 160.375 12.012 ;
			RECT	160.511 11.948 160.543 12.012 ;
			RECT	160.679 11.948 160.711 12.012 ;
			RECT	160.847 11.948 160.879 12.012 ;
			RECT	161.015 11.948 161.047 12.012 ;
			RECT	161.183 11.948 161.215 12.012 ;
			RECT	161.351 11.948 161.383 12.012 ;
			RECT	161.519 11.948 161.551 12.012 ;
			RECT	161.687 11.948 161.719 12.012 ;
			RECT	161.855 11.948 161.887 12.012 ;
			RECT	162.023 11.948 162.055 12.012 ;
			RECT	162.191 11.948 162.223 12.012 ;
			RECT	162.359 11.948 162.391 12.012 ;
			RECT	162.527 11.948 162.559 12.012 ;
			RECT	162.695 11.948 162.727 12.012 ;
			RECT	162.863 11.948 162.895 12.012 ;
			RECT	163.031 11.948 163.063 12.012 ;
			RECT	163.199 11.948 163.231 12.012 ;
			RECT	163.367 11.948 163.399 12.012 ;
			RECT	163.535 11.948 163.567 12.012 ;
			RECT	163.703 11.948 163.735 12.012 ;
			RECT	163.871 11.948 163.903 12.012 ;
			RECT	164.039 11.948 164.071 12.012 ;
			RECT	164.207 11.948 164.239 12.012 ;
			RECT	164.375 11.948 164.407 12.012 ;
			RECT	164.543 11.948 164.575 12.012 ;
			RECT	164.711 11.948 164.743 12.012 ;
			RECT	164.879 11.948 164.911 12.012 ;
			RECT	165.047 11.948 165.079 12.012 ;
			RECT	165.215 11.948 165.247 12.012 ;
			RECT	165.383 11.948 165.415 12.012 ;
			RECT	165.551 11.948 165.583 12.012 ;
			RECT	165.719 11.948 165.751 12.012 ;
			RECT	165.887 11.948 165.919 12.012 ;
			RECT	166.055 11.948 166.087 12.012 ;
			RECT	166.223 11.948 166.255 12.012 ;
			RECT	166.391 11.948 166.423 12.012 ;
			RECT	166.559 11.948 166.591 12.012 ;
			RECT	166.727 11.948 166.759 12.012 ;
			RECT	166.895 11.948 166.927 12.012 ;
			RECT	167.063 11.948 167.095 12.012 ;
			RECT	167.231 11.948 167.263 12.012 ;
			RECT	167.399 11.948 167.431 12.012 ;
			RECT	167.567 11.948 167.599 12.012 ;
			RECT	167.735 11.948 167.767 12.012 ;
			RECT	167.903 11.948 167.935 12.012 ;
			RECT	168.071 11.948 168.103 12.012 ;
			RECT	168.239 11.948 168.271 12.012 ;
			RECT	168.407 11.948 168.439 12.012 ;
			RECT	168.575 11.948 168.607 12.012 ;
			RECT	168.743 11.948 168.775 12.012 ;
			RECT	168.911 11.948 168.943 12.012 ;
			RECT	169.079 11.948 169.111 12.012 ;
			RECT	169.247 11.948 169.279 12.012 ;
			RECT	169.415 11.948 169.447 12.012 ;
			RECT	169.583 11.948 169.615 12.012 ;
			RECT	169.751 11.948 169.783 12.012 ;
			RECT	169.919 11.948 169.951 12.012 ;
			RECT	170.087 11.948 170.119 12.012 ;
			RECT	170.255 11.948 170.287 12.012 ;
			RECT	170.423 11.948 170.455 12.012 ;
			RECT	170.591 11.948 170.623 12.012 ;
			RECT	170.759 11.948 170.791 12.012 ;
			RECT	170.927 11.948 170.959 12.012 ;
			RECT	171.095 11.948 171.127 12.012 ;
			RECT	171.263 11.948 171.295 12.012 ;
			RECT	171.431 11.948 171.463 12.012 ;
			RECT	171.599 11.948 171.631 12.012 ;
			RECT	171.767 11.948 171.799 12.012 ;
			RECT	171.935 11.948 171.967 12.012 ;
			RECT	172.103 11.948 172.135 12.012 ;
			RECT	172.271 11.948 172.303 12.012 ;
			RECT	172.439 11.948 172.471 12.012 ;
			RECT	172.607 11.948 172.639 12.012 ;
			RECT	172.775 11.948 172.807 12.012 ;
			RECT	172.943 11.948 172.975 12.012 ;
			RECT	173.111 11.948 173.143 12.012 ;
			RECT	173.279 11.948 173.311 12.012 ;
			RECT	173.447 11.948 173.479 12.012 ;
			RECT	173.615 11.948 173.647 12.012 ;
			RECT	173.783 11.948 173.815 12.012 ;
			RECT	173.951 11.948 173.983 12.012 ;
			RECT	174.119 11.948 174.151 12.012 ;
			RECT	174.287 11.948 174.319 12.012 ;
			RECT	174.455 11.948 174.487 12.012 ;
			RECT	174.623 11.948 174.655 12.012 ;
			RECT	174.791 11.948 174.823 12.012 ;
			RECT	174.959 11.948 174.991 12.012 ;
			RECT	175.127 11.948 175.159 12.012 ;
			RECT	175.295 11.948 175.327 12.012 ;
			RECT	175.463 11.948 175.495 12.012 ;
			RECT	175.631 11.948 175.663 12.012 ;
			RECT	175.799 11.948 175.831 12.012 ;
			RECT	175.967 11.948 175.999 12.012 ;
			RECT	176.135 11.948 176.167 12.012 ;
			RECT	176.303 11.948 176.335 12.012 ;
			RECT	176.471 11.948 176.503 12.012 ;
			RECT	176.639 11.948 176.671 12.012 ;
			RECT	176.807 11.948 176.839 12.012 ;
			RECT	176.975 11.948 177.007 12.012 ;
			RECT	177.143 11.948 177.175 12.012 ;
			RECT	177.311 11.948 177.343 12.012 ;
			RECT	177.479 11.948 177.511 12.012 ;
			RECT	177.647 11.948 177.679 12.012 ;
			RECT	177.815 11.948 177.847 12.012 ;
			RECT	177.983 11.948 178.015 12.012 ;
			RECT	178.151 11.948 178.183 12.012 ;
			RECT	178.319 11.948 178.351 12.012 ;
			RECT	178.487 11.948 178.519 12.012 ;
			RECT	178.655 11.948 178.687 12.012 ;
			RECT	178.823 11.948 178.855 12.012 ;
			RECT	178.991 11.948 179.023 12.012 ;
			RECT	179.159 11.948 179.191 12.012 ;
			RECT	179.327 11.948 179.359 12.012 ;
			RECT	179.495 11.948 179.527 12.012 ;
			RECT	179.663 11.948 179.695 12.012 ;
			RECT	179.831 11.948 179.863 12.012 ;
			RECT	179.999 11.948 180.031 12.012 ;
			RECT	180.167 11.948 180.199 12.012 ;
			RECT	180.335 11.948 180.367 12.012 ;
			RECT	180.503 11.948 180.535 12.012 ;
			RECT	180.671 11.948 180.703 12.012 ;
			RECT	180.839 11.948 180.871 12.012 ;
			RECT	181.007 11.948 181.039 12.012 ;
			RECT	181.175 11.948 181.207 12.012 ;
			RECT	181.343 11.948 181.375 12.012 ;
			RECT	181.511 11.948 181.543 12.012 ;
			RECT	181.679 11.948 181.711 12.012 ;
			RECT	181.847 11.948 181.879 12.012 ;
			RECT	182.015 11.948 182.047 12.012 ;
			RECT	182.183 11.948 182.215 12.012 ;
			RECT	182.351 11.948 182.383 12.012 ;
			RECT	182.519 11.948 182.551 12.012 ;
			RECT	182.687 11.948 182.719 12.012 ;
			RECT	182.855 11.948 182.887 12.012 ;
			RECT	183.023 11.948 183.055 12.012 ;
			RECT	183.191 11.948 183.223 12.012 ;
			RECT	183.359 11.948 183.391 12.012 ;
			RECT	183.527 11.948 183.559 12.012 ;
			RECT	183.695 11.948 183.727 12.012 ;
			RECT	183.863 11.948 183.895 12.012 ;
			RECT	184.031 11.948 184.063 12.012 ;
			RECT	184.199 11.948 184.231 12.012 ;
			RECT	184.367 11.948 184.399 12.012 ;
			RECT	184.535 11.948 184.567 12.012 ;
			RECT	184.703 11.948 184.735 12.012 ;
			RECT	184.871 11.948 184.903 12.012 ;
			RECT	185.039 11.948 185.071 12.012 ;
			RECT	185.207 11.948 185.239 12.012 ;
			RECT	185.375 11.948 185.407 12.012 ;
			RECT	185.543 11.948 185.575 12.012 ;
			RECT	185.711 11.948 185.743 12.012 ;
			RECT	185.879 11.948 185.911 12.012 ;
			RECT	186.047 11.948 186.079 12.012 ;
			RECT	186.215 11.948 186.247 12.012 ;
			RECT	186.383 11.948 186.415 12.012 ;
			RECT	186.551 11.948 186.583 12.012 ;
			RECT	186.719 11.948 186.751 12.012 ;
			RECT	186.887 11.948 186.919 12.012 ;
			RECT	187.055 11.948 187.087 12.012 ;
			RECT	187.223 11.948 187.255 12.012 ;
			RECT	187.391 11.948 187.423 12.012 ;
			RECT	187.559 11.948 187.591 12.012 ;
			RECT	187.727 11.948 187.759 12.012 ;
			RECT	187.895 11.948 187.927 12.012 ;
			RECT	188.063 11.948 188.095 12.012 ;
			RECT	188.231 11.948 188.263 12.012 ;
			RECT	188.399 11.948 188.431 12.012 ;
			RECT	188.567 11.948 188.599 12.012 ;
			RECT	188.735 11.948 188.767 12.012 ;
			RECT	188.903 11.948 188.935 12.012 ;
			RECT	189.071 11.948 189.103 12.012 ;
			RECT	189.239 11.948 189.271 12.012 ;
			RECT	189.407 11.948 189.439 12.012 ;
			RECT	189.575 11.948 189.607 12.012 ;
			RECT	189.743 11.948 189.775 12.012 ;
			RECT	189.911 11.948 189.943 12.012 ;
			RECT	190.079 11.948 190.111 12.012 ;
			RECT	190.247 11.948 190.279 12.012 ;
			RECT	190.415 11.948 190.447 12.012 ;
			RECT	190.583 11.948 190.615 12.012 ;
			RECT	190.751 11.948 190.783 12.012 ;
			RECT	190.919 11.948 190.951 12.012 ;
			RECT	191.087 11.948 191.119 12.012 ;
			RECT	191.255 11.948 191.287 12.012 ;
			RECT	191.423 11.948 191.455 12.012 ;
			RECT	191.591 11.948 191.623 12.012 ;
			RECT	191.759 11.948 191.791 12.012 ;
			RECT	191.927 11.948 191.959 12.012 ;
			RECT	192.095 11.948 192.127 12.012 ;
			RECT	192.263 11.948 192.295 12.012 ;
			RECT	192.431 11.948 192.463 12.012 ;
			RECT	192.599 11.948 192.631 12.012 ;
			RECT	192.767 11.948 192.799 12.012 ;
			RECT	192.935 11.948 192.967 12.012 ;
			RECT	193.103 11.948 193.135 12.012 ;
			RECT	193.271 11.948 193.303 12.012 ;
			RECT	193.439 11.948 193.471 12.012 ;
			RECT	193.607 11.948 193.639 12.012 ;
			RECT	193.775 11.948 193.807 12.012 ;
			RECT	193.943 11.948 193.975 12.012 ;
			RECT	194.111 11.948 194.143 12.012 ;
			RECT	194.279 11.948 194.311 12.012 ;
			RECT	194.447 11.948 194.479 12.012 ;
			RECT	194.615 11.948 194.647 12.012 ;
			RECT	194.783 11.948 194.815 12.012 ;
			RECT	194.951 11.948 194.983 12.012 ;
			RECT	195.119 11.948 195.151 12.012 ;
			RECT	195.287 11.948 195.319 12.012 ;
			RECT	195.455 11.948 195.487 12.012 ;
			RECT	195.623 11.948 195.655 12.012 ;
			RECT	195.791 11.948 195.823 12.012 ;
			RECT	195.959 11.948 195.991 12.012 ;
			RECT	196.127 11.948 196.159 12.012 ;
			RECT	196.295 11.948 196.327 12.012 ;
			RECT	196.463 11.948 196.495 12.012 ;
			RECT	196.631 11.948 196.663 12.012 ;
			RECT	196.799 11.948 196.831 12.012 ;
			RECT	196.967 11.948 196.999 12.012 ;
			RECT	197.135 11.948 197.167 12.012 ;
			RECT	197.303 11.948 197.335 12.012 ;
			RECT	197.471 11.948 197.503 12.012 ;
			RECT	197.639 11.948 197.671 12.012 ;
			RECT	197.807 11.948 197.839 12.012 ;
			RECT	197.975 11.948 198.007 12.012 ;
			RECT	198.143 11.948 198.175 12.012 ;
			RECT	198.311 11.948 198.343 12.012 ;
			RECT	198.479 11.948 198.511 12.012 ;
			RECT	198.647 11.948 198.679 12.012 ;
			RECT	198.815 11.948 198.847 12.012 ;
			RECT	198.983 11.948 199.015 12.012 ;
			RECT	199.151 11.948 199.183 12.012 ;
			RECT	199.319 11.948 199.351 12.012 ;
			RECT	199.487 11.948 199.519 12.012 ;
			RECT	199.655 11.948 199.687 12.012 ;
			RECT	199.823 11.948 199.855 12.012 ;
			RECT	199.991 11.948 200.023 12.012 ;
			RECT	200.121 11.964 200.153 11.996 ;
			RECT	200.243 11.969 200.275 12.001 ;
			RECT	200.373 11.948 200.405 12.012 ;
			RECT	200.9 11.948 200.932 12.012 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 10 201.665 10.12 ;
			LAYER	J3 ;
			RECT	0.755 10.028 0.787 10.092 ;
			RECT	1.645 10.028 1.709 10.092 ;
			RECT	2.323 10.028 2.387 10.092 ;
			RECT	3.438 10.028 3.47 10.092 ;
			RECT	3.585 10.028 3.617 10.092 ;
			RECT	4.195 10.028 4.227 10.092 ;
			RECT	4.72 10.028 4.752 10.092 ;
			RECT	4.944 10.028 5.008 10.092 ;
			RECT	5.267 10.028 5.299 10.092 ;
			RECT	5.797 10.028 5.829 10.092 ;
			RECT	5.927 10.049 5.959 10.081 ;
			RECT	6.049 10.044 6.081 10.076 ;
			RECT	6.179 10.028 6.211 10.092 ;
			RECT	6.347 10.028 6.379 10.092 ;
			RECT	6.515 10.028 6.547 10.092 ;
			RECT	6.683 10.028 6.715 10.092 ;
			RECT	6.851 10.028 6.883 10.092 ;
			RECT	7.019 10.028 7.051 10.092 ;
			RECT	7.187 10.028 7.219 10.092 ;
			RECT	7.355 10.028 7.387 10.092 ;
			RECT	7.523 10.028 7.555 10.092 ;
			RECT	7.691 10.028 7.723 10.092 ;
			RECT	7.859 10.028 7.891 10.092 ;
			RECT	8.027 10.028 8.059 10.092 ;
			RECT	8.195 10.028 8.227 10.092 ;
			RECT	8.363 10.028 8.395 10.092 ;
			RECT	8.531 10.028 8.563 10.092 ;
			RECT	8.699 10.028 8.731 10.092 ;
			RECT	8.867 10.028 8.899 10.092 ;
			RECT	9.035 10.028 9.067 10.092 ;
			RECT	9.203 10.028 9.235 10.092 ;
			RECT	9.371 10.028 9.403 10.092 ;
			RECT	9.539 10.028 9.571 10.092 ;
			RECT	9.707 10.028 9.739 10.092 ;
			RECT	9.875 10.028 9.907 10.092 ;
			RECT	10.043 10.028 10.075 10.092 ;
			RECT	10.211 10.028 10.243 10.092 ;
			RECT	10.379 10.028 10.411 10.092 ;
			RECT	10.547 10.028 10.579 10.092 ;
			RECT	10.715 10.028 10.747 10.092 ;
			RECT	10.883 10.028 10.915 10.092 ;
			RECT	11.051 10.028 11.083 10.092 ;
			RECT	11.219 10.028 11.251 10.092 ;
			RECT	11.387 10.028 11.419 10.092 ;
			RECT	11.555 10.028 11.587 10.092 ;
			RECT	11.723 10.028 11.755 10.092 ;
			RECT	11.891 10.028 11.923 10.092 ;
			RECT	12.059 10.028 12.091 10.092 ;
			RECT	12.227 10.028 12.259 10.092 ;
			RECT	12.395 10.028 12.427 10.092 ;
			RECT	12.563 10.028 12.595 10.092 ;
			RECT	12.731 10.028 12.763 10.092 ;
			RECT	12.899 10.028 12.931 10.092 ;
			RECT	13.067 10.028 13.099 10.092 ;
			RECT	13.235 10.028 13.267 10.092 ;
			RECT	13.403 10.028 13.435 10.092 ;
			RECT	13.571 10.028 13.603 10.092 ;
			RECT	13.739 10.028 13.771 10.092 ;
			RECT	13.907 10.028 13.939 10.092 ;
			RECT	14.075 10.028 14.107 10.092 ;
			RECT	14.243 10.028 14.275 10.092 ;
			RECT	14.411 10.028 14.443 10.092 ;
			RECT	14.579 10.028 14.611 10.092 ;
			RECT	14.747 10.028 14.779 10.092 ;
			RECT	14.915 10.028 14.947 10.092 ;
			RECT	15.083 10.028 15.115 10.092 ;
			RECT	15.251 10.028 15.283 10.092 ;
			RECT	15.419 10.028 15.451 10.092 ;
			RECT	15.587 10.028 15.619 10.092 ;
			RECT	15.755 10.028 15.787 10.092 ;
			RECT	15.923 10.028 15.955 10.092 ;
			RECT	16.091 10.028 16.123 10.092 ;
			RECT	16.259 10.028 16.291 10.092 ;
			RECT	16.427 10.028 16.459 10.092 ;
			RECT	16.595 10.028 16.627 10.092 ;
			RECT	16.763 10.028 16.795 10.092 ;
			RECT	16.931 10.028 16.963 10.092 ;
			RECT	17.099 10.028 17.131 10.092 ;
			RECT	17.267 10.028 17.299 10.092 ;
			RECT	17.435 10.028 17.467 10.092 ;
			RECT	17.603 10.028 17.635 10.092 ;
			RECT	17.771 10.028 17.803 10.092 ;
			RECT	17.939 10.028 17.971 10.092 ;
			RECT	18.107 10.028 18.139 10.092 ;
			RECT	18.275 10.028 18.307 10.092 ;
			RECT	18.443 10.028 18.475 10.092 ;
			RECT	18.611 10.028 18.643 10.092 ;
			RECT	18.779 10.028 18.811 10.092 ;
			RECT	18.947 10.028 18.979 10.092 ;
			RECT	19.115 10.028 19.147 10.092 ;
			RECT	19.283 10.028 19.315 10.092 ;
			RECT	19.451 10.028 19.483 10.092 ;
			RECT	19.619 10.028 19.651 10.092 ;
			RECT	19.787 10.028 19.819 10.092 ;
			RECT	19.955 10.028 19.987 10.092 ;
			RECT	20.123 10.028 20.155 10.092 ;
			RECT	20.291 10.028 20.323 10.092 ;
			RECT	20.459 10.028 20.491 10.092 ;
			RECT	20.627 10.028 20.659 10.092 ;
			RECT	20.795 10.028 20.827 10.092 ;
			RECT	20.963 10.028 20.995 10.092 ;
			RECT	21.131 10.028 21.163 10.092 ;
			RECT	21.299 10.028 21.331 10.092 ;
			RECT	21.467 10.028 21.499 10.092 ;
			RECT	21.635 10.028 21.667 10.092 ;
			RECT	21.803 10.028 21.835 10.092 ;
			RECT	21.971 10.028 22.003 10.092 ;
			RECT	22.139 10.028 22.171 10.092 ;
			RECT	22.307 10.028 22.339 10.092 ;
			RECT	22.475 10.028 22.507 10.092 ;
			RECT	22.643 10.028 22.675 10.092 ;
			RECT	22.811 10.028 22.843 10.092 ;
			RECT	22.979 10.028 23.011 10.092 ;
			RECT	23.147 10.028 23.179 10.092 ;
			RECT	23.315 10.028 23.347 10.092 ;
			RECT	23.483 10.028 23.515 10.092 ;
			RECT	23.651 10.028 23.683 10.092 ;
			RECT	23.819 10.028 23.851 10.092 ;
			RECT	23.987 10.028 24.019 10.092 ;
			RECT	24.155 10.028 24.187 10.092 ;
			RECT	24.323 10.028 24.355 10.092 ;
			RECT	24.491 10.028 24.523 10.092 ;
			RECT	24.659 10.028 24.691 10.092 ;
			RECT	24.827 10.028 24.859 10.092 ;
			RECT	24.995 10.028 25.027 10.092 ;
			RECT	25.163 10.028 25.195 10.092 ;
			RECT	25.331 10.028 25.363 10.092 ;
			RECT	25.499 10.028 25.531 10.092 ;
			RECT	25.667 10.028 25.699 10.092 ;
			RECT	25.835 10.028 25.867 10.092 ;
			RECT	26.003 10.028 26.035 10.092 ;
			RECT	26.171 10.028 26.203 10.092 ;
			RECT	26.339 10.028 26.371 10.092 ;
			RECT	26.507 10.028 26.539 10.092 ;
			RECT	26.675 10.028 26.707 10.092 ;
			RECT	26.843 10.028 26.875 10.092 ;
			RECT	27.011 10.028 27.043 10.092 ;
			RECT	27.179 10.028 27.211 10.092 ;
			RECT	27.347 10.028 27.379 10.092 ;
			RECT	27.515 10.028 27.547 10.092 ;
			RECT	27.683 10.028 27.715 10.092 ;
			RECT	27.851 10.028 27.883 10.092 ;
			RECT	28.019 10.028 28.051 10.092 ;
			RECT	28.187 10.028 28.219 10.092 ;
			RECT	28.355 10.028 28.387 10.092 ;
			RECT	28.523 10.028 28.555 10.092 ;
			RECT	28.691 10.028 28.723 10.092 ;
			RECT	28.859 10.028 28.891 10.092 ;
			RECT	29.027 10.028 29.059 10.092 ;
			RECT	29.195 10.028 29.227 10.092 ;
			RECT	29.363 10.028 29.395 10.092 ;
			RECT	29.531 10.028 29.563 10.092 ;
			RECT	29.699 10.028 29.731 10.092 ;
			RECT	29.867 10.028 29.899 10.092 ;
			RECT	30.035 10.028 30.067 10.092 ;
			RECT	30.203 10.028 30.235 10.092 ;
			RECT	30.371 10.028 30.403 10.092 ;
			RECT	30.539 10.028 30.571 10.092 ;
			RECT	30.707 10.028 30.739 10.092 ;
			RECT	30.875 10.028 30.907 10.092 ;
			RECT	31.043 10.028 31.075 10.092 ;
			RECT	31.211 10.028 31.243 10.092 ;
			RECT	31.379 10.028 31.411 10.092 ;
			RECT	31.547 10.028 31.579 10.092 ;
			RECT	31.715 10.028 31.747 10.092 ;
			RECT	31.883 10.028 31.915 10.092 ;
			RECT	32.051 10.028 32.083 10.092 ;
			RECT	32.219 10.028 32.251 10.092 ;
			RECT	32.387 10.028 32.419 10.092 ;
			RECT	32.555 10.028 32.587 10.092 ;
			RECT	32.723 10.028 32.755 10.092 ;
			RECT	32.891 10.028 32.923 10.092 ;
			RECT	33.059 10.028 33.091 10.092 ;
			RECT	33.227 10.028 33.259 10.092 ;
			RECT	33.395 10.028 33.427 10.092 ;
			RECT	33.563 10.028 33.595 10.092 ;
			RECT	33.731 10.028 33.763 10.092 ;
			RECT	33.899 10.028 33.931 10.092 ;
			RECT	34.067 10.028 34.099 10.092 ;
			RECT	34.235 10.028 34.267 10.092 ;
			RECT	34.403 10.028 34.435 10.092 ;
			RECT	34.571 10.028 34.603 10.092 ;
			RECT	34.739 10.028 34.771 10.092 ;
			RECT	34.907 10.028 34.939 10.092 ;
			RECT	35.075 10.028 35.107 10.092 ;
			RECT	35.243 10.028 35.275 10.092 ;
			RECT	35.411 10.028 35.443 10.092 ;
			RECT	35.579 10.028 35.611 10.092 ;
			RECT	35.747 10.028 35.779 10.092 ;
			RECT	35.915 10.028 35.947 10.092 ;
			RECT	36.083 10.028 36.115 10.092 ;
			RECT	36.251 10.028 36.283 10.092 ;
			RECT	36.419 10.028 36.451 10.092 ;
			RECT	36.587 10.028 36.619 10.092 ;
			RECT	36.755 10.028 36.787 10.092 ;
			RECT	36.923 10.028 36.955 10.092 ;
			RECT	37.091 10.028 37.123 10.092 ;
			RECT	37.259 10.028 37.291 10.092 ;
			RECT	37.427 10.028 37.459 10.092 ;
			RECT	37.595 10.028 37.627 10.092 ;
			RECT	37.763 10.028 37.795 10.092 ;
			RECT	37.931 10.028 37.963 10.092 ;
			RECT	38.099 10.028 38.131 10.092 ;
			RECT	38.267 10.028 38.299 10.092 ;
			RECT	38.435 10.028 38.467 10.092 ;
			RECT	38.603 10.028 38.635 10.092 ;
			RECT	38.771 10.028 38.803 10.092 ;
			RECT	38.939 10.028 38.971 10.092 ;
			RECT	39.107 10.028 39.139 10.092 ;
			RECT	39.275 10.028 39.307 10.092 ;
			RECT	39.443 10.028 39.475 10.092 ;
			RECT	39.611 10.028 39.643 10.092 ;
			RECT	39.779 10.028 39.811 10.092 ;
			RECT	39.947 10.028 39.979 10.092 ;
			RECT	40.115 10.028 40.147 10.092 ;
			RECT	40.283 10.028 40.315 10.092 ;
			RECT	40.451 10.028 40.483 10.092 ;
			RECT	40.619 10.028 40.651 10.092 ;
			RECT	40.787 10.028 40.819 10.092 ;
			RECT	40.955 10.028 40.987 10.092 ;
			RECT	41.123 10.028 41.155 10.092 ;
			RECT	41.291 10.028 41.323 10.092 ;
			RECT	41.459 10.028 41.491 10.092 ;
			RECT	41.627 10.028 41.659 10.092 ;
			RECT	41.795 10.028 41.827 10.092 ;
			RECT	41.963 10.028 41.995 10.092 ;
			RECT	42.131 10.028 42.163 10.092 ;
			RECT	42.299 10.028 42.331 10.092 ;
			RECT	42.467 10.028 42.499 10.092 ;
			RECT	42.635 10.028 42.667 10.092 ;
			RECT	42.803 10.028 42.835 10.092 ;
			RECT	42.971 10.028 43.003 10.092 ;
			RECT	43.139 10.028 43.171 10.092 ;
			RECT	43.307 10.028 43.339 10.092 ;
			RECT	43.475 10.028 43.507 10.092 ;
			RECT	43.643 10.028 43.675 10.092 ;
			RECT	43.811 10.028 43.843 10.092 ;
			RECT	43.979 10.028 44.011 10.092 ;
			RECT	44.147 10.028 44.179 10.092 ;
			RECT	44.315 10.028 44.347 10.092 ;
			RECT	44.483 10.028 44.515 10.092 ;
			RECT	44.651 10.028 44.683 10.092 ;
			RECT	44.819 10.028 44.851 10.092 ;
			RECT	44.987 10.028 45.019 10.092 ;
			RECT	45.155 10.028 45.187 10.092 ;
			RECT	45.323 10.028 45.355 10.092 ;
			RECT	45.491 10.028 45.523 10.092 ;
			RECT	45.659 10.028 45.691 10.092 ;
			RECT	45.827 10.028 45.859 10.092 ;
			RECT	45.995 10.028 46.027 10.092 ;
			RECT	46.163 10.028 46.195 10.092 ;
			RECT	46.331 10.028 46.363 10.092 ;
			RECT	46.499 10.028 46.531 10.092 ;
			RECT	46.667 10.028 46.699 10.092 ;
			RECT	46.835 10.028 46.867 10.092 ;
			RECT	47.003 10.028 47.035 10.092 ;
			RECT	47.171 10.028 47.203 10.092 ;
			RECT	47.339 10.028 47.371 10.092 ;
			RECT	47.507 10.028 47.539 10.092 ;
			RECT	47.675 10.028 47.707 10.092 ;
			RECT	47.843 10.028 47.875 10.092 ;
			RECT	48.011 10.028 48.043 10.092 ;
			RECT	48.179 10.028 48.211 10.092 ;
			RECT	48.347 10.028 48.379 10.092 ;
			RECT	48.515 10.028 48.547 10.092 ;
			RECT	48.683 10.028 48.715 10.092 ;
			RECT	48.851 10.028 48.883 10.092 ;
			RECT	49.019 10.028 49.051 10.092 ;
			RECT	49.187 10.028 49.219 10.092 ;
			RECT	49.318 10.044 49.35 10.076 ;
			RECT	49.439 10.044 49.471 10.076 ;
			RECT	49.569 10.028 49.601 10.092 ;
			RECT	51.881 10.028 51.913 10.092 ;
			RECT	53.132 10.028 53.196 10.092 ;
			RECT	53.812 10.028 53.844 10.092 ;
			RECT	54.251 10.028 54.283 10.092 ;
			RECT	55.562 10.028 55.626 10.092 ;
			RECT	58.603 10.028 58.635 10.092 ;
			RECT	58.733 10.044 58.765 10.076 ;
			RECT	58.854 10.044 58.886 10.076 ;
			RECT	58.985 10.028 59.017 10.092 ;
			RECT	59.153 10.028 59.185 10.092 ;
			RECT	59.321 10.028 59.353 10.092 ;
			RECT	59.489 10.028 59.521 10.092 ;
			RECT	59.657 10.028 59.689 10.092 ;
			RECT	59.825 10.028 59.857 10.092 ;
			RECT	59.993 10.028 60.025 10.092 ;
			RECT	60.161 10.028 60.193 10.092 ;
			RECT	60.329 10.028 60.361 10.092 ;
			RECT	60.497 10.028 60.529 10.092 ;
			RECT	60.665 10.028 60.697 10.092 ;
			RECT	60.833 10.028 60.865 10.092 ;
			RECT	61.001 10.028 61.033 10.092 ;
			RECT	61.169 10.028 61.201 10.092 ;
			RECT	61.337 10.028 61.369 10.092 ;
			RECT	61.505 10.028 61.537 10.092 ;
			RECT	61.673 10.028 61.705 10.092 ;
			RECT	61.841 10.028 61.873 10.092 ;
			RECT	62.009 10.028 62.041 10.092 ;
			RECT	62.177 10.028 62.209 10.092 ;
			RECT	62.345 10.028 62.377 10.092 ;
			RECT	62.513 10.028 62.545 10.092 ;
			RECT	62.681 10.028 62.713 10.092 ;
			RECT	62.849 10.028 62.881 10.092 ;
			RECT	63.017 10.028 63.049 10.092 ;
			RECT	63.185 10.028 63.217 10.092 ;
			RECT	63.353 10.028 63.385 10.092 ;
			RECT	63.521 10.028 63.553 10.092 ;
			RECT	63.689 10.028 63.721 10.092 ;
			RECT	63.857 10.028 63.889 10.092 ;
			RECT	64.025 10.028 64.057 10.092 ;
			RECT	64.193 10.028 64.225 10.092 ;
			RECT	64.361 10.028 64.393 10.092 ;
			RECT	64.529 10.028 64.561 10.092 ;
			RECT	64.697 10.028 64.729 10.092 ;
			RECT	64.865 10.028 64.897 10.092 ;
			RECT	65.033 10.028 65.065 10.092 ;
			RECT	65.201 10.028 65.233 10.092 ;
			RECT	65.369 10.028 65.401 10.092 ;
			RECT	65.537 10.028 65.569 10.092 ;
			RECT	65.705 10.028 65.737 10.092 ;
			RECT	65.873 10.028 65.905 10.092 ;
			RECT	66.041 10.028 66.073 10.092 ;
			RECT	66.209 10.028 66.241 10.092 ;
			RECT	66.377 10.028 66.409 10.092 ;
			RECT	66.545 10.028 66.577 10.092 ;
			RECT	66.713 10.028 66.745 10.092 ;
			RECT	66.881 10.028 66.913 10.092 ;
			RECT	67.049 10.028 67.081 10.092 ;
			RECT	67.217 10.028 67.249 10.092 ;
			RECT	67.385 10.028 67.417 10.092 ;
			RECT	67.553 10.028 67.585 10.092 ;
			RECT	67.721 10.028 67.753 10.092 ;
			RECT	67.889 10.028 67.921 10.092 ;
			RECT	68.057 10.028 68.089 10.092 ;
			RECT	68.225 10.028 68.257 10.092 ;
			RECT	68.393 10.028 68.425 10.092 ;
			RECT	68.561 10.028 68.593 10.092 ;
			RECT	68.729 10.028 68.761 10.092 ;
			RECT	68.897 10.028 68.929 10.092 ;
			RECT	69.065 10.028 69.097 10.092 ;
			RECT	69.233 10.028 69.265 10.092 ;
			RECT	69.401 10.028 69.433 10.092 ;
			RECT	69.569 10.028 69.601 10.092 ;
			RECT	69.737 10.028 69.769 10.092 ;
			RECT	69.905 10.028 69.937 10.092 ;
			RECT	70.073 10.028 70.105 10.092 ;
			RECT	70.241 10.028 70.273 10.092 ;
			RECT	70.409 10.028 70.441 10.092 ;
			RECT	70.577 10.028 70.609 10.092 ;
			RECT	70.745 10.028 70.777 10.092 ;
			RECT	70.913 10.028 70.945 10.092 ;
			RECT	71.081 10.028 71.113 10.092 ;
			RECT	71.249 10.028 71.281 10.092 ;
			RECT	71.417 10.028 71.449 10.092 ;
			RECT	71.585 10.028 71.617 10.092 ;
			RECT	71.753 10.028 71.785 10.092 ;
			RECT	71.921 10.028 71.953 10.092 ;
			RECT	72.089 10.028 72.121 10.092 ;
			RECT	72.257 10.028 72.289 10.092 ;
			RECT	72.425 10.028 72.457 10.092 ;
			RECT	72.593 10.028 72.625 10.092 ;
			RECT	72.761 10.028 72.793 10.092 ;
			RECT	72.929 10.028 72.961 10.092 ;
			RECT	73.097 10.028 73.129 10.092 ;
			RECT	73.265 10.028 73.297 10.092 ;
			RECT	73.433 10.028 73.465 10.092 ;
			RECT	73.601 10.028 73.633 10.092 ;
			RECT	73.769 10.028 73.801 10.092 ;
			RECT	73.937 10.028 73.969 10.092 ;
			RECT	74.105 10.028 74.137 10.092 ;
			RECT	74.273 10.028 74.305 10.092 ;
			RECT	74.441 10.028 74.473 10.092 ;
			RECT	74.609 10.028 74.641 10.092 ;
			RECT	74.777 10.028 74.809 10.092 ;
			RECT	74.945 10.028 74.977 10.092 ;
			RECT	75.113 10.028 75.145 10.092 ;
			RECT	75.281 10.028 75.313 10.092 ;
			RECT	75.449 10.028 75.481 10.092 ;
			RECT	75.617 10.028 75.649 10.092 ;
			RECT	75.785 10.028 75.817 10.092 ;
			RECT	75.953 10.028 75.985 10.092 ;
			RECT	76.121 10.028 76.153 10.092 ;
			RECT	76.289 10.028 76.321 10.092 ;
			RECT	76.457 10.028 76.489 10.092 ;
			RECT	76.625 10.028 76.657 10.092 ;
			RECT	76.793 10.028 76.825 10.092 ;
			RECT	76.961 10.028 76.993 10.092 ;
			RECT	77.129 10.028 77.161 10.092 ;
			RECT	77.297 10.028 77.329 10.092 ;
			RECT	77.465 10.028 77.497 10.092 ;
			RECT	77.633 10.028 77.665 10.092 ;
			RECT	77.801 10.028 77.833 10.092 ;
			RECT	77.969 10.028 78.001 10.092 ;
			RECT	78.137 10.028 78.169 10.092 ;
			RECT	78.305 10.028 78.337 10.092 ;
			RECT	78.473 10.028 78.505 10.092 ;
			RECT	78.641 10.028 78.673 10.092 ;
			RECT	78.809 10.028 78.841 10.092 ;
			RECT	78.977 10.028 79.009 10.092 ;
			RECT	79.145 10.028 79.177 10.092 ;
			RECT	79.313 10.028 79.345 10.092 ;
			RECT	79.481 10.028 79.513 10.092 ;
			RECT	79.649 10.028 79.681 10.092 ;
			RECT	79.817 10.028 79.849 10.092 ;
			RECT	79.985 10.028 80.017 10.092 ;
			RECT	80.153 10.028 80.185 10.092 ;
			RECT	80.321 10.028 80.353 10.092 ;
			RECT	80.489 10.028 80.521 10.092 ;
			RECT	80.657 10.028 80.689 10.092 ;
			RECT	80.825 10.028 80.857 10.092 ;
			RECT	80.993 10.028 81.025 10.092 ;
			RECT	81.161 10.028 81.193 10.092 ;
			RECT	81.329 10.028 81.361 10.092 ;
			RECT	81.497 10.028 81.529 10.092 ;
			RECT	81.665 10.028 81.697 10.092 ;
			RECT	81.833 10.028 81.865 10.092 ;
			RECT	82.001 10.028 82.033 10.092 ;
			RECT	82.169 10.028 82.201 10.092 ;
			RECT	82.337 10.028 82.369 10.092 ;
			RECT	82.505 10.028 82.537 10.092 ;
			RECT	82.673 10.028 82.705 10.092 ;
			RECT	82.841 10.028 82.873 10.092 ;
			RECT	83.009 10.028 83.041 10.092 ;
			RECT	83.177 10.028 83.209 10.092 ;
			RECT	83.345 10.028 83.377 10.092 ;
			RECT	83.513 10.028 83.545 10.092 ;
			RECT	83.681 10.028 83.713 10.092 ;
			RECT	83.849 10.028 83.881 10.092 ;
			RECT	84.017 10.028 84.049 10.092 ;
			RECT	84.185 10.028 84.217 10.092 ;
			RECT	84.353 10.028 84.385 10.092 ;
			RECT	84.521 10.028 84.553 10.092 ;
			RECT	84.689 10.028 84.721 10.092 ;
			RECT	84.857 10.028 84.889 10.092 ;
			RECT	85.025 10.028 85.057 10.092 ;
			RECT	85.193 10.028 85.225 10.092 ;
			RECT	85.361 10.028 85.393 10.092 ;
			RECT	85.529 10.028 85.561 10.092 ;
			RECT	85.697 10.028 85.729 10.092 ;
			RECT	85.865 10.028 85.897 10.092 ;
			RECT	86.033 10.028 86.065 10.092 ;
			RECT	86.201 10.028 86.233 10.092 ;
			RECT	86.369 10.028 86.401 10.092 ;
			RECT	86.537 10.028 86.569 10.092 ;
			RECT	86.705 10.028 86.737 10.092 ;
			RECT	86.873 10.028 86.905 10.092 ;
			RECT	87.041 10.028 87.073 10.092 ;
			RECT	87.209 10.028 87.241 10.092 ;
			RECT	87.377 10.028 87.409 10.092 ;
			RECT	87.545 10.028 87.577 10.092 ;
			RECT	87.713 10.028 87.745 10.092 ;
			RECT	87.881 10.028 87.913 10.092 ;
			RECT	88.049 10.028 88.081 10.092 ;
			RECT	88.217 10.028 88.249 10.092 ;
			RECT	88.385 10.028 88.417 10.092 ;
			RECT	88.553 10.028 88.585 10.092 ;
			RECT	88.721 10.028 88.753 10.092 ;
			RECT	88.889 10.028 88.921 10.092 ;
			RECT	89.057 10.028 89.089 10.092 ;
			RECT	89.225 10.028 89.257 10.092 ;
			RECT	89.393 10.028 89.425 10.092 ;
			RECT	89.561 10.028 89.593 10.092 ;
			RECT	89.729 10.028 89.761 10.092 ;
			RECT	89.897 10.028 89.929 10.092 ;
			RECT	90.065 10.028 90.097 10.092 ;
			RECT	90.233 10.028 90.265 10.092 ;
			RECT	90.401 10.028 90.433 10.092 ;
			RECT	90.569 10.028 90.601 10.092 ;
			RECT	90.737 10.028 90.769 10.092 ;
			RECT	90.905 10.028 90.937 10.092 ;
			RECT	91.073 10.028 91.105 10.092 ;
			RECT	91.241 10.028 91.273 10.092 ;
			RECT	91.409 10.028 91.441 10.092 ;
			RECT	91.577 10.028 91.609 10.092 ;
			RECT	91.745 10.028 91.777 10.092 ;
			RECT	91.913 10.028 91.945 10.092 ;
			RECT	92.081 10.028 92.113 10.092 ;
			RECT	92.249 10.028 92.281 10.092 ;
			RECT	92.417 10.028 92.449 10.092 ;
			RECT	92.585 10.028 92.617 10.092 ;
			RECT	92.753 10.028 92.785 10.092 ;
			RECT	92.921 10.028 92.953 10.092 ;
			RECT	93.089 10.028 93.121 10.092 ;
			RECT	93.257 10.028 93.289 10.092 ;
			RECT	93.425 10.028 93.457 10.092 ;
			RECT	93.593 10.028 93.625 10.092 ;
			RECT	93.761 10.028 93.793 10.092 ;
			RECT	93.929 10.028 93.961 10.092 ;
			RECT	94.097 10.028 94.129 10.092 ;
			RECT	94.265 10.028 94.297 10.092 ;
			RECT	94.433 10.028 94.465 10.092 ;
			RECT	94.601 10.028 94.633 10.092 ;
			RECT	94.769 10.028 94.801 10.092 ;
			RECT	94.937 10.028 94.969 10.092 ;
			RECT	95.105 10.028 95.137 10.092 ;
			RECT	95.273 10.028 95.305 10.092 ;
			RECT	95.441 10.028 95.473 10.092 ;
			RECT	95.609 10.028 95.641 10.092 ;
			RECT	95.777 10.028 95.809 10.092 ;
			RECT	95.945 10.028 95.977 10.092 ;
			RECT	96.113 10.028 96.145 10.092 ;
			RECT	96.281 10.028 96.313 10.092 ;
			RECT	96.449 10.028 96.481 10.092 ;
			RECT	96.617 10.028 96.649 10.092 ;
			RECT	96.785 10.028 96.817 10.092 ;
			RECT	96.953 10.028 96.985 10.092 ;
			RECT	97.121 10.028 97.153 10.092 ;
			RECT	97.289 10.028 97.321 10.092 ;
			RECT	97.457 10.028 97.489 10.092 ;
			RECT	97.625 10.028 97.657 10.092 ;
			RECT	97.793 10.028 97.825 10.092 ;
			RECT	97.961 10.028 97.993 10.092 ;
			RECT	98.129 10.028 98.161 10.092 ;
			RECT	98.297 10.028 98.329 10.092 ;
			RECT	98.465 10.028 98.497 10.092 ;
			RECT	98.633 10.028 98.665 10.092 ;
			RECT	98.801 10.028 98.833 10.092 ;
			RECT	98.969 10.028 99.001 10.092 ;
			RECT	99.137 10.028 99.169 10.092 ;
			RECT	99.305 10.028 99.337 10.092 ;
			RECT	99.473 10.028 99.505 10.092 ;
			RECT	99.641 10.028 99.673 10.092 ;
			RECT	99.809 10.028 99.841 10.092 ;
			RECT	99.977 10.028 100.009 10.092 ;
			RECT	100.145 10.028 100.177 10.092 ;
			RECT	100.313 10.028 100.345 10.092 ;
			RECT	100.481 10.028 100.513 10.092 ;
			RECT	100.649 10.028 100.681 10.092 ;
			RECT	100.817 10.028 100.849 10.092 ;
			RECT	100.985 10.028 101.017 10.092 ;
			RECT	101.153 10.028 101.185 10.092 ;
			RECT	101.321 10.028 101.353 10.092 ;
			RECT	101.489 10.028 101.521 10.092 ;
			RECT	101.657 10.028 101.689 10.092 ;
			RECT	101.825 10.028 101.857 10.092 ;
			RECT	101.993 10.028 102.025 10.092 ;
			RECT	102.123 10.044 102.155 10.076 ;
			RECT	102.245 10.049 102.277 10.081 ;
			RECT	102.375 10.028 102.407 10.092 ;
			RECT	103.795 10.028 103.827 10.092 ;
			RECT	103.925 10.049 103.957 10.081 ;
			RECT	104.047 10.044 104.079 10.076 ;
			RECT	104.177 10.028 104.209 10.092 ;
			RECT	104.345 10.028 104.377 10.092 ;
			RECT	104.513 10.028 104.545 10.092 ;
			RECT	104.681 10.028 104.713 10.092 ;
			RECT	104.849 10.028 104.881 10.092 ;
			RECT	105.017 10.028 105.049 10.092 ;
			RECT	105.185 10.028 105.217 10.092 ;
			RECT	105.353 10.028 105.385 10.092 ;
			RECT	105.521 10.028 105.553 10.092 ;
			RECT	105.689 10.028 105.721 10.092 ;
			RECT	105.857 10.028 105.889 10.092 ;
			RECT	106.025 10.028 106.057 10.092 ;
			RECT	106.193 10.028 106.225 10.092 ;
			RECT	106.361 10.028 106.393 10.092 ;
			RECT	106.529 10.028 106.561 10.092 ;
			RECT	106.697 10.028 106.729 10.092 ;
			RECT	106.865 10.028 106.897 10.092 ;
			RECT	107.033 10.028 107.065 10.092 ;
			RECT	107.201 10.028 107.233 10.092 ;
			RECT	107.369 10.028 107.401 10.092 ;
			RECT	107.537 10.028 107.569 10.092 ;
			RECT	107.705 10.028 107.737 10.092 ;
			RECT	107.873 10.028 107.905 10.092 ;
			RECT	108.041 10.028 108.073 10.092 ;
			RECT	108.209 10.028 108.241 10.092 ;
			RECT	108.377 10.028 108.409 10.092 ;
			RECT	108.545 10.028 108.577 10.092 ;
			RECT	108.713 10.028 108.745 10.092 ;
			RECT	108.881 10.028 108.913 10.092 ;
			RECT	109.049 10.028 109.081 10.092 ;
			RECT	109.217 10.028 109.249 10.092 ;
			RECT	109.385 10.028 109.417 10.092 ;
			RECT	109.553 10.028 109.585 10.092 ;
			RECT	109.721 10.028 109.753 10.092 ;
			RECT	109.889 10.028 109.921 10.092 ;
			RECT	110.057 10.028 110.089 10.092 ;
			RECT	110.225 10.028 110.257 10.092 ;
			RECT	110.393 10.028 110.425 10.092 ;
			RECT	110.561 10.028 110.593 10.092 ;
			RECT	110.729 10.028 110.761 10.092 ;
			RECT	110.897 10.028 110.929 10.092 ;
			RECT	111.065 10.028 111.097 10.092 ;
			RECT	111.233 10.028 111.265 10.092 ;
			RECT	111.401 10.028 111.433 10.092 ;
			RECT	111.569 10.028 111.601 10.092 ;
			RECT	111.737 10.028 111.769 10.092 ;
			RECT	111.905 10.028 111.937 10.092 ;
			RECT	112.073 10.028 112.105 10.092 ;
			RECT	112.241 10.028 112.273 10.092 ;
			RECT	112.409 10.028 112.441 10.092 ;
			RECT	112.577 10.028 112.609 10.092 ;
			RECT	112.745 10.028 112.777 10.092 ;
			RECT	112.913 10.028 112.945 10.092 ;
			RECT	113.081 10.028 113.113 10.092 ;
			RECT	113.249 10.028 113.281 10.092 ;
			RECT	113.417 10.028 113.449 10.092 ;
			RECT	113.585 10.028 113.617 10.092 ;
			RECT	113.753 10.028 113.785 10.092 ;
			RECT	113.921 10.028 113.953 10.092 ;
			RECT	114.089 10.028 114.121 10.092 ;
			RECT	114.257 10.028 114.289 10.092 ;
			RECT	114.425 10.028 114.457 10.092 ;
			RECT	114.593 10.028 114.625 10.092 ;
			RECT	114.761 10.028 114.793 10.092 ;
			RECT	114.929 10.028 114.961 10.092 ;
			RECT	115.097 10.028 115.129 10.092 ;
			RECT	115.265 10.028 115.297 10.092 ;
			RECT	115.433 10.028 115.465 10.092 ;
			RECT	115.601 10.028 115.633 10.092 ;
			RECT	115.769 10.028 115.801 10.092 ;
			RECT	115.937 10.028 115.969 10.092 ;
			RECT	116.105 10.028 116.137 10.092 ;
			RECT	116.273 10.028 116.305 10.092 ;
			RECT	116.441 10.028 116.473 10.092 ;
			RECT	116.609 10.028 116.641 10.092 ;
			RECT	116.777 10.028 116.809 10.092 ;
			RECT	116.945 10.028 116.977 10.092 ;
			RECT	117.113 10.028 117.145 10.092 ;
			RECT	117.281 10.028 117.313 10.092 ;
			RECT	117.449 10.028 117.481 10.092 ;
			RECT	117.617 10.028 117.649 10.092 ;
			RECT	117.785 10.028 117.817 10.092 ;
			RECT	117.953 10.028 117.985 10.092 ;
			RECT	118.121 10.028 118.153 10.092 ;
			RECT	118.289 10.028 118.321 10.092 ;
			RECT	118.457 10.028 118.489 10.092 ;
			RECT	118.625 10.028 118.657 10.092 ;
			RECT	118.793 10.028 118.825 10.092 ;
			RECT	118.961 10.028 118.993 10.092 ;
			RECT	119.129 10.028 119.161 10.092 ;
			RECT	119.297 10.028 119.329 10.092 ;
			RECT	119.465 10.028 119.497 10.092 ;
			RECT	119.633 10.028 119.665 10.092 ;
			RECT	119.801 10.028 119.833 10.092 ;
			RECT	119.969 10.028 120.001 10.092 ;
			RECT	120.137 10.028 120.169 10.092 ;
			RECT	120.305 10.028 120.337 10.092 ;
			RECT	120.473 10.028 120.505 10.092 ;
			RECT	120.641 10.028 120.673 10.092 ;
			RECT	120.809 10.028 120.841 10.092 ;
			RECT	120.977 10.028 121.009 10.092 ;
			RECT	121.145 10.028 121.177 10.092 ;
			RECT	121.313 10.028 121.345 10.092 ;
			RECT	121.481 10.028 121.513 10.092 ;
			RECT	121.649 10.028 121.681 10.092 ;
			RECT	121.817 10.028 121.849 10.092 ;
			RECT	121.985 10.028 122.017 10.092 ;
			RECT	122.153 10.028 122.185 10.092 ;
			RECT	122.321 10.028 122.353 10.092 ;
			RECT	122.489 10.028 122.521 10.092 ;
			RECT	122.657 10.028 122.689 10.092 ;
			RECT	122.825 10.028 122.857 10.092 ;
			RECT	122.993 10.028 123.025 10.092 ;
			RECT	123.161 10.028 123.193 10.092 ;
			RECT	123.329 10.028 123.361 10.092 ;
			RECT	123.497 10.028 123.529 10.092 ;
			RECT	123.665 10.028 123.697 10.092 ;
			RECT	123.833 10.028 123.865 10.092 ;
			RECT	124.001 10.028 124.033 10.092 ;
			RECT	124.169 10.028 124.201 10.092 ;
			RECT	124.337 10.028 124.369 10.092 ;
			RECT	124.505 10.028 124.537 10.092 ;
			RECT	124.673 10.028 124.705 10.092 ;
			RECT	124.841 10.028 124.873 10.092 ;
			RECT	125.009 10.028 125.041 10.092 ;
			RECT	125.177 10.028 125.209 10.092 ;
			RECT	125.345 10.028 125.377 10.092 ;
			RECT	125.513 10.028 125.545 10.092 ;
			RECT	125.681 10.028 125.713 10.092 ;
			RECT	125.849 10.028 125.881 10.092 ;
			RECT	126.017 10.028 126.049 10.092 ;
			RECT	126.185 10.028 126.217 10.092 ;
			RECT	126.353 10.028 126.385 10.092 ;
			RECT	126.521 10.028 126.553 10.092 ;
			RECT	126.689 10.028 126.721 10.092 ;
			RECT	126.857 10.028 126.889 10.092 ;
			RECT	127.025 10.028 127.057 10.092 ;
			RECT	127.193 10.028 127.225 10.092 ;
			RECT	127.361 10.028 127.393 10.092 ;
			RECT	127.529 10.028 127.561 10.092 ;
			RECT	127.697 10.028 127.729 10.092 ;
			RECT	127.865 10.028 127.897 10.092 ;
			RECT	128.033 10.028 128.065 10.092 ;
			RECT	128.201 10.028 128.233 10.092 ;
			RECT	128.369 10.028 128.401 10.092 ;
			RECT	128.537 10.028 128.569 10.092 ;
			RECT	128.705 10.028 128.737 10.092 ;
			RECT	128.873 10.028 128.905 10.092 ;
			RECT	129.041 10.028 129.073 10.092 ;
			RECT	129.209 10.028 129.241 10.092 ;
			RECT	129.377 10.028 129.409 10.092 ;
			RECT	129.545 10.028 129.577 10.092 ;
			RECT	129.713 10.028 129.745 10.092 ;
			RECT	129.881 10.028 129.913 10.092 ;
			RECT	130.049 10.028 130.081 10.092 ;
			RECT	130.217 10.028 130.249 10.092 ;
			RECT	130.385 10.028 130.417 10.092 ;
			RECT	130.553 10.028 130.585 10.092 ;
			RECT	130.721 10.028 130.753 10.092 ;
			RECT	130.889 10.028 130.921 10.092 ;
			RECT	131.057 10.028 131.089 10.092 ;
			RECT	131.225 10.028 131.257 10.092 ;
			RECT	131.393 10.028 131.425 10.092 ;
			RECT	131.561 10.028 131.593 10.092 ;
			RECT	131.729 10.028 131.761 10.092 ;
			RECT	131.897 10.028 131.929 10.092 ;
			RECT	132.065 10.028 132.097 10.092 ;
			RECT	132.233 10.028 132.265 10.092 ;
			RECT	132.401 10.028 132.433 10.092 ;
			RECT	132.569 10.028 132.601 10.092 ;
			RECT	132.737 10.028 132.769 10.092 ;
			RECT	132.905 10.028 132.937 10.092 ;
			RECT	133.073 10.028 133.105 10.092 ;
			RECT	133.241 10.028 133.273 10.092 ;
			RECT	133.409 10.028 133.441 10.092 ;
			RECT	133.577 10.028 133.609 10.092 ;
			RECT	133.745 10.028 133.777 10.092 ;
			RECT	133.913 10.028 133.945 10.092 ;
			RECT	134.081 10.028 134.113 10.092 ;
			RECT	134.249 10.028 134.281 10.092 ;
			RECT	134.417 10.028 134.449 10.092 ;
			RECT	134.585 10.028 134.617 10.092 ;
			RECT	134.753 10.028 134.785 10.092 ;
			RECT	134.921 10.028 134.953 10.092 ;
			RECT	135.089 10.028 135.121 10.092 ;
			RECT	135.257 10.028 135.289 10.092 ;
			RECT	135.425 10.028 135.457 10.092 ;
			RECT	135.593 10.028 135.625 10.092 ;
			RECT	135.761 10.028 135.793 10.092 ;
			RECT	135.929 10.028 135.961 10.092 ;
			RECT	136.097 10.028 136.129 10.092 ;
			RECT	136.265 10.028 136.297 10.092 ;
			RECT	136.433 10.028 136.465 10.092 ;
			RECT	136.601 10.028 136.633 10.092 ;
			RECT	136.769 10.028 136.801 10.092 ;
			RECT	136.937 10.028 136.969 10.092 ;
			RECT	137.105 10.028 137.137 10.092 ;
			RECT	137.273 10.028 137.305 10.092 ;
			RECT	137.441 10.028 137.473 10.092 ;
			RECT	137.609 10.028 137.641 10.092 ;
			RECT	137.777 10.028 137.809 10.092 ;
			RECT	137.945 10.028 137.977 10.092 ;
			RECT	138.113 10.028 138.145 10.092 ;
			RECT	138.281 10.028 138.313 10.092 ;
			RECT	138.449 10.028 138.481 10.092 ;
			RECT	138.617 10.028 138.649 10.092 ;
			RECT	138.785 10.028 138.817 10.092 ;
			RECT	138.953 10.028 138.985 10.092 ;
			RECT	139.121 10.028 139.153 10.092 ;
			RECT	139.289 10.028 139.321 10.092 ;
			RECT	139.457 10.028 139.489 10.092 ;
			RECT	139.625 10.028 139.657 10.092 ;
			RECT	139.793 10.028 139.825 10.092 ;
			RECT	139.961 10.028 139.993 10.092 ;
			RECT	140.129 10.028 140.161 10.092 ;
			RECT	140.297 10.028 140.329 10.092 ;
			RECT	140.465 10.028 140.497 10.092 ;
			RECT	140.633 10.028 140.665 10.092 ;
			RECT	140.801 10.028 140.833 10.092 ;
			RECT	140.969 10.028 141.001 10.092 ;
			RECT	141.137 10.028 141.169 10.092 ;
			RECT	141.305 10.028 141.337 10.092 ;
			RECT	141.473 10.028 141.505 10.092 ;
			RECT	141.641 10.028 141.673 10.092 ;
			RECT	141.809 10.028 141.841 10.092 ;
			RECT	141.977 10.028 142.009 10.092 ;
			RECT	142.145 10.028 142.177 10.092 ;
			RECT	142.313 10.028 142.345 10.092 ;
			RECT	142.481 10.028 142.513 10.092 ;
			RECT	142.649 10.028 142.681 10.092 ;
			RECT	142.817 10.028 142.849 10.092 ;
			RECT	142.985 10.028 143.017 10.092 ;
			RECT	143.153 10.028 143.185 10.092 ;
			RECT	143.321 10.028 143.353 10.092 ;
			RECT	143.489 10.028 143.521 10.092 ;
			RECT	143.657 10.028 143.689 10.092 ;
			RECT	143.825 10.028 143.857 10.092 ;
			RECT	143.993 10.028 144.025 10.092 ;
			RECT	144.161 10.028 144.193 10.092 ;
			RECT	144.329 10.028 144.361 10.092 ;
			RECT	144.497 10.028 144.529 10.092 ;
			RECT	144.665 10.028 144.697 10.092 ;
			RECT	144.833 10.028 144.865 10.092 ;
			RECT	145.001 10.028 145.033 10.092 ;
			RECT	145.169 10.028 145.201 10.092 ;
			RECT	145.337 10.028 145.369 10.092 ;
			RECT	145.505 10.028 145.537 10.092 ;
			RECT	145.673 10.028 145.705 10.092 ;
			RECT	145.841 10.028 145.873 10.092 ;
			RECT	146.009 10.028 146.041 10.092 ;
			RECT	146.177 10.028 146.209 10.092 ;
			RECT	146.345 10.028 146.377 10.092 ;
			RECT	146.513 10.028 146.545 10.092 ;
			RECT	146.681 10.028 146.713 10.092 ;
			RECT	146.849 10.028 146.881 10.092 ;
			RECT	147.017 10.028 147.049 10.092 ;
			RECT	147.185 10.028 147.217 10.092 ;
			RECT	147.316 10.044 147.348 10.076 ;
			RECT	147.437 10.044 147.469 10.076 ;
			RECT	147.567 10.028 147.599 10.092 ;
			RECT	149.879 10.028 149.911 10.092 ;
			RECT	151.13 10.028 151.194 10.092 ;
			RECT	151.81 10.028 151.842 10.092 ;
			RECT	152.249 10.028 152.281 10.092 ;
			RECT	153.56 10.028 153.624 10.092 ;
			RECT	156.601 10.028 156.633 10.092 ;
			RECT	156.731 10.044 156.763 10.076 ;
			RECT	156.852 10.044 156.884 10.076 ;
			RECT	156.983 10.028 157.015 10.092 ;
			RECT	157.151 10.028 157.183 10.092 ;
			RECT	157.319 10.028 157.351 10.092 ;
			RECT	157.487 10.028 157.519 10.092 ;
			RECT	157.655 10.028 157.687 10.092 ;
			RECT	157.823 10.028 157.855 10.092 ;
			RECT	157.991 10.028 158.023 10.092 ;
			RECT	158.159 10.028 158.191 10.092 ;
			RECT	158.327 10.028 158.359 10.092 ;
			RECT	158.495 10.028 158.527 10.092 ;
			RECT	158.663 10.028 158.695 10.092 ;
			RECT	158.831 10.028 158.863 10.092 ;
			RECT	158.999 10.028 159.031 10.092 ;
			RECT	159.167 10.028 159.199 10.092 ;
			RECT	159.335 10.028 159.367 10.092 ;
			RECT	159.503 10.028 159.535 10.092 ;
			RECT	159.671 10.028 159.703 10.092 ;
			RECT	159.839 10.028 159.871 10.092 ;
			RECT	160.007 10.028 160.039 10.092 ;
			RECT	160.175 10.028 160.207 10.092 ;
			RECT	160.343 10.028 160.375 10.092 ;
			RECT	160.511 10.028 160.543 10.092 ;
			RECT	160.679 10.028 160.711 10.092 ;
			RECT	160.847 10.028 160.879 10.092 ;
			RECT	161.015 10.028 161.047 10.092 ;
			RECT	161.183 10.028 161.215 10.092 ;
			RECT	161.351 10.028 161.383 10.092 ;
			RECT	161.519 10.028 161.551 10.092 ;
			RECT	161.687 10.028 161.719 10.092 ;
			RECT	161.855 10.028 161.887 10.092 ;
			RECT	162.023 10.028 162.055 10.092 ;
			RECT	162.191 10.028 162.223 10.092 ;
			RECT	162.359 10.028 162.391 10.092 ;
			RECT	162.527 10.028 162.559 10.092 ;
			RECT	162.695 10.028 162.727 10.092 ;
			RECT	162.863 10.028 162.895 10.092 ;
			RECT	163.031 10.028 163.063 10.092 ;
			RECT	163.199 10.028 163.231 10.092 ;
			RECT	163.367 10.028 163.399 10.092 ;
			RECT	163.535 10.028 163.567 10.092 ;
			RECT	163.703 10.028 163.735 10.092 ;
			RECT	163.871 10.028 163.903 10.092 ;
			RECT	164.039 10.028 164.071 10.092 ;
			RECT	164.207 10.028 164.239 10.092 ;
			RECT	164.375 10.028 164.407 10.092 ;
			RECT	164.543 10.028 164.575 10.092 ;
			RECT	164.711 10.028 164.743 10.092 ;
			RECT	164.879 10.028 164.911 10.092 ;
			RECT	165.047 10.028 165.079 10.092 ;
			RECT	165.215 10.028 165.247 10.092 ;
			RECT	165.383 10.028 165.415 10.092 ;
			RECT	165.551 10.028 165.583 10.092 ;
			RECT	165.719 10.028 165.751 10.092 ;
			RECT	165.887 10.028 165.919 10.092 ;
			RECT	166.055 10.028 166.087 10.092 ;
			RECT	166.223 10.028 166.255 10.092 ;
			RECT	166.391 10.028 166.423 10.092 ;
			RECT	166.559 10.028 166.591 10.092 ;
			RECT	166.727 10.028 166.759 10.092 ;
			RECT	166.895 10.028 166.927 10.092 ;
			RECT	167.063 10.028 167.095 10.092 ;
			RECT	167.231 10.028 167.263 10.092 ;
			RECT	167.399 10.028 167.431 10.092 ;
			RECT	167.567 10.028 167.599 10.092 ;
			RECT	167.735 10.028 167.767 10.092 ;
			RECT	167.903 10.028 167.935 10.092 ;
			RECT	168.071 10.028 168.103 10.092 ;
			RECT	168.239 10.028 168.271 10.092 ;
			RECT	168.407 10.028 168.439 10.092 ;
			RECT	168.575 10.028 168.607 10.092 ;
			RECT	168.743 10.028 168.775 10.092 ;
			RECT	168.911 10.028 168.943 10.092 ;
			RECT	169.079 10.028 169.111 10.092 ;
			RECT	169.247 10.028 169.279 10.092 ;
			RECT	169.415 10.028 169.447 10.092 ;
			RECT	169.583 10.028 169.615 10.092 ;
			RECT	169.751 10.028 169.783 10.092 ;
			RECT	169.919 10.028 169.951 10.092 ;
			RECT	170.087 10.028 170.119 10.092 ;
			RECT	170.255 10.028 170.287 10.092 ;
			RECT	170.423 10.028 170.455 10.092 ;
			RECT	170.591 10.028 170.623 10.092 ;
			RECT	170.759 10.028 170.791 10.092 ;
			RECT	170.927 10.028 170.959 10.092 ;
			RECT	171.095 10.028 171.127 10.092 ;
			RECT	171.263 10.028 171.295 10.092 ;
			RECT	171.431 10.028 171.463 10.092 ;
			RECT	171.599 10.028 171.631 10.092 ;
			RECT	171.767 10.028 171.799 10.092 ;
			RECT	171.935 10.028 171.967 10.092 ;
			RECT	172.103 10.028 172.135 10.092 ;
			RECT	172.271 10.028 172.303 10.092 ;
			RECT	172.439 10.028 172.471 10.092 ;
			RECT	172.607 10.028 172.639 10.092 ;
			RECT	172.775 10.028 172.807 10.092 ;
			RECT	172.943 10.028 172.975 10.092 ;
			RECT	173.111 10.028 173.143 10.092 ;
			RECT	173.279 10.028 173.311 10.092 ;
			RECT	173.447 10.028 173.479 10.092 ;
			RECT	173.615 10.028 173.647 10.092 ;
			RECT	173.783 10.028 173.815 10.092 ;
			RECT	173.951 10.028 173.983 10.092 ;
			RECT	174.119 10.028 174.151 10.092 ;
			RECT	174.287 10.028 174.319 10.092 ;
			RECT	174.455 10.028 174.487 10.092 ;
			RECT	174.623 10.028 174.655 10.092 ;
			RECT	174.791 10.028 174.823 10.092 ;
			RECT	174.959 10.028 174.991 10.092 ;
			RECT	175.127 10.028 175.159 10.092 ;
			RECT	175.295 10.028 175.327 10.092 ;
			RECT	175.463 10.028 175.495 10.092 ;
			RECT	175.631 10.028 175.663 10.092 ;
			RECT	175.799 10.028 175.831 10.092 ;
			RECT	175.967 10.028 175.999 10.092 ;
			RECT	176.135 10.028 176.167 10.092 ;
			RECT	176.303 10.028 176.335 10.092 ;
			RECT	176.471 10.028 176.503 10.092 ;
			RECT	176.639 10.028 176.671 10.092 ;
			RECT	176.807 10.028 176.839 10.092 ;
			RECT	176.975 10.028 177.007 10.092 ;
			RECT	177.143 10.028 177.175 10.092 ;
			RECT	177.311 10.028 177.343 10.092 ;
			RECT	177.479 10.028 177.511 10.092 ;
			RECT	177.647 10.028 177.679 10.092 ;
			RECT	177.815 10.028 177.847 10.092 ;
			RECT	177.983 10.028 178.015 10.092 ;
			RECT	178.151 10.028 178.183 10.092 ;
			RECT	178.319 10.028 178.351 10.092 ;
			RECT	178.487 10.028 178.519 10.092 ;
			RECT	178.655 10.028 178.687 10.092 ;
			RECT	178.823 10.028 178.855 10.092 ;
			RECT	178.991 10.028 179.023 10.092 ;
			RECT	179.159 10.028 179.191 10.092 ;
			RECT	179.327 10.028 179.359 10.092 ;
			RECT	179.495 10.028 179.527 10.092 ;
			RECT	179.663 10.028 179.695 10.092 ;
			RECT	179.831 10.028 179.863 10.092 ;
			RECT	179.999 10.028 180.031 10.092 ;
			RECT	180.167 10.028 180.199 10.092 ;
			RECT	180.335 10.028 180.367 10.092 ;
			RECT	180.503 10.028 180.535 10.092 ;
			RECT	180.671 10.028 180.703 10.092 ;
			RECT	180.839 10.028 180.871 10.092 ;
			RECT	181.007 10.028 181.039 10.092 ;
			RECT	181.175 10.028 181.207 10.092 ;
			RECT	181.343 10.028 181.375 10.092 ;
			RECT	181.511 10.028 181.543 10.092 ;
			RECT	181.679 10.028 181.711 10.092 ;
			RECT	181.847 10.028 181.879 10.092 ;
			RECT	182.015 10.028 182.047 10.092 ;
			RECT	182.183 10.028 182.215 10.092 ;
			RECT	182.351 10.028 182.383 10.092 ;
			RECT	182.519 10.028 182.551 10.092 ;
			RECT	182.687 10.028 182.719 10.092 ;
			RECT	182.855 10.028 182.887 10.092 ;
			RECT	183.023 10.028 183.055 10.092 ;
			RECT	183.191 10.028 183.223 10.092 ;
			RECT	183.359 10.028 183.391 10.092 ;
			RECT	183.527 10.028 183.559 10.092 ;
			RECT	183.695 10.028 183.727 10.092 ;
			RECT	183.863 10.028 183.895 10.092 ;
			RECT	184.031 10.028 184.063 10.092 ;
			RECT	184.199 10.028 184.231 10.092 ;
			RECT	184.367 10.028 184.399 10.092 ;
			RECT	184.535 10.028 184.567 10.092 ;
			RECT	184.703 10.028 184.735 10.092 ;
			RECT	184.871 10.028 184.903 10.092 ;
			RECT	185.039 10.028 185.071 10.092 ;
			RECT	185.207 10.028 185.239 10.092 ;
			RECT	185.375 10.028 185.407 10.092 ;
			RECT	185.543 10.028 185.575 10.092 ;
			RECT	185.711 10.028 185.743 10.092 ;
			RECT	185.879 10.028 185.911 10.092 ;
			RECT	186.047 10.028 186.079 10.092 ;
			RECT	186.215 10.028 186.247 10.092 ;
			RECT	186.383 10.028 186.415 10.092 ;
			RECT	186.551 10.028 186.583 10.092 ;
			RECT	186.719 10.028 186.751 10.092 ;
			RECT	186.887 10.028 186.919 10.092 ;
			RECT	187.055 10.028 187.087 10.092 ;
			RECT	187.223 10.028 187.255 10.092 ;
			RECT	187.391 10.028 187.423 10.092 ;
			RECT	187.559 10.028 187.591 10.092 ;
			RECT	187.727 10.028 187.759 10.092 ;
			RECT	187.895 10.028 187.927 10.092 ;
			RECT	188.063 10.028 188.095 10.092 ;
			RECT	188.231 10.028 188.263 10.092 ;
			RECT	188.399 10.028 188.431 10.092 ;
			RECT	188.567 10.028 188.599 10.092 ;
			RECT	188.735 10.028 188.767 10.092 ;
			RECT	188.903 10.028 188.935 10.092 ;
			RECT	189.071 10.028 189.103 10.092 ;
			RECT	189.239 10.028 189.271 10.092 ;
			RECT	189.407 10.028 189.439 10.092 ;
			RECT	189.575 10.028 189.607 10.092 ;
			RECT	189.743 10.028 189.775 10.092 ;
			RECT	189.911 10.028 189.943 10.092 ;
			RECT	190.079 10.028 190.111 10.092 ;
			RECT	190.247 10.028 190.279 10.092 ;
			RECT	190.415 10.028 190.447 10.092 ;
			RECT	190.583 10.028 190.615 10.092 ;
			RECT	190.751 10.028 190.783 10.092 ;
			RECT	190.919 10.028 190.951 10.092 ;
			RECT	191.087 10.028 191.119 10.092 ;
			RECT	191.255 10.028 191.287 10.092 ;
			RECT	191.423 10.028 191.455 10.092 ;
			RECT	191.591 10.028 191.623 10.092 ;
			RECT	191.759 10.028 191.791 10.092 ;
			RECT	191.927 10.028 191.959 10.092 ;
			RECT	192.095 10.028 192.127 10.092 ;
			RECT	192.263 10.028 192.295 10.092 ;
			RECT	192.431 10.028 192.463 10.092 ;
			RECT	192.599 10.028 192.631 10.092 ;
			RECT	192.767 10.028 192.799 10.092 ;
			RECT	192.935 10.028 192.967 10.092 ;
			RECT	193.103 10.028 193.135 10.092 ;
			RECT	193.271 10.028 193.303 10.092 ;
			RECT	193.439 10.028 193.471 10.092 ;
			RECT	193.607 10.028 193.639 10.092 ;
			RECT	193.775 10.028 193.807 10.092 ;
			RECT	193.943 10.028 193.975 10.092 ;
			RECT	194.111 10.028 194.143 10.092 ;
			RECT	194.279 10.028 194.311 10.092 ;
			RECT	194.447 10.028 194.479 10.092 ;
			RECT	194.615 10.028 194.647 10.092 ;
			RECT	194.783 10.028 194.815 10.092 ;
			RECT	194.951 10.028 194.983 10.092 ;
			RECT	195.119 10.028 195.151 10.092 ;
			RECT	195.287 10.028 195.319 10.092 ;
			RECT	195.455 10.028 195.487 10.092 ;
			RECT	195.623 10.028 195.655 10.092 ;
			RECT	195.791 10.028 195.823 10.092 ;
			RECT	195.959 10.028 195.991 10.092 ;
			RECT	196.127 10.028 196.159 10.092 ;
			RECT	196.295 10.028 196.327 10.092 ;
			RECT	196.463 10.028 196.495 10.092 ;
			RECT	196.631 10.028 196.663 10.092 ;
			RECT	196.799 10.028 196.831 10.092 ;
			RECT	196.967 10.028 196.999 10.092 ;
			RECT	197.135 10.028 197.167 10.092 ;
			RECT	197.303 10.028 197.335 10.092 ;
			RECT	197.471 10.028 197.503 10.092 ;
			RECT	197.639 10.028 197.671 10.092 ;
			RECT	197.807 10.028 197.839 10.092 ;
			RECT	197.975 10.028 198.007 10.092 ;
			RECT	198.143 10.028 198.175 10.092 ;
			RECT	198.311 10.028 198.343 10.092 ;
			RECT	198.479 10.028 198.511 10.092 ;
			RECT	198.647 10.028 198.679 10.092 ;
			RECT	198.815 10.028 198.847 10.092 ;
			RECT	198.983 10.028 199.015 10.092 ;
			RECT	199.151 10.028 199.183 10.092 ;
			RECT	199.319 10.028 199.351 10.092 ;
			RECT	199.487 10.028 199.519 10.092 ;
			RECT	199.655 10.028 199.687 10.092 ;
			RECT	199.823 10.028 199.855 10.092 ;
			RECT	199.991 10.028 200.023 10.092 ;
			RECT	200.121 10.044 200.153 10.076 ;
			RECT	200.243 10.049 200.275 10.081 ;
			RECT	200.373 10.028 200.405 10.092 ;
			RECT	200.9 10.028 200.932 10.092 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 73.976 201.665 74.096 ;
			LAYER	J3 ;
			RECT	0.755 74.004 0.787 74.068 ;
			RECT	1.645 74.004 1.709 74.068 ;
			RECT	2.323 74.004 2.387 74.068 ;
			RECT	3.438 74.004 3.47 74.068 ;
			RECT	3.585 74.004 3.617 74.068 ;
			RECT	4.195 74.004 4.227 74.068 ;
			RECT	4.72 74.004 4.752 74.068 ;
			RECT	4.944 74.004 5.008 74.068 ;
			RECT	5.267 74.004 5.299 74.068 ;
			RECT	5.797 74.004 5.829 74.068 ;
			RECT	5.927 74.015 5.959 74.047 ;
			RECT	6.049 74.02 6.081 74.052 ;
			RECT	6.179 74.004 6.211 74.068 ;
			RECT	6.347 74.004 6.379 74.068 ;
			RECT	6.515 74.004 6.547 74.068 ;
			RECT	6.683 74.004 6.715 74.068 ;
			RECT	6.851 74.004 6.883 74.068 ;
			RECT	7.019 74.004 7.051 74.068 ;
			RECT	7.187 74.004 7.219 74.068 ;
			RECT	7.355 74.004 7.387 74.068 ;
			RECT	7.523 74.004 7.555 74.068 ;
			RECT	7.691 74.004 7.723 74.068 ;
			RECT	7.859 74.004 7.891 74.068 ;
			RECT	8.027 74.004 8.059 74.068 ;
			RECT	8.195 74.004 8.227 74.068 ;
			RECT	8.363 74.004 8.395 74.068 ;
			RECT	8.531 74.004 8.563 74.068 ;
			RECT	8.699 74.004 8.731 74.068 ;
			RECT	8.867 74.004 8.899 74.068 ;
			RECT	9.035 74.004 9.067 74.068 ;
			RECT	9.203 74.004 9.235 74.068 ;
			RECT	9.371 74.004 9.403 74.068 ;
			RECT	9.539 74.004 9.571 74.068 ;
			RECT	9.707 74.004 9.739 74.068 ;
			RECT	9.875 74.004 9.907 74.068 ;
			RECT	10.043 74.004 10.075 74.068 ;
			RECT	10.211 74.004 10.243 74.068 ;
			RECT	10.379 74.004 10.411 74.068 ;
			RECT	10.547 74.004 10.579 74.068 ;
			RECT	10.715 74.004 10.747 74.068 ;
			RECT	10.883 74.004 10.915 74.068 ;
			RECT	11.051 74.004 11.083 74.068 ;
			RECT	11.219 74.004 11.251 74.068 ;
			RECT	11.387 74.004 11.419 74.068 ;
			RECT	11.555 74.004 11.587 74.068 ;
			RECT	11.723 74.004 11.755 74.068 ;
			RECT	11.891 74.004 11.923 74.068 ;
			RECT	12.059 74.004 12.091 74.068 ;
			RECT	12.227 74.004 12.259 74.068 ;
			RECT	12.395 74.004 12.427 74.068 ;
			RECT	12.563 74.004 12.595 74.068 ;
			RECT	12.731 74.004 12.763 74.068 ;
			RECT	12.899 74.004 12.931 74.068 ;
			RECT	13.067 74.004 13.099 74.068 ;
			RECT	13.235 74.004 13.267 74.068 ;
			RECT	13.403 74.004 13.435 74.068 ;
			RECT	13.571 74.004 13.603 74.068 ;
			RECT	13.739 74.004 13.771 74.068 ;
			RECT	13.907 74.004 13.939 74.068 ;
			RECT	14.075 74.004 14.107 74.068 ;
			RECT	14.243 74.004 14.275 74.068 ;
			RECT	14.411 74.004 14.443 74.068 ;
			RECT	14.579 74.004 14.611 74.068 ;
			RECT	14.747 74.004 14.779 74.068 ;
			RECT	14.915 74.004 14.947 74.068 ;
			RECT	15.083 74.004 15.115 74.068 ;
			RECT	15.251 74.004 15.283 74.068 ;
			RECT	15.419 74.004 15.451 74.068 ;
			RECT	15.587 74.004 15.619 74.068 ;
			RECT	15.755 74.004 15.787 74.068 ;
			RECT	15.923 74.004 15.955 74.068 ;
			RECT	16.091 74.004 16.123 74.068 ;
			RECT	16.259 74.004 16.291 74.068 ;
			RECT	16.427 74.004 16.459 74.068 ;
			RECT	16.595 74.004 16.627 74.068 ;
			RECT	16.763 74.004 16.795 74.068 ;
			RECT	16.931 74.004 16.963 74.068 ;
			RECT	17.099 74.004 17.131 74.068 ;
			RECT	17.267 74.004 17.299 74.068 ;
			RECT	17.435 74.004 17.467 74.068 ;
			RECT	17.603 74.004 17.635 74.068 ;
			RECT	17.771 74.004 17.803 74.068 ;
			RECT	17.939 74.004 17.971 74.068 ;
			RECT	18.107 74.004 18.139 74.068 ;
			RECT	18.275 74.004 18.307 74.068 ;
			RECT	18.443 74.004 18.475 74.068 ;
			RECT	18.611 74.004 18.643 74.068 ;
			RECT	18.779 74.004 18.811 74.068 ;
			RECT	18.947 74.004 18.979 74.068 ;
			RECT	19.115 74.004 19.147 74.068 ;
			RECT	19.283 74.004 19.315 74.068 ;
			RECT	19.451 74.004 19.483 74.068 ;
			RECT	19.619 74.004 19.651 74.068 ;
			RECT	19.787 74.004 19.819 74.068 ;
			RECT	19.955 74.004 19.987 74.068 ;
			RECT	20.123 74.004 20.155 74.068 ;
			RECT	20.291 74.004 20.323 74.068 ;
			RECT	20.459 74.004 20.491 74.068 ;
			RECT	20.627 74.004 20.659 74.068 ;
			RECT	20.795 74.004 20.827 74.068 ;
			RECT	20.963 74.004 20.995 74.068 ;
			RECT	21.131 74.004 21.163 74.068 ;
			RECT	21.299 74.004 21.331 74.068 ;
			RECT	21.467 74.004 21.499 74.068 ;
			RECT	21.635 74.004 21.667 74.068 ;
			RECT	21.803 74.004 21.835 74.068 ;
			RECT	21.971 74.004 22.003 74.068 ;
			RECT	22.139 74.004 22.171 74.068 ;
			RECT	22.307 74.004 22.339 74.068 ;
			RECT	22.475 74.004 22.507 74.068 ;
			RECT	22.643 74.004 22.675 74.068 ;
			RECT	22.811 74.004 22.843 74.068 ;
			RECT	22.979 74.004 23.011 74.068 ;
			RECT	23.147 74.004 23.179 74.068 ;
			RECT	23.315 74.004 23.347 74.068 ;
			RECT	23.483 74.004 23.515 74.068 ;
			RECT	23.651 74.004 23.683 74.068 ;
			RECT	23.819 74.004 23.851 74.068 ;
			RECT	23.987 74.004 24.019 74.068 ;
			RECT	24.155 74.004 24.187 74.068 ;
			RECT	24.323 74.004 24.355 74.068 ;
			RECT	24.491 74.004 24.523 74.068 ;
			RECT	24.659 74.004 24.691 74.068 ;
			RECT	24.827 74.004 24.859 74.068 ;
			RECT	24.995 74.004 25.027 74.068 ;
			RECT	25.163 74.004 25.195 74.068 ;
			RECT	25.331 74.004 25.363 74.068 ;
			RECT	25.499 74.004 25.531 74.068 ;
			RECT	25.667 74.004 25.699 74.068 ;
			RECT	25.835 74.004 25.867 74.068 ;
			RECT	26.003 74.004 26.035 74.068 ;
			RECT	26.171 74.004 26.203 74.068 ;
			RECT	26.339 74.004 26.371 74.068 ;
			RECT	26.507 74.004 26.539 74.068 ;
			RECT	26.675 74.004 26.707 74.068 ;
			RECT	26.843 74.004 26.875 74.068 ;
			RECT	27.011 74.004 27.043 74.068 ;
			RECT	27.179 74.004 27.211 74.068 ;
			RECT	27.347 74.004 27.379 74.068 ;
			RECT	27.515 74.004 27.547 74.068 ;
			RECT	27.683 74.004 27.715 74.068 ;
			RECT	27.851 74.004 27.883 74.068 ;
			RECT	28.019 74.004 28.051 74.068 ;
			RECT	28.187 74.004 28.219 74.068 ;
			RECT	28.355 74.004 28.387 74.068 ;
			RECT	28.523 74.004 28.555 74.068 ;
			RECT	28.691 74.004 28.723 74.068 ;
			RECT	28.859 74.004 28.891 74.068 ;
			RECT	29.027 74.004 29.059 74.068 ;
			RECT	29.195 74.004 29.227 74.068 ;
			RECT	29.363 74.004 29.395 74.068 ;
			RECT	29.531 74.004 29.563 74.068 ;
			RECT	29.699 74.004 29.731 74.068 ;
			RECT	29.867 74.004 29.899 74.068 ;
			RECT	30.035 74.004 30.067 74.068 ;
			RECT	30.203 74.004 30.235 74.068 ;
			RECT	30.371 74.004 30.403 74.068 ;
			RECT	30.539 74.004 30.571 74.068 ;
			RECT	30.707 74.004 30.739 74.068 ;
			RECT	30.875 74.004 30.907 74.068 ;
			RECT	31.043 74.004 31.075 74.068 ;
			RECT	31.211 74.004 31.243 74.068 ;
			RECT	31.379 74.004 31.411 74.068 ;
			RECT	31.547 74.004 31.579 74.068 ;
			RECT	31.715 74.004 31.747 74.068 ;
			RECT	31.883 74.004 31.915 74.068 ;
			RECT	32.051 74.004 32.083 74.068 ;
			RECT	32.219 74.004 32.251 74.068 ;
			RECT	32.387 74.004 32.419 74.068 ;
			RECT	32.555 74.004 32.587 74.068 ;
			RECT	32.723 74.004 32.755 74.068 ;
			RECT	32.891 74.004 32.923 74.068 ;
			RECT	33.059 74.004 33.091 74.068 ;
			RECT	33.227 74.004 33.259 74.068 ;
			RECT	33.395 74.004 33.427 74.068 ;
			RECT	33.563 74.004 33.595 74.068 ;
			RECT	33.731 74.004 33.763 74.068 ;
			RECT	33.899 74.004 33.931 74.068 ;
			RECT	34.067 74.004 34.099 74.068 ;
			RECT	34.235 74.004 34.267 74.068 ;
			RECT	34.403 74.004 34.435 74.068 ;
			RECT	34.571 74.004 34.603 74.068 ;
			RECT	34.739 74.004 34.771 74.068 ;
			RECT	34.907 74.004 34.939 74.068 ;
			RECT	35.075 74.004 35.107 74.068 ;
			RECT	35.243 74.004 35.275 74.068 ;
			RECT	35.411 74.004 35.443 74.068 ;
			RECT	35.579 74.004 35.611 74.068 ;
			RECT	35.747 74.004 35.779 74.068 ;
			RECT	35.915 74.004 35.947 74.068 ;
			RECT	36.083 74.004 36.115 74.068 ;
			RECT	36.251 74.004 36.283 74.068 ;
			RECT	36.419 74.004 36.451 74.068 ;
			RECT	36.587 74.004 36.619 74.068 ;
			RECT	36.755 74.004 36.787 74.068 ;
			RECT	36.923 74.004 36.955 74.068 ;
			RECT	37.091 74.004 37.123 74.068 ;
			RECT	37.259 74.004 37.291 74.068 ;
			RECT	37.427 74.004 37.459 74.068 ;
			RECT	37.595 74.004 37.627 74.068 ;
			RECT	37.763 74.004 37.795 74.068 ;
			RECT	37.931 74.004 37.963 74.068 ;
			RECT	38.099 74.004 38.131 74.068 ;
			RECT	38.267 74.004 38.299 74.068 ;
			RECT	38.435 74.004 38.467 74.068 ;
			RECT	38.603 74.004 38.635 74.068 ;
			RECT	38.771 74.004 38.803 74.068 ;
			RECT	38.939 74.004 38.971 74.068 ;
			RECT	39.107 74.004 39.139 74.068 ;
			RECT	39.275 74.004 39.307 74.068 ;
			RECT	39.443 74.004 39.475 74.068 ;
			RECT	39.611 74.004 39.643 74.068 ;
			RECT	39.779 74.004 39.811 74.068 ;
			RECT	39.947 74.004 39.979 74.068 ;
			RECT	40.115 74.004 40.147 74.068 ;
			RECT	40.283 74.004 40.315 74.068 ;
			RECT	40.451 74.004 40.483 74.068 ;
			RECT	40.619 74.004 40.651 74.068 ;
			RECT	40.787 74.004 40.819 74.068 ;
			RECT	40.955 74.004 40.987 74.068 ;
			RECT	41.123 74.004 41.155 74.068 ;
			RECT	41.291 74.004 41.323 74.068 ;
			RECT	41.459 74.004 41.491 74.068 ;
			RECT	41.627 74.004 41.659 74.068 ;
			RECT	41.795 74.004 41.827 74.068 ;
			RECT	41.963 74.004 41.995 74.068 ;
			RECT	42.131 74.004 42.163 74.068 ;
			RECT	42.299 74.004 42.331 74.068 ;
			RECT	42.467 74.004 42.499 74.068 ;
			RECT	42.635 74.004 42.667 74.068 ;
			RECT	42.803 74.004 42.835 74.068 ;
			RECT	42.971 74.004 43.003 74.068 ;
			RECT	43.139 74.004 43.171 74.068 ;
			RECT	43.307 74.004 43.339 74.068 ;
			RECT	43.475 74.004 43.507 74.068 ;
			RECT	43.643 74.004 43.675 74.068 ;
			RECT	43.811 74.004 43.843 74.068 ;
			RECT	43.979 74.004 44.011 74.068 ;
			RECT	44.147 74.004 44.179 74.068 ;
			RECT	44.315 74.004 44.347 74.068 ;
			RECT	44.483 74.004 44.515 74.068 ;
			RECT	44.651 74.004 44.683 74.068 ;
			RECT	44.819 74.004 44.851 74.068 ;
			RECT	44.987 74.004 45.019 74.068 ;
			RECT	45.155 74.004 45.187 74.068 ;
			RECT	45.323 74.004 45.355 74.068 ;
			RECT	45.491 74.004 45.523 74.068 ;
			RECT	45.659 74.004 45.691 74.068 ;
			RECT	45.827 74.004 45.859 74.068 ;
			RECT	45.995 74.004 46.027 74.068 ;
			RECT	46.163 74.004 46.195 74.068 ;
			RECT	46.331 74.004 46.363 74.068 ;
			RECT	46.499 74.004 46.531 74.068 ;
			RECT	46.667 74.004 46.699 74.068 ;
			RECT	46.835 74.004 46.867 74.068 ;
			RECT	47.003 74.004 47.035 74.068 ;
			RECT	47.171 74.004 47.203 74.068 ;
			RECT	47.339 74.004 47.371 74.068 ;
			RECT	47.507 74.004 47.539 74.068 ;
			RECT	47.675 74.004 47.707 74.068 ;
			RECT	47.843 74.004 47.875 74.068 ;
			RECT	48.011 74.004 48.043 74.068 ;
			RECT	48.179 74.004 48.211 74.068 ;
			RECT	48.347 74.004 48.379 74.068 ;
			RECT	48.515 74.004 48.547 74.068 ;
			RECT	48.683 74.004 48.715 74.068 ;
			RECT	48.851 74.004 48.883 74.068 ;
			RECT	49.019 74.004 49.051 74.068 ;
			RECT	49.187 74.004 49.219 74.068 ;
			RECT	49.318 74.02 49.35 74.052 ;
			RECT	49.439 74.02 49.471 74.052 ;
			RECT	49.569 74.004 49.601 74.068 ;
			RECT	51.881 74.004 51.913 74.068 ;
			RECT	53.132 74.004 53.196 74.068 ;
			RECT	53.812 74.004 53.844 74.068 ;
			RECT	54.251 74.004 54.283 74.068 ;
			RECT	55.562 74.004 55.626 74.068 ;
			RECT	58.603 74.004 58.635 74.068 ;
			RECT	58.733 74.02 58.765 74.052 ;
			RECT	58.854 74.02 58.886 74.052 ;
			RECT	58.985 74.004 59.017 74.068 ;
			RECT	59.153 74.004 59.185 74.068 ;
			RECT	59.321 74.004 59.353 74.068 ;
			RECT	59.489 74.004 59.521 74.068 ;
			RECT	59.657 74.004 59.689 74.068 ;
			RECT	59.825 74.004 59.857 74.068 ;
			RECT	59.993 74.004 60.025 74.068 ;
			RECT	60.161 74.004 60.193 74.068 ;
			RECT	60.329 74.004 60.361 74.068 ;
			RECT	60.497 74.004 60.529 74.068 ;
			RECT	60.665 74.004 60.697 74.068 ;
			RECT	60.833 74.004 60.865 74.068 ;
			RECT	61.001 74.004 61.033 74.068 ;
			RECT	61.169 74.004 61.201 74.068 ;
			RECT	61.337 74.004 61.369 74.068 ;
			RECT	61.505 74.004 61.537 74.068 ;
			RECT	61.673 74.004 61.705 74.068 ;
			RECT	61.841 74.004 61.873 74.068 ;
			RECT	62.009 74.004 62.041 74.068 ;
			RECT	62.177 74.004 62.209 74.068 ;
			RECT	62.345 74.004 62.377 74.068 ;
			RECT	62.513 74.004 62.545 74.068 ;
			RECT	62.681 74.004 62.713 74.068 ;
			RECT	62.849 74.004 62.881 74.068 ;
			RECT	63.017 74.004 63.049 74.068 ;
			RECT	63.185 74.004 63.217 74.068 ;
			RECT	63.353 74.004 63.385 74.068 ;
			RECT	63.521 74.004 63.553 74.068 ;
			RECT	63.689 74.004 63.721 74.068 ;
			RECT	63.857 74.004 63.889 74.068 ;
			RECT	64.025 74.004 64.057 74.068 ;
			RECT	64.193 74.004 64.225 74.068 ;
			RECT	64.361 74.004 64.393 74.068 ;
			RECT	64.529 74.004 64.561 74.068 ;
			RECT	64.697 74.004 64.729 74.068 ;
			RECT	64.865 74.004 64.897 74.068 ;
			RECT	65.033 74.004 65.065 74.068 ;
			RECT	65.201 74.004 65.233 74.068 ;
			RECT	65.369 74.004 65.401 74.068 ;
			RECT	65.537 74.004 65.569 74.068 ;
			RECT	65.705 74.004 65.737 74.068 ;
			RECT	65.873 74.004 65.905 74.068 ;
			RECT	66.041 74.004 66.073 74.068 ;
			RECT	66.209 74.004 66.241 74.068 ;
			RECT	66.377 74.004 66.409 74.068 ;
			RECT	66.545 74.004 66.577 74.068 ;
			RECT	66.713 74.004 66.745 74.068 ;
			RECT	66.881 74.004 66.913 74.068 ;
			RECT	67.049 74.004 67.081 74.068 ;
			RECT	67.217 74.004 67.249 74.068 ;
			RECT	67.385 74.004 67.417 74.068 ;
			RECT	67.553 74.004 67.585 74.068 ;
			RECT	67.721 74.004 67.753 74.068 ;
			RECT	67.889 74.004 67.921 74.068 ;
			RECT	68.057 74.004 68.089 74.068 ;
			RECT	68.225 74.004 68.257 74.068 ;
			RECT	68.393 74.004 68.425 74.068 ;
			RECT	68.561 74.004 68.593 74.068 ;
			RECT	68.729 74.004 68.761 74.068 ;
			RECT	68.897 74.004 68.929 74.068 ;
			RECT	69.065 74.004 69.097 74.068 ;
			RECT	69.233 74.004 69.265 74.068 ;
			RECT	69.401 74.004 69.433 74.068 ;
			RECT	69.569 74.004 69.601 74.068 ;
			RECT	69.737 74.004 69.769 74.068 ;
			RECT	69.905 74.004 69.937 74.068 ;
			RECT	70.073 74.004 70.105 74.068 ;
			RECT	70.241 74.004 70.273 74.068 ;
			RECT	70.409 74.004 70.441 74.068 ;
			RECT	70.577 74.004 70.609 74.068 ;
			RECT	70.745 74.004 70.777 74.068 ;
			RECT	70.913 74.004 70.945 74.068 ;
			RECT	71.081 74.004 71.113 74.068 ;
			RECT	71.249 74.004 71.281 74.068 ;
			RECT	71.417 74.004 71.449 74.068 ;
			RECT	71.585 74.004 71.617 74.068 ;
			RECT	71.753 74.004 71.785 74.068 ;
			RECT	71.921 74.004 71.953 74.068 ;
			RECT	72.089 74.004 72.121 74.068 ;
			RECT	72.257 74.004 72.289 74.068 ;
			RECT	72.425 74.004 72.457 74.068 ;
			RECT	72.593 74.004 72.625 74.068 ;
			RECT	72.761 74.004 72.793 74.068 ;
			RECT	72.929 74.004 72.961 74.068 ;
			RECT	73.097 74.004 73.129 74.068 ;
			RECT	73.265 74.004 73.297 74.068 ;
			RECT	73.433 74.004 73.465 74.068 ;
			RECT	73.601 74.004 73.633 74.068 ;
			RECT	73.769 74.004 73.801 74.068 ;
			RECT	73.937 74.004 73.969 74.068 ;
			RECT	74.105 74.004 74.137 74.068 ;
			RECT	74.273 74.004 74.305 74.068 ;
			RECT	74.441 74.004 74.473 74.068 ;
			RECT	74.609 74.004 74.641 74.068 ;
			RECT	74.777 74.004 74.809 74.068 ;
			RECT	74.945 74.004 74.977 74.068 ;
			RECT	75.113 74.004 75.145 74.068 ;
			RECT	75.281 74.004 75.313 74.068 ;
			RECT	75.449 74.004 75.481 74.068 ;
			RECT	75.617 74.004 75.649 74.068 ;
			RECT	75.785 74.004 75.817 74.068 ;
			RECT	75.953 74.004 75.985 74.068 ;
			RECT	76.121 74.004 76.153 74.068 ;
			RECT	76.289 74.004 76.321 74.068 ;
			RECT	76.457 74.004 76.489 74.068 ;
			RECT	76.625 74.004 76.657 74.068 ;
			RECT	76.793 74.004 76.825 74.068 ;
			RECT	76.961 74.004 76.993 74.068 ;
			RECT	77.129 74.004 77.161 74.068 ;
			RECT	77.297 74.004 77.329 74.068 ;
			RECT	77.465 74.004 77.497 74.068 ;
			RECT	77.633 74.004 77.665 74.068 ;
			RECT	77.801 74.004 77.833 74.068 ;
			RECT	77.969 74.004 78.001 74.068 ;
			RECT	78.137 74.004 78.169 74.068 ;
			RECT	78.305 74.004 78.337 74.068 ;
			RECT	78.473 74.004 78.505 74.068 ;
			RECT	78.641 74.004 78.673 74.068 ;
			RECT	78.809 74.004 78.841 74.068 ;
			RECT	78.977 74.004 79.009 74.068 ;
			RECT	79.145 74.004 79.177 74.068 ;
			RECT	79.313 74.004 79.345 74.068 ;
			RECT	79.481 74.004 79.513 74.068 ;
			RECT	79.649 74.004 79.681 74.068 ;
			RECT	79.817 74.004 79.849 74.068 ;
			RECT	79.985 74.004 80.017 74.068 ;
			RECT	80.153 74.004 80.185 74.068 ;
			RECT	80.321 74.004 80.353 74.068 ;
			RECT	80.489 74.004 80.521 74.068 ;
			RECT	80.657 74.004 80.689 74.068 ;
			RECT	80.825 74.004 80.857 74.068 ;
			RECT	80.993 74.004 81.025 74.068 ;
			RECT	81.161 74.004 81.193 74.068 ;
			RECT	81.329 74.004 81.361 74.068 ;
			RECT	81.497 74.004 81.529 74.068 ;
			RECT	81.665 74.004 81.697 74.068 ;
			RECT	81.833 74.004 81.865 74.068 ;
			RECT	82.001 74.004 82.033 74.068 ;
			RECT	82.169 74.004 82.201 74.068 ;
			RECT	82.337 74.004 82.369 74.068 ;
			RECT	82.505 74.004 82.537 74.068 ;
			RECT	82.673 74.004 82.705 74.068 ;
			RECT	82.841 74.004 82.873 74.068 ;
			RECT	83.009 74.004 83.041 74.068 ;
			RECT	83.177 74.004 83.209 74.068 ;
			RECT	83.345 74.004 83.377 74.068 ;
			RECT	83.513 74.004 83.545 74.068 ;
			RECT	83.681 74.004 83.713 74.068 ;
			RECT	83.849 74.004 83.881 74.068 ;
			RECT	84.017 74.004 84.049 74.068 ;
			RECT	84.185 74.004 84.217 74.068 ;
			RECT	84.353 74.004 84.385 74.068 ;
			RECT	84.521 74.004 84.553 74.068 ;
			RECT	84.689 74.004 84.721 74.068 ;
			RECT	84.857 74.004 84.889 74.068 ;
			RECT	85.025 74.004 85.057 74.068 ;
			RECT	85.193 74.004 85.225 74.068 ;
			RECT	85.361 74.004 85.393 74.068 ;
			RECT	85.529 74.004 85.561 74.068 ;
			RECT	85.697 74.004 85.729 74.068 ;
			RECT	85.865 74.004 85.897 74.068 ;
			RECT	86.033 74.004 86.065 74.068 ;
			RECT	86.201 74.004 86.233 74.068 ;
			RECT	86.369 74.004 86.401 74.068 ;
			RECT	86.537 74.004 86.569 74.068 ;
			RECT	86.705 74.004 86.737 74.068 ;
			RECT	86.873 74.004 86.905 74.068 ;
			RECT	87.041 74.004 87.073 74.068 ;
			RECT	87.209 74.004 87.241 74.068 ;
			RECT	87.377 74.004 87.409 74.068 ;
			RECT	87.545 74.004 87.577 74.068 ;
			RECT	87.713 74.004 87.745 74.068 ;
			RECT	87.881 74.004 87.913 74.068 ;
			RECT	88.049 74.004 88.081 74.068 ;
			RECT	88.217 74.004 88.249 74.068 ;
			RECT	88.385 74.004 88.417 74.068 ;
			RECT	88.553 74.004 88.585 74.068 ;
			RECT	88.721 74.004 88.753 74.068 ;
			RECT	88.889 74.004 88.921 74.068 ;
			RECT	89.057 74.004 89.089 74.068 ;
			RECT	89.225 74.004 89.257 74.068 ;
			RECT	89.393 74.004 89.425 74.068 ;
			RECT	89.561 74.004 89.593 74.068 ;
			RECT	89.729 74.004 89.761 74.068 ;
			RECT	89.897 74.004 89.929 74.068 ;
			RECT	90.065 74.004 90.097 74.068 ;
			RECT	90.233 74.004 90.265 74.068 ;
			RECT	90.401 74.004 90.433 74.068 ;
			RECT	90.569 74.004 90.601 74.068 ;
			RECT	90.737 74.004 90.769 74.068 ;
			RECT	90.905 74.004 90.937 74.068 ;
			RECT	91.073 74.004 91.105 74.068 ;
			RECT	91.241 74.004 91.273 74.068 ;
			RECT	91.409 74.004 91.441 74.068 ;
			RECT	91.577 74.004 91.609 74.068 ;
			RECT	91.745 74.004 91.777 74.068 ;
			RECT	91.913 74.004 91.945 74.068 ;
			RECT	92.081 74.004 92.113 74.068 ;
			RECT	92.249 74.004 92.281 74.068 ;
			RECT	92.417 74.004 92.449 74.068 ;
			RECT	92.585 74.004 92.617 74.068 ;
			RECT	92.753 74.004 92.785 74.068 ;
			RECT	92.921 74.004 92.953 74.068 ;
			RECT	93.089 74.004 93.121 74.068 ;
			RECT	93.257 74.004 93.289 74.068 ;
			RECT	93.425 74.004 93.457 74.068 ;
			RECT	93.593 74.004 93.625 74.068 ;
			RECT	93.761 74.004 93.793 74.068 ;
			RECT	93.929 74.004 93.961 74.068 ;
			RECT	94.097 74.004 94.129 74.068 ;
			RECT	94.265 74.004 94.297 74.068 ;
			RECT	94.433 74.004 94.465 74.068 ;
			RECT	94.601 74.004 94.633 74.068 ;
			RECT	94.769 74.004 94.801 74.068 ;
			RECT	94.937 74.004 94.969 74.068 ;
			RECT	95.105 74.004 95.137 74.068 ;
			RECT	95.273 74.004 95.305 74.068 ;
			RECT	95.441 74.004 95.473 74.068 ;
			RECT	95.609 74.004 95.641 74.068 ;
			RECT	95.777 74.004 95.809 74.068 ;
			RECT	95.945 74.004 95.977 74.068 ;
			RECT	96.113 74.004 96.145 74.068 ;
			RECT	96.281 74.004 96.313 74.068 ;
			RECT	96.449 74.004 96.481 74.068 ;
			RECT	96.617 74.004 96.649 74.068 ;
			RECT	96.785 74.004 96.817 74.068 ;
			RECT	96.953 74.004 96.985 74.068 ;
			RECT	97.121 74.004 97.153 74.068 ;
			RECT	97.289 74.004 97.321 74.068 ;
			RECT	97.457 74.004 97.489 74.068 ;
			RECT	97.625 74.004 97.657 74.068 ;
			RECT	97.793 74.004 97.825 74.068 ;
			RECT	97.961 74.004 97.993 74.068 ;
			RECT	98.129 74.004 98.161 74.068 ;
			RECT	98.297 74.004 98.329 74.068 ;
			RECT	98.465 74.004 98.497 74.068 ;
			RECT	98.633 74.004 98.665 74.068 ;
			RECT	98.801 74.004 98.833 74.068 ;
			RECT	98.969 74.004 99.001 74.068 ;
			RECT	99.137 74.004 99.169 74.068 ;
			RECT	99.305 74.004 99.337 74.068 ;
			RECT	99.473 74.004 99.505 74.068 ;
			RECT	99.641 74.004 99.673 74.068 ;
			RECT	99.809 74.004 99.841 74.068 ;
			RECT	99.977 74.004 100.009 74.068 ;
			RECT	100.145 74.004 100.177 74.068 ;
			RECT	100.313 74.004 100.345 74.068 ;
			RECT	100.481 74.004 100.513 74.068 ;
			RECT	100.649 74.004 100.681 74.068 ;
			RECT	100.817 74.004 100.849 74.068 ;
			RECT	100.985 74.004 101.017 74.068 ;
			RECT	101.153 74.004 101.185 74.068 ;
			RECT	101.321 74.004 101.353 74.068 ;
			RECT	101.489 74.004 101.521 74.068 ;
			RECT	101.657 74.004 101.689 74.068 ;
			RECT	101.825 74.004 101.857 74.068 ;
			RECT	101.993 74.004 102.025 74.068 ;
			RECT	102.123 74.02 102.155 74.052 ;
			RECT	102.245 74.015 102.277 74.047 ;
			RECT	102.375 74.004 102.407 74.068 ;
			RECT	103.795 74.004 103.827 74.068 ;
			RECT	103.925 74.015 103.957 74.047 ;
			RECT	104.047 74.02 104.079 74.052 ;
			RECT	104.177 74.004 104.209 74.068 ;
			RECT	104.345 74.004 104.377 74.068 ;
			RECT	104.513 74.004 104.545 74.068 ;
			RECT	104.681 74.004 104.713 74.068 ;
			RECT	104.849 74.004 104.881 74.068 ;
			RECT	105.017 74.004 105.049 74.068 ;
			RECT	105.185 74.004 105.217 74.068 ;
			RECT	105.353 74.004 105.385 74.068 ;
			RECT	105.521 74.004 105.553 74.068 ;
			RECT	105.689 74.004 105.721 74.068 ;
			RECT	105.857 74.004 105.889 74.068 ;
			RECT	106.025 74.004 106.057 74.068 ;
			RECT	106.193 74.004 106.225 74.068 ;
			RECT	106.361 74.004 106.393 74.068 ;
			RECT	106.529 74.004 106.561 74.068 ;
			RECT	106.697 74.004 106.729 74.068 ;
			RECT	106.865 74.004 106.897 74.068 ;
			RECT	107.033 74.004 107.065 74.068 ;
			RECT	107.201 74.004 107.233 74.068 ;
			RECT	107.369 74.004 107.401 74.068 ;
			RECT	107.537 74.004 107.569 74.068 ;
			RECT	107.705 74.004 107.737 74.068 ;
			RECT	107.873 74.004 107.905 74.068 ;
			RECT	108.041 74.004 108.073 74.068 ;
			RECT	108.209 74.004 108.241 74.068 ;
			RECT	108.377 74.004 108.409 74.068 ;
			RECT	108.545 74.004 108.577 74.068 ;
			RECT	108.713 74.004 108.745 74.068 ;
			RECT	108.881 74.004 108.913 74.068 ;
			RECT	109.049 74.004 109.081 74.068 ;
			RECT	109.217 74.004 109.249 74.068 ;
			RECT	109.385 74.004 109.417 74.068 ;
			RECT	109.553 74.004 109.585 74.068 ;
			RECT	109.721 74.004 109.753 74.068 ;
			RECT	109.889 74.004 109.921 74.068 ;
			RECT	110.057 74.004 110.089 74.068 ;
			RECT	110.225 74.004 110.257 74.068 ;
			RECT	110.393 74.004 110.425 74.068 ;
			RECT	110.561 74.004 110.593 74.068 ;
			RECT	110.729 74.004 110.761 74.068 ;
			RECT	110.897 74.004 110.929 74.068 ;
			RECT	111.065 74.004 111.097 74.068 ;
			RECT	111.233 74.004 111.265 74.068 ;
			RECT	111.401 74.004 111.433 74.068 ;
			RECT	111.569 74.004 111.601 74.068 ;
			RECT	111.737 74.004 111.769 74.068 ;
			RECT	111.905 74.004 111.937 74.068 ;
			RECT	112.073 74.004 112.105 74.068 ;
			RECT	112.241 74.004 112.273 74.068 ;
			RECT	112.409 74.004 112.441 74.068 ;
			RECT	112.577 74.004 112.609 74.068 ;
			RECT	112.745 74.004 112.777 74.068 ;
			RECT	112.913 74.004 112.945 74.068 ;
			RECT	113.081 74.004 113.113 74.068 ;
			RECT	113.249 74.004 113.281 74.068 ;
			RECT	113.417 74.004 113.449 74.068 ;
			RECT	113.585 74.004 113.617 74.068 ;
			RECT	113.753 74.004 113.785 74.068 ;
			RECT	113.921 74.004 113.953 74.068 ;
			RECT	114.089 74.004 114.121 74.068 ;
			RECT	114.257 74.004 114.289 74.068 ;
			RECT	114.425 74.004 114.457 74.068 ;
			RECT	114.593 74.004 114.625 74.068 ;
			RECT	114.761 74.004 114.793 74.068 ;
			RECT	114.929 74.004 114.961 74.068 ;
			RECT	115.097 74.004 115.129 74.068 ;
			RECT	115.265 74.004 115.297 74.068 ;
			RECT	115.433 74.004 115.465 74.068 ;
			RECT	115.601 74.004 115.633 74.068 ;
			RECT	115.769 74.004 115.801 74.068 ;
			RECT	115.937 74.004 115.969 74.068 ;
			RECT	116.105 74.004 116.137 74.068 ;
			RECT	116.273 74.004 116.305 74.068 ;
			RECT	116.441 74.004 116.473 74.068 ;
			RECT	116.609 74.004 116.641 74.068 ;
			RECT	116.777 74.004 116.809 74.068 ;
			RECT	116.945 74.004 116.977 74.068 ;
			RECT	117.113 74.004 117.145 74.068 ;
			RECT	117.281 74.004 117.313 74.068 ;
			RECT	117.449 74.004 117.481 74.068 ;
			RECT	117.617 74.004 117.649 74.068 ;
			RECT	117.785 74.004 117.817 74.068 ;
			RECT	117.953 74.004 117.985 74.068 ;
			RECT	118.121 74.004 118.153 74.068 ;
			RECT	118.289 74.004 118.321 74.068 ;
			RECT	118.457 74.004 118.489 74.068 ;
			RECT	118.625 74.004 118.657 74.068 ;
			RECT	118.793 74.004 118.825 74.068 ;
			RECT	118.961 74.004 118.993 74.068 ;
			RECT	119.129 74.004 119.161 74.068 ;
			RECT	119.297 74.004 119.329 74.068 ;
			RECT	119.465 74.004 119.497 74.068 ;
			RECT	119.633 74.004 119.665 74.068 ;
			RECT	119.801 74.004 119.833 74.068 ;
			RECT	119.969 74.004 120.001 74.068 ;
			RECT	120.137 74.004 120.169 74.068 ;
			RECT	120.305 74.004 120.337 74.068 ;
			RECT	120.473 74.004 120.505 74.068 ;
			RECT	120.641 74.004 120.673 74.068 ;
			RECT	120.809 74.004 120.841 74.068 ;
			RECT	120.977 74.004 121.009 74.068 ;
			RECT	121.145 74.004 121.177 74.068 ;
			RECT	121.313 74.004 121.345 74.068 ;
			RECT	121.481 74.004 121.513 74.068 ;
			RECT	121.649 74.004 121.681 74.068 ;
			RECT	121.817 74.004 121.849 74.068 ;
			RECT	121.985 74.004 122.017 74.068 ;
			RECT	122.153 74.004 122.185 74.068 ;
			RECT	122.321 74.004 122.353 74.068 ;
			RECT	122.489 74.004 122.521 74.068 ;
			RECT	122.657 74.004 122.689 74.068 ;
			RECT	122.825 74.004 122.857 74.068 ;
			RECT	122.993 74.004 123.025 74.068 ;
			RECT	123.161 74.004 123.193 74.068 ;
			RECT	123.329 74.004 123.361 74.068 ;
			RECT	123.497 74.004 123.529 74.068 ;
			RECT	123.665 74.004 123.697 74.068 ;
			RECT	123.833 74.004 123.865 74.068 ;
			RECT	124.001 74.004 124.033 74.068 ;
			RECT	124.169 74.004 124.201 74.068 ;
			RECT	124.337 74.004 124.369 74.068 ;
			RECT	124.505 74.004 124.537 74.068 ;
			RECT	124.673 74.004 124.705 74.068 ;
			RECT	124.841 74.004 124.873 74.068 ;
			RECT	125.009 74.004 125.041 74.068 ;
			RECT	125.177 74.004 125.209 74.068 ;
			RECT	125.345 74.004 125.377 74.068 ;
			RECT	125.513 74.004 125.545 74.068 ;
			RECT	125.681 74.004 125.713 74.068 ;
			RECT	125.849 74.004 125.881 74.068 ;
			RECT	126.017 74.004 126.049 74.068 ;
			RECT	126.185 74.004 126.217 74.068 ;
			RECT	126.353 74.004 126.385 74.068 ;
			RECT	126.521 74.004 126.553 74.068 ;
			RECT	126.689 74.004 126.721 74.068 ;
			RECT	126.857 74.004 126.889 74.068 ;
			RECT	127.025 74.004 127.057 74.068 ;
			RECT	127.193 74.004 127.225 74.068 ;
			RECT	127.361 74.004 127.393 74.068 ;
			RECT	127.529 74.004 127.561 74.068 ;
			RECT	127.697 74.004 127.729 74.068 ;
			RECT	127.865 74.004 127.897 74.068 ;
			RECT	128.033 74.004 128.065 74.068 ;
			RECT	128.201 74.004 128.233 74.068 ;
			RECT	128.369 74.004 128.401 74.068 ;
			RECT	128.537 74.004 128.569 74.068 ;
			RECT	128.705 74.004 128.737 74.068 ;
			RECT	128.873 74.004 128.905 74.068 ;
			RECT	129.041 74.004 129.073 74.068 ;
			RECT	129.209 74.004 129.241 74.068 ;
			RECT	129.377 74.004 129.409 74.068 ;
			RECT	129.545 74.004 129.577 74.068 ;
			RECT	129.713 74.004 129.745 74.068 ;
			RECT	129.881 74.004 129.913 74.068 ;
			RECT	130.049 74.004 130.081 74.068 ;
			RECT	130.217 74.004 130.249 74.068 ;
			RECT	130.385 74.004 130.417 74.068 ;
			RECT	130.553 74.004 130.585 74.068 ;
			RECT	130.721 74.004 130.753 74.068 ;
			RECT	130.889 74.004 130.921 74.068 ;
			RECT	131.057 74.004 131.089 74.068 ;
			RECT	131.225 74.004 131.257 74.068 ;
			RECT	131.393 74.004 131.425 74.068 ;
			RECT	131.561 74.004 131.593 74.068 ;
			RECT	131.729 74.004 131.761 74.068 ;
			RECT	131.897 74.004 131.929 74.068 ;
			RECT	132.065 74.004 132.097 74.068 ;
			RECT	132.233 74.004 132.265 74.068 ;
			RECT	132.401 74.004 132.433 74.068 ;
			RECT	132.569 74.004 132.601 74.068 ;
			RECT	132.737 74.004 132.769 74.068 ;
			RECT	132.905 74.004 132.937 74.068 ;
			RECT	133.073 74.004 133.105 74.068 ;
			RECT	133.241 74.004 133.273 74.068 ;
			RECT	133.409 74.004 133.441 74.068 ;
			RECT	133.577 74.004 133.609 74.068 ;
			RECT	133.745 74.004 133.777 74.068 ;
			RECT	133.913 74.004 133.945 74.068 ;
			RECT	134.081 74.004 134.113 74.068 ;
			RECT	134.249 74.004 134.281 74.068 ;
			RECT	134.417 74.004 134.449 74.068 ;
			RECT	134.585 74.004 134.617 74.068 ;
			RECT	134.753 74.004 134.785 74.068 ;
			RECT	134.921 74.004 134.953 74.068 ;
			RECT	135.089 74.004 135.121 74.068 ;
			RECT	135.257 74.004 135.289 74.068 ;
			RECT	135.425 74.004 135.457 74.068 ;
			RECT	135.593 74.004 135.625 74.068 ;
			RECT	135.761 74.004 135.793 74.068 ;
			RECT	135.929 74.004 135.961 74.068 ;
			RECT	136.097 74.004 136.129 74.068 ;
			RECT	136.265 74.004 136.297 74.068 ;
			RECT	136.433 74.004 136.465 74.068 ;
			RECT	136.601 74.004 136.633 74.068 ;
			RECT	136.769 74.004 136.801 74.068 ;
			RECT	136.937 74.004 136.969 74.068 ;
			RECT	137.105 74.004 137.137 74.068 ;
			RECT	137.273 74.004 137.305 74.068 ;
			RECT	137.441 74.004 137.473 74.068 ;
			RECT	137.609 74.004 137.641 74.068 ;
			RECT	137.777 74.004 137.809 74.068 ;
			RECT	137.945 74.004 137.977 74.068 ;
			RECT	138.113 74.004 138.145 74.068 ;
			RECT	138.281 74.004 138.313 74.068 ;
			RECT	138.449 74.004 138.481 74.068 ;
			RECT	138.617 74.004 138.649 74.068 ;
			RECT	138.785 74.004 138.817 74.068 ;
			RECT	138.953 74.004 138.985 74.068 ;
			RECT	139.121 74.004 139.153 74.068 ;
			RECT	139.289 74.004 139.321 74.068 ;
			RECT	139.457 74.004 139.489 74.068 ;
			RECT	139.625 74.004 139.657 74.068 ;
			RECT	139.793 74.004 139.825 74.068 ;
			RECT	139.961 74.004 139.993 74.068 ;
			RECT	140.129 74.004 140.161 74.068 ;
			RECT	140.297 74.004 140.329 74.068 ;
			RECT	140.465 74.004 140.497 74.068 ;
			RECT	140.633 74.004 140.665 74.068 ;
			RECT	140.801 74.004 140.833 74.068 ;
			RECT	140.969 74.004 141.001 74.068 ;
			RECT	141.137 74.004 141.169 74.068 ;
			RECT	141.305 74.004 141.337 74.068 ;
			RECT	141.473 74.004 141.505 74.068 ;
			RECT	141.641 74.004 141.673 74.068 ;
			RECT	141.809 74.004 141.841 74.068 ;
			RECT	141.977 74.004 142.009 74.068 ;
			RECT	142.145 74.004 142.177 74.068 ;
			RECT	142.313 74.004 142.345 74.068 ;
			RECT	142.481 74.004 142.513 74.068 ;
			RECT	142.649 74.004 142.681 74.068 ;
			RECT	142.817 74.004 142.849 74.068 ;
			RECT	142.985 74.004 143.017 74.068 ;
			RECT	143.153 74.004 143.185 74.068 ;
			RECT	143.321 74.004 143.353 74.068 ;
			RECT	143.489 74.004 143.521 74.068 ;
			RECT	143.657 74.004 143.689 74.068 ;
			RECT	143.825 74.004 143.857 74.068 ;
			RECT	143.993 74.004 144.025 74.068 ;
			RECT	144.161 74.004 144.193 74.068 ;
			RECT	144.329 74.004 144.361 74.068 ;
			RECT	144.497 74.004 144.529 74.068 ;
			RECT	144.665 74.004 144.697 74.068 ;
			RECT	144.833 74.004 144.865 74.068 ;
			RECT	145.001 74.004 145.033 74.068 ;
			RECT	145.169 74.004 145.201 74.068 ;
			RECT	145.337 74.004 145.369 74.068 ;
			RECT	145.505 74.004 145.537 74.068 ;
			RECT	145.673 74.004 145.705 74.068 ;
			RECT	145.841 74.004 145.873 74.068 ;
			RECT	146.009 74.004 146.041 74.068 ;
			RECT	146.177 74.004 146.209 74.068 ;
			RECT	146.345 74.004 146.377 74.068 ;
			RECT	146.513 74.004 146.545 74.068 ;
			RECT	146.681 74.004 146.713 74.068 ;
			RECT	146.849 74.004 146.881 74.068 ;
			RECT	147.017 74.004 147.049 74.068 ;
			RECT	147.185 74.004 147.217 74.068 ;
			RECT	147.316 74.02 147.348 74.052 ;
			RECT	147.437 74.02 147.469 74.052 ;
			RECT	147.567 74.004 147.599 74.068 ;
			RECT	149.879 74.004 149.911 74.068 ;
			RECT	151.13 74.004 151.194 74.068 ;
			RECT	151.81 74.004 151.842 74.068 ;
			RECT	152.249 74.004 152.281 74.068 ;
			RECT	153.56 74.004 153.624 74.068 ;
			RECT	156.601 74.004 156.633 74.068 ;
			RECT	156.731 74.02 156.763 74.052 ;
			RECT	156.852 74.02 156.884 74.052 ;
			RECT	156.983 74.004 157.015 74.068 ;
			RECT	157.151 74.004 157.183 74.068 ;
			RECT	157.319 74.004 157.351 74.068 ;
			RECT	157.487 74.004 157.519 74.068 ;
			RECT	157.655 74.004 157.687 74.068 ;
			RECT	157.823 74.004 157.855 74.068 ;
			RECT	157.991 74.004 158.023 74.068 ;
			RECT	158.159 74.004 158.191 74.068 ;
			RECT	158.327 74.004 158.359 74.068 ;
			RECT	158.495 74.004 158.527 74.068 ;
			RECT	158.663 74.004 158.695 74.068 ;
			RECT	158.831 74.004 158.863 74.068 ;
			RECT	158.999 74.004 159.031 74.068 ;
			RECT	159.167 74.004 159.199 74.068 ;
			RECT	159.335 74.004 159.367 74.068 ;
			RECT	159.503 74.004 159.535 74.068 ;
			RECT	159.671 74.004 159.703 74.068 ;
			RECT	159.839 74.004 159.871 74.068 ;
			RECT	160.007 74.004 160.039 74.068 ;
			RECT	160.175 74.004 160.207 74.068 ;
			RECT	160.343 74.004 160.375 74.068 ;
			RECT	160.511 74.004 160.543 74.068 ;
			RECT	160.679 74.004 160.711 74.068 ;
			RECT	160.847 74.004 160.879 74.068 ;
			RECT	161.015 74.004 161.047 74.068 ;
			RECT	161.183 74.004 161.215 74.068 ;
			RECT	161.351 74.004 161.383 74.068 ;
			RECT	161.519 74.004 161.551 74.068 ;
			RECT	161.687 74.004 161.719 74.068 ;
			RECT	161.855 74.004 161.887 74.068 ;
			RECT	162.023 74.004 162.055 74.068 ;
			RECT	162.191 74.004 162.223 74.068 ;
			RECT	162.359 74.004 162.391 74.068 ;
			RECT	162.527 74.004 162.559 74.068 ;
			RECT	162.695 74.004 162.727 74.068 ;
			RECT	162.863 74.004 162.895 74.068 ;
			RECT	163.031 74.004 163.063 74.068 ;
			RECT	163.199 74.004 163.231 74.068 ;
			RECT	163.367 74.004 163.399 74.068 ;
			RECT	163.535 74.004 163.567 74.068 ;
			RECT	163.703 74.004 163.735 74.068 ;
			RECT	163.871 74.004 163.903 74.068 ;
			RECT	164.039 74.004 164.071 74.068 ;
			RECT	164.207 74.004 164.239 74.068 ;
			RECT	164.375 74.004 164.407 74.068 ;
			RECT	164.543 74.004 164.575 74.068 ;
			RECT	164.711 74.004 164.743 74.068 ;
			RECT	164.879 74.004 164.911 74.068 ;
			RECT	165.047 74.004 165.079 74.068 ;
			RECT	165.215 74.004 165.247 74.068 ;
			RECT	165.383 74.004 165.415 74.068 ;
			RECT	165.551 74.004 165.583 74.068 ;
			RECT	165.719 74.004 165.751 74.068 ;
			RECT	165.887 74.004 165.919 74.068 ;
			RECT	166.055 74.004 166.087 74.068 ;
			RECT	166.223 74.004 166.255 74.068 ;
			RECT	166.391 74.004 166.423 74.068 ;
			RECT	166.559 74.004 166.591 74.068 ;
			RECT	166.727 74.004 166.759 74.068 ;
			RECT	166.895 74.004 166.927 74.068 ;
			RECT	167.063 74.004 167.095 74.068 ;
			RECT	167.231 74.004 167.263 74.068 ;
			RECT	167.399 74.004 167.431 74.068 ;
			RECT	167.567 74.004 167.599 74.068 ;
			RECT	167.735 74.004 167.767 74.068 ;
			RECT	167.903 74.004 167.935 74.068 ;
			RECT	168.071 74.004 168.103 74.068 ;
			RECT	168.239 74.004 168.271 74.068 ;
			RECT	168.407 74.004 168.439 74.068 ;
			RECT	168.575 74.004 168.607 74.068 ;
			RECT	168.743 74.004 168.775 74.068 ;
			RECT	168.911 74.004 168.943 74.068 ;
			RECT	169.079 74.004 169.111 74.068 ;
			RECT	169.247 74.004 169.279 74.068 ;
			RECT	169.415 74.004 169.447 74.068 ;
			RECT	169.583 74.004 169.615 74.068 ;
			RECT	169.751 74.004 169.783 74.068 ;
			RECT	169.919 74.004 169.951 74.068 ;
			RECT	170.087 74.004 170.119 74.068 ;
			RECT	170.255 74.004 170.287 74.068 ;
			RECT	170.423 74.004 170.455 74.068 ;
			RECT	170.591 74.004 170.623 74.068 ;
			RECT	170.759 74.004 170.791 74.068 ;
			RECT	170.927 74.004 170.959 74.068 ;
			RECT	171.095 74.004 171.127 74.068 ;
			RECT	171.263 74.004 171.295 74.068 ;
			RECT	171.431 74.004 171.463 74.068 ;
			RECT	171.599 74.004 171.631 74.068 ;
			RECT	171.767 74.004 171.799 74.068 ;
			RECT	171.935 74.004 171.967 74.068 ;
			RECT	172.103 74.004 172.135 74.068 ;
			RECT	172.271 74.004 172.303 74.068 ;
			RECT	172.439 74.004 172.471 74.068 ;
			RECT	172.607 74.004 172.639 74.068 ;
			RECT	172.775 74.004 172.807 74.068 ;
			RECT	172.943 74.004 172.975 74.068 ;
			RECT	173.111 74.004 173.143 74.068 ;
			RECT	173.279 74.004 173.311 74.068 ;
			RECT	173.447 74.004 173.479 74.068 ;
			RECT	173.615 74.004 173.647 74.068 ;
			RECT	173.783 74.004 173.815 74.068 ;
			RECT	173.951 74.004 173.983 74.068 ;
			RECT	174.119 74.004 174.151 74.068 ;
			RECT	174.287 74.004 174.319 74.068 ;
			RECT	174.455 74.004 174.487 74.068 ;
			RECT	174.623 74.004 174.655 74.068 ;
			RECT	174.791 74.004 174.823 74.068 ;
			RECT	174.959 74.004 174.991 74.068 ;
			RECT	175.127 74.004 175.159 74.068 ;
			RECT	175.295 74.004 175.327 74.068 ;
			RECT	175.463 74.004 175.495 74.068 ;
			RECT	175.631 74.004 175.663 74.068 ;
			RECT	175.799 74.004 175.831 74.068 ;
			RECT	175.967 74.004 175.999 74.068 ;
			RECT	176.135 74.004 176.167 74.068 ;
			RECT	176.303 74.004 176.335 74.068 ;
			RECT	176.471 74.004 176.503 74.068 ;
			RECT	176.639 74.004 176.671 74.068 ;
			RECT	176.807 74.004 176.839 74.068 ;
			RECT	176.975 74.004 177.007 74.068 ;
			RECT	177.143 74.004 177.175 74.068 ;
			RECT	177.311 74.004 177.343 74.068 ;
			RECT	177.479 74.004 177.511 74.068 ;
			RECT	177.647 74.004 177.679 74.068 ;
			RECT	177.815 74.004 177.847 74.068 ;
			RECT	177.983 74.004 178.015 74.068 ;
			RECT	178.151 74.004 178.183 74.068 ;
			RECT	178.319 74.004 178.351 74.068 ;
			RECT	178.487 74.004 178.519 74.068 ;
			RECT	178.655 74.004 178.687 74.068 ;
			RECT	178.823 74.004 178.855 74.068 ;
			RECT	178.991 74.004 179.023 74.068 ;
			RECT	179.159 74.004 179.191 74.068 ;
			RECT	179.327 74.004 179.359 74.068 ;
			RECT	179.495 74.004 179.527 74.068 ;
			RECT	179.663 74.004 179.695 74.068 ;
			RECT	179.831 74.004 179.863 74.068 ;
			RECT	179.999 74.004 180.031 74.068 ;
			RECT	180.167 74.004 180.199 74.068 ;
			RECT	180.335 74.004 180.367 74.068 ;
			RECT	180.503 74.004 180.535 74.068 ;
			RECT	180.671 74.004 180.703 74.068 ;
			RECT	180.839 74.004 180.871 74.068 ;
			RECT	181.007 74.004 181.039 74.068 ;
			RECT	181.175 74.004 181.207 74.068 ;
			RECT	181.343 74.004 181.375 74.068 ;
			RECT	181.511 74.004 181.543 74.068 ;
			RECT	181.679 74.004 181.711 74.068 ;
			RECT	181.847 74.004 181.879 74.068 ;
			RECT	182.015 74.004 182.047 74.068 ;
			RECT	182.183 74.004 182.215 74.068 ;
			RECT	182.351 74.004 182.383 74.068 ;
			RECT	182.519 74.004 182.551 74.068 ;
			RECT	182.687 74.004 182.719 74.068 ;
			RECT	182.855 74.004 182.887 74.068 ;
			RECT	183.023 74.004 183.055 74.068 ;
			RECT	183.191 74.004 183.223 74.068 ;
			RECT	183.359 74.004 183.391 74.068 ;
			RECT	183.527 74.004 183.559 74.068 ;
			RECT	183.695 74.004 183.727 74.068 ;
			RECT	183.863 74.004 183.895 74.068 ;
			RECT	184.031 74.004 184.063 74.068 ;
			RECT	184.199 74.004 184.231 74.068 ;
			RECT	184.367 74.004 184.399 74.068 ;
			RECT	184.535 74.004 184.567 74.068 ;
			RECT	184.703 74.004 184.735 74.068 ;
			RECT	184.871 74.004 184.903 74.068 ;
			RECT	185.039 74.004 185.071 74.068 ;
			RECT	185.207 74.004 185.239 74.068 ;
			RECT	185.375 74.004 185.407 74.068 ;
			RECT	185.543 74.004 185.575 74.068 ;
			RECT	185.711 74.004 185.743 74.068 ;
			RECT	185.879 74.004 185.911 74.068 ;
			RECT	186.047 74.004 186.079 74.068 ;
			RECT	186.215 74.004 186.247 74.068 ;
			RECT	186.383 74.004 186.415 74.068 ;
			RECT	186.551 74.004 186.583 74.068 ;
			RECT	186.719 74.004 186.751 74.068 ;
			RECT	186.887 74.004 186.919 74.068 ;
			RECT	187.055 74.004 187.087 74.068 ;
			RECT	187.223 74.004 187.255 74.068 ;
			RECT	187.391 74.004 187.423 74.068 ;
			RECT	187.559 74.004 187.591 74.068 ;
			RECT	187.727 74.004 187.759 74.068 ;
			RECT	187.895 74.004 187.927 74.068 ;
			RECT	188.063 74.004 188.095 74.068 ;
			RECT	188.231 74.004 188.263 74.068 ;
			RECT	188.399 74.004 188.431 74.068 ;
			RECT	188.567 74.004 188.599 74.068 ;
			RECT	188.735 74.004 188.767 74.068 ;
			RECT	188.903 74.004 188.935 74.068 ;
			RECT	189.071 74.004 189.103 74.068 ;
			RECT	189.239 74.004 189.271 74.068 ;
			RECT	189.407 74.004 189.439 74.068 ;
			RECT	189.575 74.004 189.607 74.068 ;
			RECT	189.743 74.004 189.775 74.068 ;
			RECT	189.911 74.004 189.943 74.068 ;
			RECT	190.079 74.004 190.111 74.068 ;
			RECT	190.247 74.004 190.279 74.068 ;
			RECT	190.415 74.004 190.447 74.068 ;
			RECT	190.583 74.004 190.615 74.068 ;
			RECT	190.751 74.004 190.783 74.068 ;
			RECT	190.919 74.004 190.951 74.068 ;
			RECT	191.087 74.004 191.119 74.068 ;
			RECT	191.255 74.004 191.287 74.068 ;
			RECT	191.423 74.004 191.455 74.068 ;
			RECT	191.591 74.004 191.623 74.068 ;
			RECT	191.759 74.004 191.791 74.068 ;
			RECT	191.927 74.004 191.959 74.068 ;
			RECT	192.095 74.004 192.127 74.068 ;
			RECT	192.263 74.004 192.295 74.068 ;
			RECT	192.431 74.004 192.463 74.068 ;
			RECT	192.599 74.004 192.631 74.068 ;
			RECT	192.767 74.004 192.799 74.068 ;
			RECT	192.935 74.004 192.967 74.068 ;
			RECT	193.103 74.004 193.135 74.068 ;
			RECT	193.271 74.004 193.303 74.068 ;
			RECT	193.439 74.004 193.471 74.068 ;
			RECT	193.607 74.004 193.639 74.068 ;
			RECT	193.775 74.004 193.807 74.068 ;
			RECT	193.943 74.004 193.975 74.068 ;
			RECT	194.111 74.004 194.143 74.068 ;
			RECT	194.279 74.004 194.311 74.068 ;
			RECT	194.447 74.004 194.479 74.068 ;
			RECT	194.615 74.004 194.647 74.068 ;
			RECT	194.783 74.004 194.815 74.068 ;
			RECT	194.951 74.004 194.983 74.068 ;
			RECT	195.119 74.004 195.151 74.068 ;
			RECT	195.287 74.004 195.319 74.068 ;
			RECT	195.455 74.004 195.487 74.068 ;
			RECT	195.623 74.004 195.655 74.068 ;
			RECT	195.791 74.004 195.823 74.068 ;
			RECT	195.959 74.004 195.991 74.068 ;
			RECT	196.127 74.004 196.159 74.068 ;
			RECT	196.295 74.004 196.327 74.068 ;
			RECT	196.463 74.004 196.495 74.068 ;
			RECT	196.631 74.004 196.663 74.068 ;
			RECT	196.799 74.004 196.831 74.068 ;
			RECT	196.967 74.004 196.999 74.068 ;
			RECT	197.135 74.004 197.167 74.068 ;
			RECT	197.303 74.004 197.335 74.068 ;
			RECT	197.471 74.004 197.503 74.068 ;
			RECT	197.639 74.004 197.671 74.068 ;
			RECT	197.807 74.004 197.839 74.068 ;
			RECT	197.975 74.004 198.007 74.068 ;
			RECT	198.143 74.004 198.175 74.068 ;
			RECT	198.311 74.004 198.343 74.068 ;
			RECT	198.479 74.004 198.511 74.068 ;
			RECT	198.647 74.004 198.679 74.068 ;
			RECT	198.815 74.004 198.847 74.068 ;
			RECT	198.983 74.004 199.015 74.068 ;
			RECT	199.151 74.004 199.183 74.068 ;
			RECT	199.319 74.004 199.351 74.068 ;
			RECT	199.487 74.004 199.519 74.068 ;
			RECT	199.655 74.004 199.687 74.068 ;
			RECT	199.823 74.004 199.855 74.068 ;
			RECT	199.991 74.004 200.023 74.068 ;
			RECT	200.121 74.02 200.153 74.052 ;
			RECT	200.243 74.015 200.275 74.047 ;
			RECT	200.373 74.004 200.405 74.068 ;
			RECT	200.9 74.004 200.932 74.068 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 8.08 201.665 8.2 ;
			LAYER	J3 ;
			RECT	0.755 8.108 0.787 8.172 ;
			RECT	1.645 8.108 1.709 8.172 ;
			RECT	2.323 8.108 2.387 8.172 ;
			RECT	3.438 8.108 3.47 8.172 ;
			RECT	3.585 8.108 3.617 8.172 ;
			RECT	4.195 8.108 4.227 8.172 ;
			RECT	4.72 8.108 4.752 8.172 ;
			RECT	4.944 8.108 5.008 8.172 ;
			RECT	5.267 8.108 5.299 8.172 ;
			RECT	5.797 8.108 5.829 8.172 ;
			RECT	5.927 8.129 5.959 8.161 ;
			RECT	6.049 8.124 6.081 8.156 ;
			RECT	6.179 8.108 6.211 8.172 ;
			RECT	6.347 8.108 6.379 8.172 ;
			RECT	6.515 8.108 6.547 8.172 ;
			RECT	6.683 8.108 6.715 8.172 ;
			RECT	6.851 8.108 6.883 8.172 ;
			RECT	7.019 8.108 7.051 8.172 ;
			RECT	7.187 8.108 7.219 8.172 ;
			RECT	7.355 8.108 7.387 8.172 ;
			RECT	7.523 8.108 7.555 8.172 ;
			RECT	7.691 8.108 7.723 8.172 ;
			RECT	7.859 8.108 7.891 8.172 ;
			RECT	8.027 8.108 8.059 8.172 ;
			RECT	8.195 8.108 8.227 8.172 ;
			RECT	8.363 8.108 8.395 8.172 ;
			RECT	8.531 8.108 8.563 8.172 ;
			RECT	8.699 8.108 8.731 8.172 ;
			RECT	8.867 8.108 8.899 8.172 ;
			RECT	9.035 8.108 9.067 8.172 ;
			RECT	9.203 8.108 9.235 8.172 ;
			RECT	9.371 8.108 9.403 8.172 ;
			RECT	9.539 8.108 9.571 8.172 ;
			RECT	9.707 8.108 9.739 8.172 ;
			RECT	9.875 8.108 9.907 8.172 ;
			RECT	10.043 8.108 10.075 8.172 ;
			RECT	10.211 8.108 10.243 8.172 ;
			RECT	10.379 8.108 10.411 8.172 ;
			RECT	10.547 8.108 10.579 8.172 ;
			RECT	10.715 8.108 10.747 8.172 ;
			RECT	10.883 8.108 10.915 8.172 ;
			RECT	11.051 8.108 11.083 8.172 ;
			RECT	11.219 8.108 11.251 8.172 ;
			RECT	11.387 8.108 11.419 8.172 ;
			RECT	11.555 8.108 11.587 8.172 ;
			RECT	11.723 8.108 11.755 8.172 ;
			RECT	11.891 8.108 11.923 8.172 ;
			RECT	12.059 8.108 12.091 8.172 ;
			RECT	12.227 8.108 12.259 8.172 ;
			RECT	12.395 8.108 12.427 8.172 ;
			RECT	12.563 8.108 12.595 8.172 ;
			RECT	12.731 8.108 12.763 8.172 ;
			RECT	12.899 8.108 12.931 8.172 ;
			RECT	13.067 8.108 13.099 8.172 ;
			RECT	13.235 8.108 13.267 8.172 ;
			RECT	13.403 8.108 13.435 8.172 ;
			RECT	13.571 8.108 13.603 8.172 ;
			RECT	13.739 8.108 13.771 8.172 ;
			RECT	13.907 8.108 13.939 8.172 ;
			RECT	14.075 8.108 14.107 8.172 ;
			RECT	14.243 8.108 14.275 8.172 ;
			RECT	14.411 8.108 14.443 8.172 ;
			RECT	14.579 8.108 14.611 8.172 ;
			RECT	14.747 8.108 14.779 8.172 ;
			RECT	14.915 8.108 14.947 8.172 ;
			RECT	15.083 8.108 15.115 8.172 ;
			RECT	15.251 8.108 15.283 8.172 ;
			RECT	15.419 8.108 15.451 8.172 ;
			RECT	15.587 8.108 15.619 8.172 ;
			RECT	15.755 8.108 15.787 8.172 ;
			RECT	15.923 8.108 15.955 8.172 ;
			RECT	16.091 8.108 16.123 8.172 ;
			RECT	16.259 8.108 16.291 8.172 ;
			RECT	16.427 8.108 16.459 8.172 ;
			RECT	16.595 8.108 16.627 8.172 ;
			RECT	16.763 8.108 16.795 8.172 ;
			RECT	16.931 8.108 16.963 8.172 ;
			RECT	17.099 8.108 17.131 8.172 ;
			RECT	17.267 8.108 17.299 8.172 ;
			RECT	17.435 8.108 17.467 8.172 ;
			RECT	17.603 8.108 17.635 8.172 ;
			RECT	17.771 8.108 17.803 8.172 ;
			RECT	17.939 8.108 17.971 8.172 ;
			RECT	18.107 8.108 18.139 8.172 ;
			RECT	18.275 8.108 18.307 8.172 ;
			RECT	18.443 8.108 18.475 8.172 ;
			RECT	18.611 8.108 18.643 8.172 ;
			RECT	18.779 8.108 18.811 8.172 ;
			RECT	18.947 8.108 18.979 8.172 ;
			RECT	19.115 8.108 19.147 8.172 ;
			RECT	19.283 8.108 19.315 8.172 ;
			RECT	19.451 8.108 19.483 8.172 ;
			RECT	19.619 8.108 19.651 8.172 ;
			RECT	19.787 8.108 19.819 8.172 ;
			RECT	19.955 8.108 19.987 8.172 ;
			RECT	20.123 8.108 20.155 8.172 ;
			RECT	20.291 8.108 20.323 8.172 ;
			RECT	20.459 8.108 20.491 8.172 ;
			RECT	20.627 8.108 20.659 8.172 ;
			RECT	20.795 8.108 20.827 8.172 ;
			RECT	20.963 8.108 20.995 8.172 ;
			RECT	21.131 8.108 21.163 8.172 ;
			RECT	21.299 8.108 21.331 8.172 ;
			RECT	21.467 8.108 21.499 8.172 ;
			RECT	21.635 8.108 21.667 8.172 ;
			RECT	21.803 8.108 21.835 8.172 ;
			RECT	21.971 8.108 22.003 8.172 ;
			RECT	22.139 8.108 22.171 8.172 ;
			RECT	22.307 8.108 22.339 8.172 ;
			RECT	22.475 8.108 22.507 8.172 ;
			RECT	22.643 8.108 22.675 8.172 ;
			RECT	22.811 8.108 22.843 8.172 ;
			RECT	22.979 8.108 23.011 8.172 ;
			RECT	23.147 8.108 23.179 8.172 ;
			RECT	23.315 8.108 23.347 8.172 ;
			RECT	23.483 8.108 23.515 8.172 ;
			RECT	23.651 8.108 23.683 8.172 ;
			RECT	23.819 8.108 23.851 8.172 ;
			RECT	23.987 8.108 24.019 8.172 ;
			RECT	24.155 8.108 24.187 8.172 ;
			RECT	24.323 8.108 24.355 8.172 ;
			RECT	24.491 8.108 24.523 8.172 ;
			RECT	24.659 8.108 24.691 8.172 ;
			RECT	24.827 8.108 24.859 8.172 ;
			RECT	24.995 8.108 25.027 8.172 ;
			RECT	25.163 8.108 25.195 8.172 ;
			RECT	25.331 8.108 25.363 8.172 ;
			RECT	25.499 8.108 25.531 8.172 ;
			RECT	25.667 8.108 25.699 8.172 ;
			RECT	25.835 8.108 25.867 8.172 ;
			RECT	26.003 8.108 26.035 8.172 ;
			RECT	26.171 8.108 26.203 8.172 ;
			RECT	26.339 8.108 26.371 8.172 ;
			RECT	26.507 8.108 26.539 8.172 ;
			RECT	26.675 8.108 26.707 8.172 ;
			RECT	26.843 8.108 26.875 8.172 ;
			RECT	27.011 8.108 27.043 8.172 ;
			RECT	27.179 8.108 27.211 8.172 ;
			RECT	27.347 8.108 27.379 8.172 ;
			RECT	27.515 8.108 27.547 8.172 ;
			RECT	27.683 8.108 27.715 8.172 ;
			RECT	27.851 8.108 27.883 8.172 ;
			RECT	28.019 8.108 28.051 8.172 ;
			RECT	28.187 8.108 28.219 8.172 ;
			RECT	28.355 8.108 28.387 8.172 ;
			RECT	28.523 8.108 28.555 8.172 ;
			RECT	28.691 8.108 28.723 8.172 ;
			RECT	28.859 8.108 28.891 8.172 ;
			RECT	29.027 8.108 29.059 8.172 ;
			RECT	29.195 8.108 29.227 8.172 ;
			RECT	29.363 8.108 29.395 8.172 ;
			RECT	29.531 8.108 29.563 8.172 ;
			RECT	29.699 8.108 29.731 8.172 ;
			RECT	29.867 8.108 29.899 8.172 ;
			RECT	30.035 8.108 30.067 8.172 ;
			RECT	30.203 8.108 30.235 8.172 ;
			RECT	30.371 8.108 30.403 8.172 ;
			RECT	30.539 8.108 30.571 8.172 ;
			RECT	30.707 8.108 30.739 8.172 ;
			RECT	30.875 8.108 30.907 8.172 ;
			RECT	31.043 8.108 31.075 8.172 ;
			RECT	31.211 8.108 31.243 8.172 ;
			RECT	31.379 8.108 31.411 8.172 ;
			RECT	31.547 8.108 31.579 8.172 ;
			RECT	31.715 8.108 31.747 8.172 ;
			RECT	31.883 8.108 31.915 8.172 ;
			RECT	32.051 8.108 32.083 8.172 ;
			RECT	32.219 8.108 32.251 8.172 ;
			RECT	32.387 8.108 32.419 8.172 ;
			RECT	32.555 8.108 32.587 8.172 ;
			RECT	32.723 8.108 32.755 8.172 ;
			RECT	32.891 8.108 32.923 8.172 ;
			RECT	33.059 8.108 33.091 8.172 ;
			RECT	33.227 8.108 33.259 8.172 ;
			RECT	33.395 8.108 33.427 8.172 ;
			RECT	33.563 8.108 33.595 8.172 ;
			RECT	33.731 8.108 33.763 8.172 ;
			RECT	33.899 8.108 33.931 8.172 ;
			RECT	34.067 8.108 34.099 8.172 ;
			RECT	34.235 8.108 34.267 8.172 ;
			RECT	34.403 8.108 34.435 8.172 ;
			RECT	34.571 8.108 34.603 8.172 ;
			RECT	34.739 8.108 34.771 8.172 ;
			RECT	34.907 8.108 34.939 8.172 ;
			RECT	35.075 8.108 35.107 8.172 ;
			RECT	35.243 8.108 35.275 8.172 ;
			RECT	35.411 8.108 35.443 8.172 ;
			RECT	35.579 8.108 35.611 8.172 ;
			RECT	35.747 8.108 35.779 8.172 ;
			RECT	35.915 8.108 35.947 8.172 ;
			RECT	36.083 8.108 36.115 8.172 ;
			RECT	36.251 8.108 36.283 8.172 ;
			RECT	36.419 8.108 36.451 8.172 ;
			RECT	36.587 8.108 36.619 8.172 ;
			RECT	36.755 8.108 36.787 8.172 ;
			RECT	36.923 8.108 36.955 8.172 ;
			RECT	37.091 8.108 37.123 8.172 ;
			RECT	37.259 8.108 37.291 8.172 ;
			RECT	37.427 8.108 37.459 8.172 ;
			RECT	37.595 8.108 37.627 8.172 ;
			RECT	37.763 8.108 37.795 8.172 ;
			RECT	37.931 8.108 37.963 8.172 ;
			RECT	38.099 8.108 38.131 8.172 ;
			RECT	38.267 8.108 38.299 8.172 ;
			RECT	38.435 8.108 38.467 8.172 ;
			RECT	38.603 8.108 38.635 8.172 ;
			RECT	38.771 8.108 38.803 8.172 ;
			RECT	38.939 8.108 38.971 8.172 ;
			RECT	39.107 8.108 39.139 8.172 ;
			RECT	39.275 8.108 39.307 8.172 ;
			RECT	39.443 8.108 39.475 8.172 ;
			RECT	39.611 8.108 39.643 8.172 ;
			RECT	39.779 8.108 39.811 8.172 ;
			RECT	39.947 8.108 39.979 8.172 ;
			RECT	40.115 8.108 40.147 8.172 ;
			RECT	40.283 8.108 40.315 8.172 ;
			RECT	40.451 8.108 40.483 8.172 ;
			RECT	40.619 8.108 40.651 8.172 ;
			RECT	40.787 8.108 40.819 8.172 ;
			RECT	40.955 8.108 40.987 8.172 ;
			RECT	41.123 8.108 41.155 8.172 ;
			RECT	41.291 8.108 41.323 8.172 ;
			RECT	41.459 8.108 41.491 8.172 ;
			RECT	41.627 8.108 41.659 8.172 ;
			RECT	41.795 8.108 41.827 8.172 ;
			RECT	41.963 8.108 41.995 8.172 ;
			RECT	42.131 8.108 42.163 8.172 ;
			RECT	42.299 8.108 42.331 8.172 ;
			RECT	42.467 8.108 42.499 8.172 ;
			RECT	42.635 8.108 42.667 8.172 ;
			RECT	42.803 8.108 42.835 8.172 ;
			RECT	42.971 8.108 43.003 8.172 ;
			RECT	43.139 8.108 43.171 8.172 ;
			RECT	43.307 8.108 43.339 8.172 ;
			RECT	43.475 8.108 43.507 8.172 ;
			RECT	43.643 8.108 43.675 8.172 ;
			RECT	43.811 8.108 43.843 8.172 ;
			RECT	43.979 8.108 44.011 8.172 ;
			RECT	44.147 8.108 44.179 8.172 ;
			RECT	44.315 8.108 44.347 8.172 ;
			RECT	44.483 8.108 44.515 8.172 ;
			RECT	44.651 8.108 44.683 8.172 ;
			RECT	44.819 8.108 44.851 8.172 ;
			RECT	44.987 8.108 45.019 8.172 ;
			RECT	45.155 8.108 45.187 8.172 ;
			RECT	45.323 8.108 45.355 8.172 ;
			RECT	45.491 8.108 45.523 8.172 ;
			RECT	45.659 8.108 45.691 8.172 ;
			RECT	45.827 8.108 45.859 8.172 ;
			RECT	45.995 8.108 46.027 8.172 ;
			RECT	46.163 8.108 46.195 8.172 ;
			RECT	46.331 8.108 46.363 8.172 ;
			RECT	46.499 8.108 46.531 8.172 ;
			RECT	46.667 8.108 46.699 8.172 ;
			RECT	46.835 8.108 46.867 8.172 ;
			RECT	47.003 8.108 47.035 8.172 ;
			RECT	47.171 8.108 47.203 8.172 ;
			RECT	47.339 8.108 47.371 8.172 ;
			RECT	47.507 8.108 47.539 8.172 ;
			RECT	47.675 8.108 47.707 8.172 ;
			RECT	47.843 8.108 47.875 8.172 ;
			RECT	48.011 8.108 48.043 8.172 ;
			RECT	48.179 8.108 48.211 8.172 ;
			RECT	48.347 8.108 48.379 8.172 ;
			RECT	48.515 8.108 48.547 8.172 ;
			RECT	48.683 8.108 48.715 8.172 ;
			RECT	48.851 8.108 48.883 8.172 ;
			RECT	49.019 8.108 49.051 8.172 ;
			RECT	49.187 8.108 49.219 8.172 ;
			RECT	49.318 8.124 49.35 8.156 ;
			RECT	49.439 8.124 49.471 8.156 ;
			RECT	49.569 8.108 49.601 8.172 ;
			RECT	51.881 8.108 51.913 8.172 ;
			RECT	53.132 8.108 53.196 8.172 ;
			RECT	53.812 8.108 53.844 8.172 ;
			RECT	54.251 8.108 54.283 8.172 ;
			RECT	55.562 8.108 55.626 8.172 ;
			RECT	58.603 8.108 58.635 8.172 ;
			RECT	58.733 8.124 58.765 8.156 ;
			RECT	58.854 8.124 58.886 8.156 ;
			RECT	58.985 8.108 59.017 8.172 ;
			RECT	59.153 8.108 59.185 8.172 ;
			RECT	59.321 8.108 59.353 8.172 ;
			RECT	59.489 8.108 59.521 8.172 ;
			RECT	59.657 8.108 59.689 8.172 ;
			RECT	59.825 8.108 59.857 8.172 ;
			RECT	59.993 8.108 60.025 8.172 ;
			RECT	60.161 8.108 60.193 8.172 ;
			RECT	60.329 8.108 60.361 8.172 ;
			RECT	60.497 8.108 60.529 8.172 ;
			RECT	60.665 8.108 60.697 8.172 ;
			RECT	60.833 8.108 60.865 8.172 ;
			RECT	61.001 8.108 61.033 8.172 ;
			RECT	61.169 8.108 61.201 8.172 ;
			RECT	61.337 8.108 61.369 8.172 ;
			RECT	61.505 8.108 61.537 8.172 ;
			RECT	61.673 8.108 61.705 8.172 ;
			RECT	61.841 8.108 61.873 8.172 ;
			RECT	62.009 8.108 62.041 8.172 ;
			RECT	62.177 8.108 62.209 8.172 ;
			RECT	62.345 8.108 62.377 8.172 ;
			RECT	62.513 8.108 62.545 8.172 ;
			RECT	62.681 8.108 62.713 8.172 ;
			RECT	62.849 8.108 62.881 8.172 ;
			RECT	63.017 8.108 63.049 8.172 ;
			RECT	63.185 8.108 63.217 8.172 ;
			RECT	63.353 8.108 63.385 8.172 ;
			RECT	63.521 8.108 63.553 8.172 ;
			RECT	63.689 8.108 63.721 8.172 ;
			RECT	63.857 8.108 63.889 8.172 ;
			RECT	64.025 8.108 64.057 8.172 ;
			RECT	64.193 8.108 64.225 8.172 ;
			RECT	64.361 8.108 64.393 8.172 ;
			RECT	64.529 8.108 64.561 8.172 ;
			RECT	64.697 8.108 64.729 8.172 ;
			RECT	64.865 8.108 64.897 8.172 ;
			RECT	65.033 8.108 65.065 8.172 ;
			RECT	65.201 8.108 65.233 8.172 ;
			RECT	65.369 8.108 65.401 8.172 ;
			RECT	65.537 8.108 65.569 8.172 ;
			RECT	65.705 8.108 65.737 8.172 ;
			RECT	65.873 8.108 65.905 8.172 ;
			RECT	66.041 8.108 66.073 8.172 ;
			RECT	66.209 8.108 66.241 8.172 ;
			RECT	66.377 8.108 66.409 8.172 ;
			RECT	66.545 8.108 66.577 8.172 ;
			RECT	66.713 8.108 66.745 8.172 ;
			RECT	66.881 8.108 66.913 8.172 ;
			RECT	67.049 8.108 67.081 8.172 ;
			RECT	67.217 8.108 67.249 8.172 ;
			RECT	67.385 8.108 67.417 8.172 ;
			RECT	67.553 8.108 67.585 8.172 ;
			RECT	67.721 8.108 67.753 8.172 ;
			RECT	67.889 8.108 67.921 8.172 ;
			RECT	68.057 8.108 68.089 8.172 ;
			RECT	68.225 8.108 68.257 8.172 ;
			RECT	68.393 8.108 68.425 8.172 ;
			RECT	68.561 8.108 68.593 8.172 ;
			RECT	68.729 8.108 68.761 8.172 ;
			RECT	68.897 8.108 68.929 8.172 ;
			RECT	69.065 8.108 69.097 8.172 ;
			RECT	69.233 8.108 69.265 8.172 ;
			RECT	69.401 8.108 69.433 8.172 ;
			RECT	69.569 8.108 69.601 8.172 ;
			RECT	69.737 8.108 69.769 8.172 ;
			RECT	69.905 8.108 69.937 8.172 ;
			RECT	70.073 8.108 70.105 8.172 ;
			RECT	70.241 8.108 70.273 8.172 ;
			RECT	70.409 8.108 70.441 8.172 ;
			RECT	70.577 8.108 70.609 8.172 ;
			RECT	70.745 8.108 70.777 8.172 ;
			RECT	70.913 8.108 70.945 8.172 ;
			RECT	71.081 8.108 71.113 8.172 ;
			RECT	71.249 8.108 71.281 8.172 ;
			RECT	71.417 8.108 71.449 8.172 ;
			RECT	71.585 8.108 71.617 8.172 ;
			RECT	71.753 8.108 71.785 8.172 ;
			RECT	71.921 8.108 71.953 8.172 ;
			RECT	72.089 8.108 72.121 8.172 ;
			RECT	72.257 8.108 72.289 8.172 ;
			RECT	72.425 8.108 72.457 8.172 ;
			RECT	72.593 8.108 72.625 8.172 ;
			RECT	72.761 8.108 72.793 8.172 ;
			RECT	72.929 8.108 72.961 8.172 ;
			RECT	73.097 8.108 73.129 8.172 ;
			RECT	73.265 8.108 73.297 8.172 ;
			RECT	73.433 8.108 73.465 8.172 ;
			RECT	73.601 8.108 73.633 8.172 ;
			RECT	73.769 8.108 73.801 8.172 ;
			RECT	73.937 8.108 73.969 8.172 ;
			RECT	74.105 8.108 74.137 8.172 ;
			RECT	74.273 8.108 74.305 8.172 ;
			RECT	74.441 8.108 74.473 8.172 ;
			RECT	74.609 8.108 74.641 8.172 ;
			RECT	74.777 8.108 74.809 8.172 ;
			RECT	74.945 8.108 74.977 8.172 ;
			RECT	75.113 8.108 75.145 8.172 ;
			RECT	75.281 8.108 75.313 8.172 ;
			RECT	75.449 8.108 75.481 8.172 ;
			RECT	75.617 8.108 75.649 8.172 ;
			RECT	75.785 8.108 75.817 8.172 ;
			RECT	75.953 8.108 75.985 8.172 ;
			RECT	76.121 8.108 76.153 8.172 ;
			RECT	76.289 8.108 76.321 8.172 ;
			RECT	76.457 8.108 76.489 8.172 ;
			RECT	76.625 8.108 76.657 8.172 ;
			RECT	76.793 8.108 76.825 8.172 ;
			RECT	76.961 8.108 76.993 8.172 ;
			RECT	77.129 8.108 77.161 8.172 ;
			RECT	77.297 8.108 77.329 8.172 ;
			RECT	77.465 8.108 77.497 8.172 ;
			RECT	77.633 8.108 77.665 8.172 ;
			RECT	77.801 8.108 77.833 8.172 ;
			RECT	77.969 8.108 78.001 8.172 ;
			RECT	78.137 8.108 78.169 8.172 ;
			RECT	78.305 8.108 78.337 8.172 ;
			RECT	78.473 8.108 78.505 8.172 ;
			RECT	78.641 8.108 78.673 8.172 ;
			RECT	78.809 8.108 78.841 8.172 ;
			RECT	78.977 8.108 79.009 8.172 ;
			RECT	79.145 8.108 79.177 8.172 ;
			RECT	79.313 8.108 79.345 8.172 ;
			RECT	79.481 8.108 79.513 8.172 ;
			RECT	79.649 8.108 79.681 8.172 ;
			RECT	79.817 8.108 79.849 8.172 ;
			RECT	79.985 8.108 80.017 8.172 ;
			RECT	80.153 8.108 80.185 8.172 ;
			RECT	80.321 8.108 80.353 8.172 ;
			RECT	80.489 8.108 80.521 8.172 ;
			RECT	80.657 8.108 80.689 8.172 ;
			RECT	80.825 8.108 80.857 8.172 ;
			RECT	80.993 8.108 81.025 8.172 ;
			RECT	81.161 8.108 81.193 8.172 ;
			RECT	81.329 8.108 81.361 8.172 ;
			RECT	81.497 8.108 81.529 8.172 ;
			RECT	81.665 8.108 81.697 8.172 ;
			RECT	81.833 8.108 81.865 8.172 ;
			RECT	82.001 8.108 82.033 8.172 ;
			RECT	82.169 8.108 82.201 8.172 ;
			RECT	82.337 8.108 82.369 8.172 ;
			RECT	82.505 8.108 82.537 8.172 ;
			RECT	82.673 8.108 82.705 8.172 ;
			RECT	82.841 8.108 82.873 8.172 ;
			RECT	83.009 8.108 83.041 8.172 ;
			RECT	83.177 8.108 83.209 8.172 ;
			RECT	83.345 8.108 83.377 8.172 ;
			RECT	83.513 8.108 83.545 8.172 ;
			RECT	83.681 8.108 83.713 8.172 ;
			RECT	83.849 8.108 83.881 8.172 ;
			RECT	84.017 8.108 84.049 8.172 ;
			RECT	84.185 8.108 84.217 8.172 ;
			RECT	84.353 8.108 84.385 8.172 ;
			RECT	84.521 8.108 84.553 8.172 ;
			RECT	84.689 8.108 84.721 8.172 ;
			RECT	84.857 8.108 84.889 8.172 ;
			RECT	85.025 8.108 85.057 8.172 ;
			RECT	85.193 8.108 85.225 8.172 ;
			RECT	85.361 8.108 85.393 8.172 ;
			RECT	85.529 8.108 85.561 8.172 ;
			RECT	85.697 8.108 85.729 8.172 ;
			RECT	85.865 8.108 85.897 8.172 ;
			RECT	86.033 8.108 86.065 8.172 ;
			RECT	86.201 8.108 86.233 8.172 ;
			RECT	86.369 8.108 86.401 8.172 ;
			RECT	86.537 8.108 86.569 8.172 ;
			RECT	86.705 8.108 86.737 8.172 ;
			RECT	86.873 8.108 86.905 8.172 ;
			RECT	87.041 8.108 87.073 8.172 ;
			RECT	87.209 8.108 87.241 8.172 ;
			RECT	87.377 8.108 87.409 8.172 ;
			RECT	87.545 8.108 87.577 8.172 ;
			RECT	87.713 8.108 87.745 8.172 ;
			RECT	87.881 8.108 87.913 8.172 ;
			RECT	88.049 8.108 88.081 8.172 ;
			RECT	88.217 8.108 88.249 8.172 ;
			RECT	88.385 8.108 88.417 8.172 ;
			RECT	88.553 8.108 88.585 8.172 ;
			RECT	88.721 8.108 88.753 8.172 ;
			RECT	88.889 8.108 88.921 8.172 ;
			RECT	89.057 8.108 89.089 8.172 ;
			RECT	89.225 8.108 89.257 8.172 ;
			RECT	89.393 8.108 89.425 8.172 ;
			RECT	89.561 8.108 89.593 8.172 ;
			RECT	89.729 8.108 89.761 8.172 ;
			RECT	89.897 8.108 89.929 8.172 ;
			RECT	90.065 8.108 90.097 8.172 ;
			RECT	90.233 8.108 90.265 8.172 ;
			RECT	90.401 8.108 90.433 8.172 ;
			RECT	90.569 8.108 90.601 8.172 ;
			RECT	90.737 8.108 90.769 8.172 ;
			RECT	90.905 8.108 90.937 8.172 ;
			RECT	91.073 8.108 91.105 8.172 ;
			RECT	91.241 8.108 91.273 8.172 ;
			RECT	91.409 8.108 91.441 8.172 ;
			RECT	91.577 8.108 91.609 8.172 ;
			RECT	91.745 8.108 91.777 8.172 ;
			RECT	91.913 8.108 91.945 8.172 ;
			RECT	92.081 8.108 92.113 8.172 ;
			RECT	92.249 8.108 92.281 8.172 ;
			RECT	92.417 8.108 92.449 8.172 ;
			RECT	92.585 8.108 92.617 8.172 ;
			RECT	92.753 8.108 92.785 8.172 ;
			RECT	92.921 8.108 92.953 8.172 ;
			RECT	93.089 8.108 93.121 8.172 ;
			RECT	93.257 8.108 93.289 8.172 ;
			RECT	93.425 8.108 93.457 8.172 ;
			RECT	93.593 8.108 93.625 8.172 ;
			RECT	93.761 8.108 93.793 8.172 ;
			RECT	93.929 8.108 93.961 8.172 ;
			RECT	94.097 8.108 94.129 8.172 ;
			RECT	94.265 8.108 94.297 8.172 ;
			RECT	94.433 8.108 94.465 8.172 ;
			RECT	94.601 8.108 94.633 8.172 ;
			RECT	94.769 8.108 94.801 8.172 ;
			RECT	94.937 8.108 94.969 8.172 ;
			RECT	95.105 8.108 95.137 8.172 ;
			RECT	95.273 8.108 95.305 8.172 ;
			RECT	95.441 8.108 95.473 8.172 ;
			RECT	95.609 8.108 95.641 8.172 ;
			RECT	95.777 8.108 95.809 8.172 ;
			RECT	95.945 8.108 95.977 8.172 ;
			RECT	96.113 8.108 96.145 8.172 ;
			RECT	96.281 8.108 96.313 8.172 ;
			RECT	96.449 8.108 96.481 8.172 ;
			RECT	96.617 8.108 96.649 8.172 ;
			RECT	96.785 8.108 96.817 8.172 ;
			RECT	96.953 8.108 96.985 8.172 ;
			RECT	97.121 8.108 97.153 8.172 ;
			RECT	97.289 8.108 97.321 8.172 ;
			RECT	97.457 8.108 97.489 8.172 ;
			RECT	97.625 8.108 97.657 8.172 ;
			RECT	97.793 8.108 97.825 8.172 ;
			RECT	97.961 8.108 97.993 8.172 ;
			RECT	98.129 8.108 98.161 8.172 ;
			RECT	98.297 8.108 98.329 8.172 ;
			RECT	98.465 8.108 98.497 8.172 ;
			RECT	98.633 8.108 98.665 8.172 ;
			RECT	98.801 8.108 98.833 8.172 ;
			RECT	98.969 8.108 99.001 8.172 ;
			RECT	99.137 8.108 99.169 8.172 ;
			RECT	99.305 8.108 99.337 8.172 ;
			RECT	99.473 8.108 99.505 8.172 ;
			RECT	99.641 8.108 99.673 8.172 ;
			RECT	99.809 8.108 99.841 8.172 ;
			RECT	99.977 8.108 100.009 8.172 ;
			RECT	100.145 8.108 100.177 8.172 ;
			RECT	100.313 8.108 100.345 8.172 ;
			RECT	100.481 8.108 100.513 8.172 ;
			RECT	100.649 8.108 100.681 8.172 ;
			RECT	100.817 8.108 100.849 8.172 ;
			RECT	100.985 8.108 101.017 8.172 ;
			RECT	101.153 8.108 101.185 8.172 ;
			RECT	101.321 8.108 101.353 8.172 ;
			RECT	101.489 8.108 101.521 8.172 ;
			RECT	101.657 8.108 101.689 8.172 ;
			RECT	101.825 8.108 101.857 8.172 ;
			RECT	101.993 8.108 102.025 8.172 ;
			RECT	102.123 8.124 102.155 8.156 ;
			RECT	102.245 8.129 102.277 8.161 ;
			RECT	102.375 8.108 102.407 8.172 ;
			RECT	103.795 8.108 103.827 8.172 ;
			RECT	103.925 8.129 103.957 8.161 ;
			RECT	104.047 8.124 104.079 8.156 ;
			RECT	104.177 8.108 104.209 8.172 ;
			RECT	104.345 8.108 104.377 8.172 ;
			RECT	104.513 8.108 104.545 8.172 ;
			RECT	104.681 8.108 104.713 8.172 ;
			RECT	104.849 8.108 104.881 8.172 ;
			RECT	105.017 8.108 105.049 8.172 ;
			RECT	105.185 8.108 105.217 8.172 ;
			RECT	105.353 8.108 105.385 8.172 ;
			RECT	105.521 8.108 105.553 8.172 ;
			RECT	105.689 8.108 105.721 8.172 ;
			RECT	105.857 8.108 105.889 8.172 ;
			RECT	106.025 8.108 106.057 8.172 ;
			RECT	106.193 8.108 106.225 8.172 ;
			RECT	106.361 8.108 106.393 8.172 ;
			RECT	106.529 8.108 106.561 8.172 ;
			RECT	106.697 8.108 106.729 8.172 ;
			RECT	106.865 8.108 106.897 8.172 ;
			RECT	107.033 8.108 107.065 8.172 ;
			RECT	107.201 8.108 107.233 8.172 ;
			RECT	107.369 8.108 107.401 8.172 ;
			RECT	107.537 8.108 107.569 8.172 ;
			RECT	107.705 8.108 107.737 8.172 ;
			RECT	107.873 8.108 107.905 8.172 ;
			RECT	108.041 8.108 108.073 8.172 ;
			RECT	108.209 8.108 108.241 8.172 ;
			RECT	108.377 8.108 108.409 8.172 ;
			RECT	108.545 8.108 108.577 8.172 ;
			RECT	108.713 8.108 108.745 8.172 ;
			RECT	108.881 8.108 108.913 8.172 ;
			RECT	109.049 8.108 109.081 8.172 ;
			RECT	109.217 8.108 109.249 8.172 ;
			RECT	109.385 8.108 109.417 8.172 ;
			RECT	109.553 8.108 109.585 8.172 ;
			RECT	109.721 8.108 109.753 8.172 ;
			RECT	109.889 8.108 109.921 8.172 ;
			RECT	110.057 8.108 110.089 8.172 ;
			RECT	110.225 8.108 110.257 8.172 ;
			RECT	110.393 8.108 110.425 8.172 ;
			RECT	110.561 8.108 110.593 8.172 ;
			RECT	110.729 8.108 110.761 8.172 ;
			RECT	110.897 8.108 110.929 8.172 ;
			RECT	111.065 8.108 111.097 8.172 ;
			RECT	111.233 8.108 111.265 8.172 ;
			RECT	111.401 8.108 111.433 8.172 ;
			RECT	111.569 8.108 111.601 8.172 ;
			RECT	111.737 8.108 111.769 8.172 ;
			RECT	111.905 8.108 111.937 8.172 ;
			RECT	112.073 8.108 112.105 8.172 ;
			RECT	112.241 8.108 112.273 8.172 ;
			RECT	112.409 8.108 112.441 8.172 ;
			RECT	112.577 8.108 112.609 8.172 ;
			RECT	112.745 8.108 112.777 8.172 ;
			RECT	112.913 8.108 112.945 8.172 ;
			RECT	113.081 8.108 113.113 8.172 ;
			RECT	113.249 8.108 113.281 8.172 ;
			RECT	113.417 8.108 113.449 8.172 ;
			RECT	113.585 8.108 113.617 8.172 ;
			RECT	113.753 8.108 113.785 8.172 ;
			RECT	113.921 8.108 113.953 8.172 ;
			RECT	114.089 8.108 114.121 8.172 ;
			RECT	114.257 8.108 114.289 8.172 ;
			RECT	114.425 8.108 114.457 8.172 ;
			RECT	114.593 8.108 114.625 8.172 ;
			RECT	114.761 8.108 114.793 8.172 ;
			RECT	114.929 8.108 114.961 8.172 ;
			RECT	115.097 8.108 115.129 8.172 ;
			RECT	115.265 8.108 115.297 8.172 ;
			RECT	115.433 8.108 115.465 8.172 ;
			RECT	115.601 8.108 115.633 8.172 ;
			RECT	115.769 8.108 115.801 8.172 ;
			RECT	115.937 8.108 115.969 8.172 ;
			RECT	116.105 8.108 116.137 8.172 ;
			RECT	116.273 8.108 116.305 8.172 ;
			RECT	116.441 8.108 116.473 8.172 ;
			RECT	116.609 8.108 116.641 8.172 ;
			RECT	116.777 8.108 116.809 8.172 ;
			RECT	116.945 8.108 116.977 8.172 ;
			RECT	117.113 8.108 117.145 8.172 ;
			RECT	117.281 8.108 117.313 8.172 ;
			RECT	117.449 8.108 117.481 8.172 ;
			RECT	117.617 8.108 117.649 8.172 ;
			RECT	117.785 8.108 117.817 8.172 ;
			RECT	117.953 8.108 117.985 8.172 ;
			RECT	118.121 8.108 118.153 8.172 ;
			RECT	118.289 8.108 118.321 8.172 ;
			RECT	118.457 8.108 118.489 8.172 ;
			RECT	118.625 8.108 118.657 8.172 ;
			RECT	118.793 8.108 118.825 8.172 ;
			RECT	118.961 8.108 118.993 8.172 ;
			RECT	119.129 8.108 119.161 8.172 ;
			RECT	119.297 8.108 119.329 8.172 ;
			RECT	119.465 8.108 119.497 8.172 ;
			RECT	119.633 8.108 119.665 8.172 ;
			RECT	119.801 8.108 119.833 8.172 ;
			RECT	119.969 8.108 120.001 8.172 ;
			RECT	120.137 8.108 120.169 8.172 ;
			RECT	120.305 8.108 120.337 8.172 ;
			RECT	120.473 8.108 120.505 8.172 ;
			RECT	120.641 8.108 120.673 8.172 ;
			RECT	120.809 8.108 120.841 8.172 ;
			RECT	120.977 8.108 121.009 8.172 ;
			RECT	121.145 8.108 121.177 8.172 ;
			RECT	121.313 8.108 121.345 8.172 ;
			RECT	121.481 8.108 121.513 8.172 ;
			RECT	121.649 8.108 121.681 8.172 ;
			RECT	121.817 8.108 121.849 8.172 ;
			RECT	121.985 8.108 122.017 8.172 ;
			RECT	122.153 8.108 122.185 8.172 ;
			RECT	122.321 8.108 122.353 8.172 ;
			RECT	122.489 8.108 122.521 8.172 ;
			RECT	122.657 8.108 122.689 8.172 ;
			RECT	122.825 8.108 122.857 8.172 ;
			RECT	122.993 8.108 123.025 8.172 ;
			RECT	123.161 8.108 123.193 8.172 ;
			RECT	123.329 8.108 123.361 8.172 ;
			RECT	123.497 8.108 123.529 8.172 ;
			RECT	123.665 8.108 123.697 8.172 ;
			RECT	123.833 8.108 123.865 8.172 ;
			RECT	124.001 8.108 124.033 8.172 ;
			RECT	124.169 8.108 124.201 8.172 ;
			RECT	124.337 8.108 124.369 8.172 ;
			RECT	124.505 8.108 124.537 8.172 ;
			RECT	124.673 8.108 124.705 8.172 ;
			RECT	124.841 8.108 124.873 8.172 ;
			RECT	125.009 8.108 125.041 8.172 ;
			RECT	125.177 8.108 125.209 8.172 ;
			RECT	125.345 8.108 125.377 8.172 ;
			RECT	125.513 8.108 125.545 8.172 ;
			RECT	125.681 8.108 125.713 8.172 ;
			RECT	125.849 8.108 125.881 8.172 ;
			RECT	126.017 8.108 126.049 8.172 ;
			RECT	126.185 8.108 126.217 8.172 ;
			RECT	126.353 8.108 126.385 8.172 ;
			RECT	126.521 8.108 126.553 8.172 ;
			RECT	126.689 8.108 126.721 8.172 ;
			RECT	126.857 8.108 126.889 8.172 ;
			RECT	127.025 8.108 127.057 8.172 ;
			RECT	127.193 8.108 127.225 8.172 ;
			RECT	127.361 8.108 127.393 8.172 ;
			RECT	127.529 8.108 127.561 8.172 ;
			RECT	127.697 8.108 127.729 8.172 ;
			RECT	127.865 8.108 127.897 8.172 ;
			RECT	128.033 8.108 128.065 8.172 ;
			RECT	128.201 8.108 128.233 8.172 ;
			RECT	128.369 8.108 128.401 8.172 ;
			RECT	128.537 8.108 128.569 8.172 ;
			RECT	128.705 8.108 128.737 8.172 ;
			RECT	128.873 8.108 128.905 8.172 ;
			RECT	129.041 8.108 129.073 8.172 ;
			RECT	129.209 8.108 129.241 8.172 ;
			RECT	129.377 8.108 129.409 8.172 ;
			RECT	129.545 8.108 129.577 8.172 ;
			RECT	129.713 8.108 129.745 8.172 ;
			RECT	129.881 8.108 129.913 8.172 ;
			RECT	130.049 8.108 130.081 8.172 ;
			RECT	130.217 8.108 130.249 8.172 ;
			RECT	130.385 8.108 130.417 8.172 ;
			RECT	130.553 8.108 130.585 8.172 ;
			RECT	130.721 8.108 130.753 8.172 ;
			RECT	130.889 8.108 130.921 8.172 ;
			RECT	131.057 8.108 131.089 8.172 ;
			RECT	131.225 8.108 131.257 8.172 ;
			RECT	131.393 8.108 131.425 8.172 ;
			RECT	131.561 8.108 131.593 8.172 ;
			RECT	131.729 8.108 131.761 8.172 ;
			RECT	131.897 8.108 131.929 8.172 ;
			RECT	132.065 8.108 132.097 8.172 ;
			RECT	132.233 8.108 132.265 8.172 ;
			RECT	132.401 8.108 132.433 8.172 ;
			RECT	132.569 8.108 132.601 8.172 ;
			RECT	132.737 8.108 132.769 8.172 ;
			RECT	132.905 8.108 132.937 8.172 ;
			RECT	133.073 8.108 133.105 8.172 ;
			RECT	133.241 8.108 133.273 8.172 ;
			RECT	133.409 8.108 133.441 8.172 ;
			RECT	133.577 8.108 133.609 8.172 ;
			RECT	133.745 8.108 133.777 8.172 ;
			RECT	133.913 8.108 133.945 8.172 ;
			RECT	134.081 8.108 134.113 8.172 ;
			RECT	134.249 8.108 134.281 8.172 ;
			RECT	134.417 8.108 134.449 8.172 ;
			RECT	134.585 8.108 134.617 8.172 ;
			RECT	134.753 8.108 134.785 8.172 ;
			RECT	134.921 8.108 134.953 8.172 ;
			RECT	135.089 8.108 135.121 8.172 ;
			RECT	135.257 8.108 135.289 8.172 ;
			RECT	135.425 8.108 135.457 8.172 ;
			RECT	135.593 8.108 135.625 8.172 ;
			RECT	135.761 8.108 135.793 8.172 ;
			RECT	135.929 8.108 135.961 8.172 ;
			RECT	136.097 8.108 136.129 8.172 ;
			RECT	136.265 8.108 136.297 8.172 ;
			RECT	136.433 8.108 136.465 8.172 ;
			RECT	136.601 8.108 136.633 8.172 ;
			RECT	136.769 8.108 136.801 8.172 ;
			RECT	136.937 8.108 136.969 8.172 ;
			RECT	137.105 8.108 137.137 8.172 ;
			RECT	137.273 8.108 137.305 8.172 ;
			RECT	137.441 8.108 137.473 8.172 ;
			RECT	137.609 8.108 137.641 8.172 ;
			RECT	137.777 8.108 137.809 8.172 ;
			RECT	137.945 8.108 137.977 8.172 ;
			RECT	138.113 8.108 138.145 8.172 ;
			RECT	138.281 8.108 138.313 8.172 ;
			RECT	138.449 8.108 138.481 8.172 ;
			RECT	138.617 8.108 138.649 8.172 ;
			RECT	138.785 8.108 138.817 8.172 ;
			RECT	138.953 8.108 138.985 8.172 ;
			RECT	139.121 8.108 139.153 8.172 ;
			RECT	139.289 8.108 139.321 8.172 ;
			RECT	139.457 8.108 139.489 8.172 ;
			RECT	139.625 8.108 139.657 8.172 ;
			RECT	139.793 8.108 139.825 8.172 ;
			RECT	139.961 8.108 139.993 8.172 ;
			RECT	140.129 8.108 140.161 8.172 ;
			RECT	140.297 8.108 140.329 8.172 ;
			RECT	140.465 8.108 140.497 8.172 ;
			RECT	140.633 8.108 140.665 8.172 ;
			RECT	140.801 8.108 140.833 8.172 ;
			RECT	140.969 8.108 141.001 8.172 ;
			RECT	141.137 8.108 141.169 8.172 ;
			RECT	141.305 8.108 141.337 8.172 ;
			RECT	141.473 8.108 141.505 8.172 ;
			RECT	141.641 8.108 141.673 8.172 ;
			RECT	141.809 8.108 141.841 8.172 ;
			RECT	141.977 8.108 142.009 8.172 ;
			RECT	142.145 8.108 142.177 8.172 ;
			RECT	142.313 8.108 142.345 8.172 ;
			RECT	142.481 8.108 142.513 8.172 ;
			RECT	142.649 8.108 142.681 8.172 ;
			RECT	142.817 8.108 142.849 8.172 ;
			RECT	142.985 8.108 143.017 8.172 ;
			RECT	143.153 8.108 143.185 8.172 ;
			RECT	143.321 8.108 143.353 8.172 ;
			RECT	143.489 8.108 143.521 8.172 ;
			RECT	143.657 8.108 143.689 8.172 ;
			RECT	143.825 8.108 143.857 8.172 ;
			RECT	143.993 8.108 144.025 8.172 ;
			RECT	144.161 8.108 144.193 8.172 ;
			RECT	144.329 8.108 144.361 8.172 ;
			RECT	144.497 8.108 144.529 8.172 ;
			RECT	144.665 8.108 144.697 8.172 ;
			RECT	144.833 8.108 144.865 8.172 ;
			RECT	145.001 8.108 145.033 8.172 ;
			RECT	145.169 8.108 145.201 8.172 ;
			RECT	145.337 8.108 145.369 8.172 ;
			RECT	145.505 8.108 145.537 8.172 ;
			RECT	145.673 8.108 145.705 8.172 ;
			RECT	145.841 8.108 145.873 8.172 ;
			RECT	146.009 8.108 146.041 8.172 ;
			RECT	146.177 8.108 146.209 8.172 ;
			RECT	146.345 8.108 146.377 8.172 ;
			RECT	146.513 8.108 146.545 8.172 ;
			RECT	146.681 8.108 146.713 8.172 ;
			RECT	146.849 8.108 146.881 8.172 ;
			RECT	147.017 8.108 147.049 8.172 ;
			RECT	147.185 8.108 147.217 8.172 ;
			RECT	147.316 8.124 147.348 8.156 ;
			RECT	147.437 8.124 147.469 8.156 ;
			RECT	147.567 8.108 147.599 8.172 ;
			RECT	149.879 8.108 149.911 8.172 ;
			RECT	151.13 8.108 151.194 8.172 ;
			RECT	151.81 8.108 151.842 8.172 ;
			RECT	152.249 8.108 152.281 8.172 ;
			RECT	153.56 8.108 153.624 8.172 ;
			RECT	156.601 8.108 156.633 8.172 ;
			RECT	156.731 8.124 156.763 8.156 ;
			RECT	156.852 8.124 156.884 8.156 ;
			RECT	156.983 8.108 157.015 8.172 ;
			RECT	157.151 8.108 157.183 8.172 ;
			RECT	157.319 8.108 157.351 8.172 ;
			RECT	157.487 8.108 157.519 8.172 ;
			RECT	157.655 8.108 157.687 8.172 ;
			RECT	157.823 8.108 157.855 8.172 ;
			RECT	157.991 8.108 158.023 8.172 ;
			RECT	158.159 8.108 158.191 8.172 ;
			RECT	158.327 8.108 158.359 8.172 ;
			RECT	158.495 8.108 158.527 8.172 ;
			RECT	158.663 8.108 158.695 8.172 ;
			RECT	158.831 8.108 158.863 8.172 ;
			RECT	158.999 8.108 159.031 8.172 ;
			RECT	159.167 8.108 159.199 8.172 ;
			RECT	159.335 8.108 159.367 8.172 ;
			RECT	159.503 8.108 159.535 8.172 ;
			RECT	159.671 8.108 159.703 8.172 ;
			RECT	159.839 8.108 159.871 8.172 ;
			RECT	160.007 8.108 160.039 8.172 ;
			RECT	160.175 8.108 160.207 8.172 ;
			RECT	160.343 8.108 160.375 8.172 ;
			RECT	160.511 8.108 160.543 8.172 ;
			RECT	160.679 8.108 160.711 8.172 ;
			RECT	160.847 8.108 160.879 8.172 ;
			RECT	161.015 8.108 161.047 8.172 ;
			RECT	161.183 8.108 161.215 8.172 ;
			RECT	161.351 8.108 161.383 8.172 ;
			RECT	161.519 8.108 161.551 8.172 ;
			RECT	161.687 8.108 161.719 8.172 ;
			RECT	161.855 8.108 161.887 8.172 ;
			RECT	162.023 8.108 162.055 8.172 ;
			RECT	162.191 8.108 162.223 8.172 ;
			RECT	162.359 8.108 162.391 8.172 ;
			RECT	162.527 8.108 162.559 8.172 ;
			RECT	162.695 8.108 162.727 8.172 ;
			RECT	162.863 8.108 162.895 8.172 ;
			RECT	163.031 8.108 163.063 8.172 ;
			RECT	163.199 8.108 163.231 8.172 ;
			RECT	163.367 8.108 163.399 8.172 ;
			RECT	163.535 8.108 163.567 8.172 ;
			RECT	163.703 8.108 163.735 8.172 ;
			RECT	163.871 8.108 163.903 8.172 ;
			RECT	164.039 8.108 164.071 8.172 ;
			RECT	164.207 8.108 164.239 8.172 ;
			RECT	164.375 8.108 164.407 8.172 ;
			RECT	164.543 8.108 164.575 8.172 ;
			RECT	164.711 8.108 164.743 8.172 ;
			RECT	164.879 8.108 164.911 8.172 ;
			RECT	165.047 8.108 165.079 8.172 ;
			RECT	165.215 8.108 165.247 8.172 ;
			RECT	165.383 8.108 165.415 8.172 ;
			RECT	165.551 8.108 165.583 8.172 ;
			RECT	165.719 8.108 165.751 8.172 ;
			RECT	165.887 8.108 165.919 8.172 ;
			RECT	166.055 8.108 166.087 8.172 ;
			RECT	166.223 8.108 166.255 8.172 ;
			RECT	166.391 8.108 166.423 8.172 ;
			RECT	166.559 8.108 166.591 8.172 ;
			RECT	166.727 8.108 166.759 8.172 ;
			RECT	166.895 8.108 166.927 8.172 ;
			RECT	167.063 8.108 167.095 8.172 ;
			RECT	167.231 8.108 167.263 8.172 ;
			RECT	167.399 8.108 167.431 8.172 ;
			RECT	167.567 8.108 167.599 8.172 ;
			RECT	167.735 8.108 167.767 8.172 ;
			RECT	167.903 8.108 167.935 8.172 ;
			RECT	168.071 8.108 168.103 8.172 ;
			RECT	168.239 8.108 168.271 8.172 ;
			RECT	168.407 8.108 168.439 8.172 ;
			RECT	168.575 8.108 168.607 8.172 ;
			RECT	168.743 8.108 168.775 8.172 ;
			RECT	168.911 8.108 168.943 8.172 ;
			RECT	169.079 8.108 169.111 8.172 ;
			RECT	169.247 8.108 169.279 8.172 ;
			RECT	169.415 8.108 169.447 8.172 ;
			RECT	169.583 8.108 169.615 8.172 ;
			RECT	169.751 8.108 169.783 8.172 ;
			RECT	169.919 8.108 169.951 8.172 ;
			RECT	170.087 8.108 170.119 8.172 ;
			RECT	170.255 8.108 170.287 8.172 ;
			RECT	170.423 8.108 170.455 8.172 ;
			RECT	170.591 8.108 170.623 8.172 ;
			RECT	170.759 8.108 170.791 8.172 ;
			RECT	170.927 8.108 170.959 8.172 ;
			RECT	171.095 8.108 171.127 8.172 ;
			RECT	171.263 8.108 171.295 8.172 ;
			RECT	171.431 8.108 171.463 8.172 ;
			RECT	171.599 8.108 171.631 8.172 ;
			RECT	171.767 8.108 171.799 8.172 ;
			RECT	171.935 8.108 171.967 8.172 ;
			RECT	172.103 8.108 172.135 8.172 ;
			RECT	172.271 8.108 172.303 8.172 ;
			RECT	172.439 8.108 172.471 8.172 ;
			RECT	172.607 8.108 172.639 8.172 ;
			RECT	172.775 8.108 172.807 8.172 ;
			RECT	172.943 8.108 172.975 8.172 ;
			RECT	173.111 8.108 173.143 8.172 ;
			RECT	173.279 8.108 173.311 8.172 ;
			RECT	173.447 8.108 173.479 8.172 ;
			RECT	173.615 8.108 173.647 8.172 ;
			RECT	173.783 8.108 173.815 8.172 ;
			RECT	173.951 8.108 173.983 8.172 ;
			RECT	174.119 8.108 174.151 8.172 ;
			RECT	174.287 8.108 174.319 8.172 ;
			RECT	174.455 8.108 174.487 8.172 ;
			RECT	174.623 8.108 174.655 8.172 ;
			RECT	174.791 8.108 174.823 8.172 ;
			RECT	174.959 8.108 174.991 8.172 ;
			RECT	175.127 8.108 175.159 8.172 ;
			RECT	175.295 8.108 175.327 8.172 ;
			RECT	175.463 8.108 175.495 8.172 ;
			RECT	175.631 8.108 175.663 8.172 ;
			RECT	175.799 8.108 175.831 8.172 ;
			RECT	175.967 8.108 175.999 8.172 ;
			RECT	176.135 8.108 176.167 8.172 ;
			RECT	176.303 8.108 176.335 8.172 ;
			RECT	176.471 8.108 176.503 8.172 ;
			RECT	176.639 8.108 176.671 8.172 ;
			RECT	176.807 8.108 176.839 8.172 ;
			RECT	176.975 8.108 177.007 8.172 ;
			RECT	177.143 8.108 177.175 8.172 ;
			RECT	177.311 8.108 177.343 8.172 ;
			RECT	177.479 8.108 177.511 8.172 ;
			RECT	177.647 8.108 177.679 8.172 ;
			RECT	177.815 8.108 177.847 8.172 ;
			RECT	177.983 8.108 178.015 8.172 ;
			RECT	178.151 8.108 178.183 8.172 ;
			RECT	178.319 8.108 178.351 8.172 ;
			RECT	178.487 8.108 178.519 8.172 ;
			RECT	178.655 8.108 178.687 8.172 ;
			RECT	178.823 8.108 178.855 8.172 ;
			RECT	178.991 8.108 179.023 8.172 ;
			RECT	179.159 8.108 179.191 8.172 ;
			RECT	179.327 8.108 179.359 8.172 ;
			RECT	179.495 8.108 179.527 8.172 ;
			RECT	179.663 8.108 179.695 8.172 ;
			RECT	179.831 8.108 179.863 8.172 ;
			RECT	179.999 8.108 180.031 8.172 ;
			RECT	180.167 8.108 180.199 8.172 ;
			RECT	180.335 8.108 180.367 8.172 ;
			RECT	180.503 8.108 180.535 8.172 ;
			RECT	180.671 8.108 180.703 8.172 ;
			RECT	180.839 8.108 180.871 8.172 ;
			RECT	181.007 8.108 181.039 8.172 ;
			RECT	181.175 8.108 181.207 8.172 ;
			RECT	181.343 8.108 181.375 8.172 ;
			RECT	181.511 8.108 181.543 8.172 ;
			RECT	181.679 8.108 181.711 8.172 ;
			RECT	181.847 8.108 181.879 8.172 ;
			RECT	182.015 8.108 182.047 8.172 ;
			RECT	182.183 8.108 182.215 8.172 ;
			RECT	182.351 8.108 182.383 8.172 ;
			RECT	182.519 8.108 182.551 8.172 ;
			RECT	182.687 8.108 182.719 8.172 ;
			RECT	182.855 8.108 182.887 8.172 ;
			RECT	183.023 8.108 183.055 8.172 ;
			RECT	183.191 8.108 183.223 8.172 ;
			RECT	183.359 8.108 183.391 8.172 ;
			RECT	183.527 8.108 183.559 8.172 ;
			RECT	183.695 8.108 183.727 8.172 ;
			RECT	183.863 8.108 183.895 8.172 ;
			RECT	184.031 8.108 184.063 8.172 ;
			RECT	184.199 8.108 184.231 8.172 ;
			RECT	184.367 8.108 184.399 8.172 ;
			RECT	184.535 8.108 184.567 8.172 ;
			RECT	184.703 8.108 184.735 8.172 ;
			RECT	184.871 8.108 184.903 8.172 ;
			RECT	185.039 8.108 185.071 8.172 ;
			RECT	185.207 8.108 185.239 8.172 ;
			RECT	185.375 8.108 185.407 8.172 ;
			RECT	185.543 8.108 185.575 8.172 ;
			RECT	185.711 8.108 185.743 8.172 ;
			RECT	185.879 8.108 185.911 8.172 ;
			RECT	186.047 8.108 186.079 8.172 ;
			RECT	186.215 8.108 186.247 8.172 ;
			RECT	186.383 8.108 186.415 8.172 ;
			RECT	186.551 8.108 186.583 8.172 ;
			RECT	186.719 8.108 186.751 8.172 ;
			RECT	186.887 8.108 186.919 8.172 ;
			RECT	187.055 8.108 187.087 8.172 ;
			RECT	187.223 8.108 187.255 8.172 ;
			RECT	187.391 8.108 187.423 8.172 ;
			RECT	187.559 8.108 187.591 8.172 ;
			RECT	187.727 8.108 187.759 8.172 ;
			RECT	187.895 8.108 187.927 8.172 ;
			RECT	188.063 8.108 188.095 8.172 ;
			RECT	188.231 8.108 188.263 8.172 ;
			RECT	188.399 8.108 188.431 8.172 ;
			RECT	188.567 8.108 188.599 8.172 ;
			RECT	188.735 8.108 188.767 8.172 ;
			RECT	188.903 8.108 188.935 8.172 ;
			RECT	189.071 8.108 189.103 8.172 ;
			RECT	189.239 8.108 189.271 8.172 ;
			RECT	189.407 8.108 189.439 8.172 ;
			RECT	189.575 8.108 189.607 8.172 ;
			RECT	189.743 8.108 189.775 8.172 ;
			RECT	189.911 8.108 189.943 8.172 ;
			RECT	190.079 8.108 190.111 8.172 ;
			RECT	190.247 8.108 190.279 8.172 ;
			RECT	190.415 8.108 190.447 8.172 ;
			RECT	190.583 8.108 190.615 8.172 ;
			RECT	190.751 8.108 190.783 8.172 ;
			RECT	190.919 8.108 190.951 8.172 ;
			RECT	191.087 8.108 191.119 8.172 ;
			RECT	191.255 8.108 191.287 8.172 ;
			RECT	191.423 8.108 191.455 8.172 ;
			RECT	191.591 8.108 191.623 8.172 ;
			RECT	191.759 8.108 191.791 8.172 ;
			RECT	191.927 8.108 191.959 8.172 ;
			RECT	192.095 8.108 192.127 8.172 ;
			RECT	192.263 8.108 192.295 8.172 ;
			RECT	192.431 8.108 192.463 8.172 ;
			RECT	192.599 8.108 192.631 8.172 ;
			RECT	192.767 8.108 192.799 8.172 ;
			RECT	192.935 8.108 192.967 8.172 ;
			RECT	193.103 8.108 193.135 8.172 ;
			RECT	193.271 8.108 193.303 8.172 ;
			RECT	193.439 8.108 193.471 8.172 ;
			RECT	193.607 8.108 193.639 8.172 ;
			RECT	193.775 8.108 193.807 8.172 ;
			RECT	193.943 8.108 193.975 8.172 ;
			RECT	194.111 8.108 194.143 8.172 ;
			RECT	194.279 8.108 194.311 8.172 ;
			RECT	194.447 8.108 194.479 8.172 ;
			RECT	194.615 8.108 194.647 8.172 ;
			RECT	194.783 8.108 194.815 8.172 ;
			RECT	194.951 8.108 194.983 8.172 ;
			RECT	195.119 8.108 195.151 8.172 ;
			RECT	195.287 8.108 195.319 8.172 ;
			RECT	195.455 8.108 195.487 8.172 ;
			RECT	195.623 8.108 195.655 8.172 ;
			RECT	195.791 8.108 195.823 8.172 ;
			RECT	195.959 8.108 195.991 8.172 ;
			RECT	196.127 8.108 196.159 8.172 ;
			RECT	196.295 8.108 196.327 8.172 ;
			RECT	196.463 8.108 196.495 8.172 ;
			RECT	196.631 8.108 196.663 8.172 ;
			RECT	196.799 8.108 196.831 8.172 ;
			RECT	196.967 8.108 196.999 8.172 ;
			RECT	197.135 8.108 197.167 8.172 ;
			RECT	197.303 8.108 197.335 8.172 ;
			RECT	197.471 8.108 197.503 8.172 ;
			RECT	197.639 8.108 197.671 8.172 ;
			RECT	197.807 8.108 197.839 8.172 ;
			RECT	197.975 8.108 198.007 8.172 ;
			RECT	198.143 8.108 198.175 8.172 ;
			RECT	198.311 8.108 198.343 8.172 ;
			RECT	198.479 8.108 198.511 8.172 ;
			RECT	198.647 8.108 198.679 8.172 ;
			RECT	198.815 8.108 198.847 8.172 ;
			RECT	198.983 8.108 199.015 8.172 ;
			RECT	199.151 8.108 199.183 8.172 ;
			RECT	199.319 8.108 199.351 8.172 ;
			RECT	199.487 8.108 199.519 8.172 ;
			RECT	199.655 8.108 199.687 8.172 ;
			RECT	199.823 8.108 199.855 8.172 ;
			RECT	199.991 8.108 200.023 8.172 ;
			RECT	200.121 8.124 200.153 8.156 ;
			RECT	200.243 8.129 200.275 8.161 ;
			RECT	200.373 8.108 200.405 8.172 ;
			RECT	200.9 8.108 200.932 8.172 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 6.16 201.665 6.28 ;
			LAYER	J3 ;
			RECT	0.755 6.188 0.787 6.252 ;
			RECT	1.645 6.188 1.709 6.252 ;
			RECT	2.323 6.188 2.387 6.252 ;
			RECT	3.438 6.188 3.47 6.252 ;
			RECT	3.585 6.188 3.617 6.252 ;
			RECT	4.195 6.188 4.227 6.252 ;
			RECT	4.72 6.188 4.752 6.252 ;
			RECT	4.944 6.188 5.008 6.252 ;
			RECT	5.267 6.188 5.299 6.252 ;
			RECT	5.797 6.188 5.829 6.252 ;
			RECT	5.927 6.209 5.959 6.241 ;
			RECT	6.049 6.204 6.081 6.236 ;
			RECT	6.179 6.188 6.211 6.252 ;
			RECT	6.347 6.188 6.379 6.252 ;
			RECT	6.515 6.188 6.547 6.252 ;
			RECT	6.683 6.188 6.715 6.252 ;
			RECT	6.851 6.188 6.883 6.252 ;
			RECT	7.019 6.188 7.051 6.252 ;
			RECT	7.187 6.188 7.219 6.252 ;
			RECT	7.355 6.188 7.387 6.252 ;
			RECT	7.523 6.188 7.555 6.252 ;
			RECT	7.691 6.188 7.723 6.252 ;
			RECT	7.859 6.188 7.891 6.252 ;
			RECT	8.027 6.188 8.059 6.252 ;
			RECT	8.195 6.188 8.227 6.252 ;
			RECT	8.363 6.188 8.395 6.252 ;
			RECT	8.531 6.188 8.563 6.252 ;
			RECT	8.699 6.188 8.731 6.252 ;
			RECT	8.867 6.188 8.899 6.252 ;
			RECT	9.035 6.188 9.067 6.252 ;
			RECT	9.203 6.188 9.235 6.252 ;
			RECT	9.371 6.188 9.403 6.252 ;
			RECT	9.539 6.188 9.571 6.252 ;
			RECT	9.707 6.188 9.739 6.252 ;
			RECT	9.875 6.188 9.907 6.252 ;
			RECT	10.043 6.188 10.075 6.252 ;
			RECT	10.211 6.188 10.243 6.252 ;
			RECT	10.379 6.188 10.411 6.252 ;
			RECT	10.547 6.188 10.579 6.252 ;
			RECT	10.715 6.188 10.747 6.252 ;
			RECT	10.883 6.188 10.915 6.252 ;
			RECT	11.051 6.188 11.083 6.252 ;
			RECT	11.219 6.188 11.251 6.252 ;
			RECT	11.387 6.188 11.419 6.252 ;
			RECT	11.555 6.188 11.587 6.252 ;
			RECT	11.723 6.188 11.755 6.252 ;
			RECT	11.891 6.188 11.923 6.252 ;
			RECT	12.059 6.188 12.091 6.252 ;
			RECT	12.227 6.188 12.259 6.252 ;
			RECT	12.395 6.188 12.427 6.252 ;
			RECT	12.563 6.188 12.595 6.252 ;
			RECT	12.731 6.188 12.763 6.252 ;
			RECT	12.899 6.188 12.931 6.252 ;
			RECT	13.067 6.188 13.099 6.252 ;
			RECT	13.235 6.188 13.267 6.252 ;
			RECT	13.403 6.188 13.435 6.252 ;
			RECT	13.571 6.188 13.603 6.252 ;
			RECT	13.739 6.188 13.771 6.252 ;
			RECT	13.907 6.188 13.939 6.252 ;
			RECT	14.075 6.188 14.107 6.252 ;
			RECT	14.243 6.188 14.275 6.252 ;
			RECT	14.411 6.188 14.443 6.252 ;
			RECT	14.579 6.188 14.611 6.252 ;
			RECT	14.747 6.188 14.779 6.252 ;
			RECT	14.915 6.188 14.947 6.252 ;
			RECT	15.083 6.188 15.115 6.252 ;
			RECT	15.251 6.188 15.283 6.252 ;
			RECT	15.419 6.188 15.451 6.252 ;
			RECT	15.587 6.188 15.619 6.252 ;
			RECT	15.755 6.188 15.787 6.252 ;
			RECT	15.923 6.188 15.955 6.252 ;
			RECT	16.091 6.188 16.123 6.252 ;
			RECT	16.259 6.188 16.291 6.252 ;
			RECT	16.427 6.188 16.459 6.252 ;
			RECT	16.595 6.188 16.627 6.252 ;
			RECT	16.763 6.188 16.795 6.252 ;
			RECT	16.931 6.188 16.963 6.252 ;
			RECT	17.099 6.188 17.131 6.252 ;
			RECT	17.267 6.188 17.299 6.252 ;
			RECT	17.435 6.188 17.467 6.252 ;
			RECT	17.603 6.188 17.635 6.252 ;
			RECT	17.771 6.188 17.803 6.252 ;
			RECT	17.939 6.188 17.971 6.252 ;
			RECT	18.107 6.188 18.139 6.252 ;
			RECT	18.275 6.188 18.307 6.252 ;
			RECT	18.443 6.188 18.475 6.252 ;
			RECT	18.611 6.188 18.643 6.252 ;
			RECT	18.779 6.188 18.811 6.252 ;
			RECT	18.947 6.188 18.979 6.252 ;
			RECT	19.115 6.188 19.147 6.252 ;
			RECT	19.283 6.188 19.315 6.252 ;
			RECT	19.451 6.188 19.483 6.252 ;
			RECT	19.619 6.188 19.651 6.252 ;
			RECT	19.787 6.188 19.819 6.252 ;
			RECT	19.955 6.188 19.987 6.252 ;
			RECT	20.123 6.188 20.155 6.252 ;
			RECT	20.291 6.188 20.323 6.252 ;
			RECT	20.459 6.188 20.491 6.252 ;
			RECT	20.627 6.188 20.659 6.252 ;
			RECT	20.795 6.188 20.827 6.252 ;
			RECT	20.963 6.188 20.995 6.252 ;
			RECT	21.131 6.188 21.163 6.252 ;
			RECT	21.299 6.188 21.331 6.252 ;
			RECT	21.467 6.188 21.499 6.252 ;
			RECT	21.635 6.188 21.667 6.252 ;
			RECT	21.803 6.188 21.835 6.252 ;
			RECT	21.971 6.188 22.003 6.252 ;
			RECT	22.139 6.188 22.171 6.252 ;
			RECT	22.307 6.188 22.339 6.252 ;
			RECT	22.475 6.188 22.507 6.252 ;
			RECT	22.643 6.188 22.675 6.252 ;
			RECT	22.811 6.188 22.843 6.252 ;
			RECT	22.979 6.188 23.011 6.252 ;
			RECT	23.147 6.188 23.179 6.252 ;
			RECT	23.315 6.188 23.347 6.252 ;
			RECT	23.483 6.188 23.515 6.252 ;
			RECT	23.651 6.188 23.683 6.252 ;
			RECT	23.819 6.188 23.851 6.252 ;
			RECT	23.987 6.188 24.019 6.252 ;
			RECT	24.155 6.188 24.187 6.252 ;
			RECT	24.323 6.188 24.355 6.252 ;
			RECT	24.491 6.188 24.523 6.252 ;
			RECT	24.659 6.188 24.691 6.252 ;
			RECT	24.827 6.188 24.859 6.252 ;
			RECT	24.995 6.188 25.027 6.252 ;
			RECT	25.163 6.188 25.195 6.252 ;
			RECT	25.331 6.188 25.363 6.252 ;
			RECT	25.499 6.188 25.531 6.252 ;
			RECT	25.667 6.188 25.699 6.252 ;
			RECT	25.835 6.188 25.867 6.252 ;
			RECT	26.003 6.188 26.035 6.252 ;
			RECT	26.171 6.188 26.203 6.252 ;
			RECT	26.339 6.188 26.371 6.252 ;
			RECT	26.507 6.188 26.539 6.252 ;
			RECT	26.675 6.188 26.707 6.252 ;
			RECT	26.843 6.188 26.875 6.252 ;
			RECT	27.011 6.188 27.043 6.252 ;
			RECT	27.179 6.188 27.211 6.252 ;
			RECT	27.347 6.188 27.379 6.252 ;
			RECT	27.515 6.188 27.547 6.252 ;
			RECT	27.683 6.188 27.715 6.252 ;
			RECT	27.851 6.188 27.883 6.252 ;
			RECT	28.019 6.188 28.051 6.252 ;
			RECT	28.187 6.188 28.219 6.252 ;
			RECT	28.355 6.188 28.387 6.252 ;
			RECT	28.523 6.188 28.555 6.252 ;
			RECT	28.691 6.188 28.723 6.252 ;
			RECT	28.859 6.188 28.891 6.252 ;
			RECT	29.027 6.188 29.059 6.252 ;
			RECT	29.195 6.188 29.227 6.252 ;
			RECT	29.363 6.188 29.395 6.252 ;
			RECT	29.531 6.188 29.563 6.252 ;
			RECT	29.699 6.188 29.731 6.252 ;
			RECT	29.867 6.188 29.899 6.252 ;
			RECT	30.035 6.188 30.067 6.252 ;
			RECT	30.203 6.188 30.235 6.252 ;
			RECT	30.371 6.188 30.403 6.252 ;
			RECT	30.539 6.188 30.571 6.252 ;
			RECT	30.707 6.188 30.739 6.252 ;
			RECT	30.875 6.188 30.907 6.252 ;
			RECT	31.043 6.188 31.075 6.252 ;
			RECT	31.211 6.188 31.243 6.252 ;
			RECT	31.379 6.188 31.411 6.252 ;
			RECT	31.547 6.188 31.579 6.252 ;
			RECT	31.715 6.188 31.747 6.252 ;
			RECT	31.883 6.188 31.915 6.252 ;
			RECT	32.051 6.188 32.083 6.252 ;
			RECT	32.219 6.188 32.251 6.252 ;
			RECT	32.387 6.188 32.419 6.252 ;
			RECT	32.555 6.188 32.587 6.252 ;
			RECT	32.723 6.188 32.755 6.252 ;
			RECT	32.891 6.188 32.923 6.252 ;
			RECT	33.059 6.188 33.091 6.252 ;
			RECT	33.227 6.188 33.259 6.252 ;
			RECT	33.395 6.188 33.427 6.252 ;
			RECT	33.563 6.188 33.595 6.252 ;
			RECT	33.731 6.188 33.763 6.252 ;
			RECT	33.899 6.188 33.931 6.252 ;
			RECT	34.067 6.188 34.099 6.252 ;
			RECT	34.235 6.188 34.267 6.252 ;
			RECT	34.403 6.188 34.435 6.252 ;
			RECT	34.571 6.188 34.603 6.252 ;
			RECT	34.739 6.188 34.771 6.252 ;
			RECT	34.907 6.188 34.939 6.252 ;
			RECT	35.075 6.188 35.107 6.252 ;
			RECT	35.243 6.188 35.275 6.252 ;
			RECT	35.411 6.188 35.443 6.252 ;
			RECT	35.579 6.188 35.611 6.252 ;
			RECT	35.747 6.188 35.779 6.252 ;
			RECT	35.915 6.188 35.947 6.252 ;
			RECT	36.083 6.188 36.115 6.252 ;
			RECT	36.251 6.188 36.283 6.252 ;
			RECT	36.419 6.188 36.451 6.252 ;
			RECT	36.587 6.188 36.619 6.252 ;
			RECT	36.755 6.188 36.787 6.252 ;
			RECT	36.923 6.188 36.955 6.252 ;
			RECT	37.091 6.188 37.123 6.252 ;
			RECT	37.259 6.188 37.291 6.252 ;
			RECT	37.427 6.188 37.459 6.252 ;
			RECT	37.595 6.188 37.627 6.252 ;
			RECT	37.763 6.188 37.795 6.252 ;
			RECT	37.931 6.188 37.963 6.252 ;
			RECT	38.099 6.188 38.131 6.252 ;
			RECT	38.267 6.188 38.299 6.252 ;
			RECT	38.435 6.188 38.467 6.252 ;
			RECT	38.603 6.188 38.635 6.252 ;
			RECT	38.771 6.188 38.803 6.252 ;
			RECT	38.939 6.188 38.971 6.252 ;
			RECT	39.107 6.188 39.139 6.252 ;
			RECT	39.275 6.188 39.307 6.252 ;
			RECT	39.443 6.188 39.475 6.252 ;
			RECT	39.611 6.188 39.643 6.252 ;
			RECT	39.779 6.188 39.811 6.252 ;
			RECT	39.947 6.188 39.979 6.252 ;
			RECT	40.115 6.188 40.147 6.252 ;
			RECT	40.283 6.188 40.315 6.252 ;
			RECT	40.451 6.188 40.483 6.252 ;
			RECT	40.619 6.188 40.651 6.252 ;
			RECT	40.787 6.188 40.819 6.252 ;
			RECT	40.955 6.188 40.987 6.252 ;
			RECT	41.123 6.188 41.155 6.252 ;
			RECT	41.291 6.188 41.323 6.252 ;
			RECT	41.459 6.188 41.491 6.252 ;
			RECT	41.627 6.188 41.659 6.252 ;
			RECT	41.795 6.188 41.827 6.252 ;
			RECT	41.963 6.188 41.995 6.252 ;
			RECT	42.131 6.188 42.163 6.252 ;
			RECT	42.299 6.188 42.331 6.252 ;
			RECT	42.467 6.188 42.499 6.252 ;
			RECT	42.635 6.188 42.667 6.252 ;
			RECT	42.803 6.188 42.835 6.252 ;
			RECT	42.971 6.188 43.003 6.252 ;
			RECT	43.139 6.188 43.171 6.252 ;
			RECT	43.307 6.188 43.339 6.252 ;
			RECT	43.475 6.188 43.507 6.252 ;
			RECT	43.643 6.188 43.675 6.252 ;
			RECT	43.811 6.188 43.843 6.252 ;
			RECT	43.979 6.188 44.011 6.252 ;
			RECT	44.147 6.188 44.179 6.252 ;
			RECT	44.315 6.188 44.347 6.252 ;
			RECT	44.483 6.188 44.515 6.252 ;
			RECT	44.651 6.188 44.683 6.252 ;
			RECT	44.819 6.188 44.851 6.252 ;
			RECT	44.987 6.188 45.019 6.252 ;
			RECT	45.155 6.188 45.187 6.252 ;
			RECT	45.323 6.188 45.355 6.252 ;
			RECT	45.491 6.188 45.523 6.252 ;
			RECT	45.659 6.188 45.691 6.252 ;
			RECT	45.827 6.188 45.859 6.252 ;
			RECT	45.995 6.188 46.027 6.252 ;
			RECT	46.163 6.188 46.195 6.252 ;
			RECT	46.331 6.188 46.363 6.252 ;
			RECT	46.499 6.188 46.531 6.252 ;
			RECT	46.667 6.188 46.699 6.252 ;
			RECT	46.835 6.188 46.867 6.252 ;
			RECT	47.003 6.188 47.035 6.252 ;
			RECT	47.171 6.188 47.203 6.252 ;
			RECT	47.339 6.188 47.371 6.252 ;
			RECT	47.507 6.188 47.539 6.252 ;
			RECT	47.675 6.188 47.707 6.252 ;
			RECT	47.843 6.188 47.875 6.252 ;
			RECT	48.011 6.188 48.043 6.252 ;
			RECT	48.179 6.188 48.211 6.252 ;
			RECT	48.347 6.188 48.379 6.252 ;
			RECT	48.515 6.188 48.547 6.252 ;
			RECT	48.683 6.188 48.715 6.252 ;
			RECT	48.851 6.188 48.883 6.252 ;
			RECT	49.019 6.188 49.051 6.252 ;
			RECT	49.187 6.188 49.219 6.252 ;
			RECT	49.318 6.204 49.35 6.236 ;
			RECT	49.439 6.204 49.471 6.236 ;
			RECT	49.569 6.188 49.601 6.252 ;
			RECT	51.881 6.188 51.913 6.252 ;
			RECT	53.132 6.188 53.196 6.252 ;
			RECT	53.812 6.188 53.844 6.252 ;
			RECT	54.251 6.188 54.283 6.252 ;
			RECT	55.562 6.188 55.626 6.252 ;
			RECT	58.603 6.188 58.635 6.252 ;
			RECT	58.733 6.204 58.765 6.236 ;
			RECT	58.854 6.204 58.886 6.236 ;
			RECT	58.985 6.188 59.017 6.252 ;
			RECT	59.153 6.188 59.185 6.252 ;
			RECT	59.321 6.188 59.353 6.252 ;
			RECT	59.489 6.188 59.521 6.252 ;
			RECT	59.657 6.188 59.689 6.252 ;
			RECT	59.825 6.188 59.857 6.252 ;
			RECT	59.993 6.188 60.025 6.252 ;
			RECT	60.161 6.188 60.193 6.252 ;
			RECT	60.329 6.188 60.361 6.252 ;
			RECT	60.497 6.188 60.529 6.252 ;
			RECT	60.665 6.188 60.697 6.252 ;
			RECT	60.833 6.188 60.865 6.252 ;
			RECT	61.001 6.188 61.033 6.252 ;
			RECT	61.169 6.188 61.201 6.252 ;
			RECT	61.337 6.188 61.369 6.252 ;
			RECT	61.505 6.188 61.537 6.252 ;
			RECT	61.673 6.188 61.705 6.252 ;
			RECT	61.841 6.188 61.873 6.252 ;
			RECT	62.009 6.188 62.041 6.252 ;
			RECT	62.177 6.188 62.209 6.252 ;
			RECT	62.345 6.188 62.377 6.252 ;
			RECT	62.513 6.188 62.545 6.252 ;
			RECT	62.681 6.188 62.713 6.252 ;
			RECT	62.849 6.188 62.881 6.252 ;
			RECT	63.017 6.188 63.049 6.252 ;
			RECT	63.185 6.188 63.217 6.252 ;
			RECT	63.353 6.188 63.385 6.252 ;
			RECT	63.521 6.188 63.553 6.252 ;
			RECT	63.689 6.188 63.721 6.252 ;
			RECT	63.857 6.188 63.889 6.252 ;
			RECT	64.025 6.188 64.057 6.252 ;
			RECT	64.193 6.188 64.225 6.252 ;
			RECT	64.361 6.188 64.393 6.252 ;
			RECT	64.529 6.188 64.561 6.252 ;
			RECT	64.697 6.188 64.729 6.252 ;
			RECT	64.865 6.188 64.897 6.252 ;
			RECT	65.033 6.188 65.065 6.252 ;
			RECT	65.201 6.188 65.233 6.252 ;
			RECT	65.369 6.188 65.401 6.252 ;
			RECT	65.537 6.188 65.569 6.252 ;
			RECT	65.705 6.188 65.737 6.252 ;
			RECT	65.873 6.188 65.905 6.252 ;
			RECT	66.041 6.188 66.073 6.252 ;
			RECT	66.209 6.188 66.241 6.252 ;
			RECT	66.377 6.188 66.409 6.252 ;
			RECT	66.545 6.188 66.577 6.252 ;
			RECT	66.713 6.188 66.745 6.252 ;
			RECT	66.881 6.188 66.913 6.252 ;
			RECT	67.049 6.188 67.081 6.252 ;
			RECT	67.217 6.188 67.249 6.252 ;
			RECT	67.385 6.188 67.417 6.252 ;
			RECT	67.553 6.188 67.585 6.252 ;
			RECT	67.721 6.188 67.753 6.252 ;
			RECT	67.889 6.188 67.921 6.252 ;
			RECT	68.057 6.188 68.089 6.252 ;
			RECT	68.225 6.188 68.257 6.252 ;
			RECT	68.393 6.188 68.425 6.252 ;
			RECT	68.561 6.188 68.593 6.252 ;
			RECT	68.729 6.188 68.761 6.252 ;
			RECT	68.897 6.188 68.929 6.252 ;
			RECT	69.065 6.188 69.097 6.252 ;
			RECT	69.233 6.188 69.265 6.252 ;
			RECT	69.401 6.188 69.433 6.252 ;
			RECT	69.569 6.188 69.601 6.252 ;
			RECT	69.737 6.188 69.769 6.252 ;
			RECT	69.905 6.188 69.937 6.252 ;
			RECT	70.073 6.188 70.105 6.252 ;
			RECT	70.241 6.188 70.273 6.252 ;
			RECT	70.409 6.188 70.441 6.252 ;
			RECT	70.577 6.188 70.609 6.252 ;
			RECT	70.745 6.188 70.777 6.252 ;
			RECT	70.913 6.188 70.945 6.252 ;
			RECT	71.081 6.188 71.113 6.252 ;
			RECT	71.249 6.188 71.281 6.252 ;
			RECT	71.417 6.188 71.449 6.252 ;
			RECT	71.585 6.188 71.617 6.252 ;
			RECT	71.753 6.188 71.785 6.252 ;
			RECT	71.921 6.188 71.953 6.252 ;
			RECT	72.089 6.188 72.121 6.252 ;
			RECT	72.257 6.188 72.289 6.252 ;
			RECT	72.425 6.188 72.457 6.252 ;
			RECT	72.593 6.188 72.625 6.252 ;
			RECT	72.761 6.188 72.793 6.252 ;
			RECT	72.929 6.188 72.961 6.252 ;
			RECT	73.097 6.188 73.129 6.252 ;
			RECT	73.265 6.188 73.297 6.252 ;
			RECT	73.433 6.188 73.465 6.252 ;
			RECT	73.601 6.188 73.633 6.252 ;
			RECT	73.769 6.188 73.801 6.252 ;
			RECT	73.937 6.188 73.969 6.252 ;
			RECT	74.105 6.188 74.137 6.252 ;
			RECT	74.273 6.188 74.305 6.252 ;
			RECT	74.441 6.188 74.473 6.252 ;
			RECT	74.609 6.188 74.641 6.252 ;
			RECT	74.777 6.188 74.809 6.252 ;
			RECT	74.945 6.188 74.977 6.252 ;
			RECT	75.113 6.188 75.145 6.252 ;
			RECT	75.281 6.188 75.313 6.252 ;
			RECT	75.449 6.188 75.481 6.252 ;
			RECT	75.617 6.188 75.649 6.252 ;
			RECT	75.785 6.188 75.817 6.252 ;
			RECT	75.953 6.188 75.985 6.252 ;
			RECT	76.121 6.188 76.153 6.252 ;
			RECT	76.289 6.188 76.321 6.252 ;
			RECT	76.457 6.188 76.489 6.252 ;
			RECT	76.625 6.188 76.657 6.252 ;
			RECT	76.793 6.188 76.825 6.252 ;
			RECT	76.961 6.188 76.993 6.252 ;
			RECT	77.129 6.188 77.161 6.252 ;
			RECT	77.297 6.188 77.329 6.252 ;
			RECT	77.465 6.188 77.497 6.252 ;
			RECT	77.633 6.188 77.665 6.252 ;
			RECT	77.801 6.188 77.833 6.252 ;
			RECT	77.969 6.188 78.001 6.252 ;
			RECT	78.137 6.188 78.169 6.252 ;
			RECT	78.305 6.188 78.337 6.252 ;
			RECT	78.473 6.188 78.505 6.252 ;
			RECT	78.641 6.188 78.673 6.252 ;
			RECT	78.809 6.188 78.841 6.252 ;
			RECT	78.977 6.188 79.009 6.252 ;
			RECT	79.145 6.188 79.177 6.252 ;
			RECT	79.313 6.188 79.345 6.252 ;
			RECT	79.481 6.188 79.513 6.252 ;
			RECT	79.649 6.188 79.681 6.252 ;
			RECT	79.817 6.188 79.849 6.252 ;
			RECT	79.985 6.188 80.017 6.252 ;
			RECT	80.153 6.188 80.185 6.252 ;
			RECT	80.321 6.188 80.353 6.252 ;
			RECT	80.489 6.188 80.521 6.252 ;
			RECT	80.657 6.188 80.689 6.252 ;
			RECT	80.825 6.188 80.857 6.252 ;
			RECT	80.993 6.188 81.025 6.252 ;
			RECT	81.161 6.188 81.193 6.252 ;
			RECT	81.329 6.188 81.361 6.252 ;
			RECT	81.497 6.188 81.529 6.252 ;
			RECT	81.665 6.188 81.697 6.252 ;
			RECT	81.833 6.188 81.865 6.252 ;
			RECT	82.001 6.188 82.033 6.252 ;
			RECT	82.169 6.188 82.201 6.252 ;
			RECT	82.337 6.188 82.369 6.252 ;
			RECT	82.505 6.188 82.537 6.252 ;
			RECT	82.673 6.188 82.705 6.252 ;
			RECT	82.841 6.188 82.873 6.252 ;
			RECT	83.009 6.188 83.041 6.252 ;
			RECT	83.177 6.188 83.209 6.252 ;
			RECT	83.345 6.188 83.377 6.252 ;
			RECT	83.513 6.188 83.545 6.252 ;
			RECT	83.681 6.188 83.713 6.252 ;
			RECT	83.849 6.188 83.881 6.252 ;
			RECT	84.017 6.188 84.049 6.252 ;
			RECT	84.185 6.188 84.217 6.252 ;
			RECT	84.353 6.188 84.385 6.252 ;
			RECT	84.521 6.188 84.553 6.252 ;
			RECT	84.689 6.188 84.721 6.252 ;
			RECT	84.857 6.188 84.889 6.252 ;
			RECT	85.025 6.188 85.057 6.252 ;
			RECT	85.193 6.188 85.225 6.252 ;
			RECT	85.361 6.188 85.393 6.252 ;
			RECT	85.529 6.188 85.561 6.252 ;
			RECT	85.697 6.188 85.729 6.252 ;
			RECT	85.865 6.188 85.897 6.252 ;
			RECT	86.033 6.188 86.065 6.252 ;
			RECT	86.201 6.188 86.233 6.252 ;
			RECT	86.369 6.188 86.401 6.252 ;
			RECT	86.537 6.188 86.569 6.252 ;
			RECT	86.705 6.188 86.737 6.252 ;
			RECT	86.873 6.188 86.905 6.252 ;
			RECT	87.041 6.188 87.073 6.252 ;
			RECT	87.209 6.188 87.241 6.252 ;
			RECT	87.377 6.188 87.409 6.252 ;
			RECT	87.545 6.188 87.577 6.252 ;
			RECT	87.713 6.188 87.745 6.252 ;
			RECT	87.881 6.188 87.913 6.252 ;
			RECT	88.049 6.188 88.081 6.252 ;
			RECT	88.217 6.188 88.249 6.252 ;
			RECT	88.385 6.188 88.417 6.252 ;
			RECT	88.553 6.188 88.585 6.252 ;
			RECT	88.721 6.188 88.753 6.252 ;
			RECT	88.889 6.188 88.921 6.252 ;
			RECT	89.057 6.188 89.089 6.252 ;
			RECT	89.225 6.188 89.257 6.252 ;
			RECT	89.393 6.188 89.425 6.252 ;
			RECT	89.561 6.188 89.593 6.252 ;
			RECT	89.729 6.188 89.761 6.252 ;
			RECT	89.897 6.188 89.929 6.252 ;
			RECT	90.065 6.188 90.097 6.252 ;
			RECT	90.233 6.188 90.265 6.252 ;
			RECT	90.401 6.188 90.433 6.252 ;
			RECT	90.569 6.188 90.601 6.252 ;
			RECT	90.737 6.188 90.769 6.252 ;
			RECT	90.905 6.188 90.937 6.252 ;
			RECT	91.073 6.188 91.105 6.252 ;
			RECT	91.241 6.188 91.273 6.252 ;
			RECT	91.409 6.188 91.441 6.252 ;
			RECT	91.577 6.188 91.609 6.252 ;
			RECT	91.745 6.188 91.777 6.252 ;
			RECT	91.913 6.188 91.945 6.252 ;
			RECT	92.081 6.188 92.113 6.252 ;
			RECT	92.249 6.188 92.281 6.252 ;
			RECT	92.417 6.188 92.449 6.252 ;
			RECT	92.585 6.188 92.617 6.252 ;
			RECT	92.753 6.188 92.785 6.252 ;
			RECT	92.921 6.188 92.953 6.252 ;
			RECT	93.089 6.188 93.121 6.252 ;
			RECT	93.257 6.188 93.289 6.252 ;
			RECT	93.425 6.188 93.457 6.252 ;
			RECT	93.593 6.188 93.625 6.252 ;
			RECT	93.761 6.188 93.793 6.252 ;
			RECT	93.929 6.188 93.961 6.252 ;
			RECT	94.097 6.188 94.129 6.252 ;
			RECT	94.265 6.188 94.297 6.252 ;
			RECT	94.433 6.188 94.465 6.252 ;
			RECT	94.601 6.188 94.633 6.252 ;
			RECT	94.769 6.188 94.801 6.252 ;
			RECT	94.937 6.188 94.969 6.252 ;
			RECT	95.105 6.188 95.137 6.252 ;
			RECT	95.273 6.188 95.305 6.252 ;
			RECT	95.441 6.188 95.473 6.252 ;
			RECT	95.609 6.188 95.641 6.252 ;
			RECT	95.777 6.188 95.809 6.252 ;
			RECT	95.945 6.188 95.977 6.252 ;
			RECT	96.113 6.188 96.145 6.252 ;
			RECT	96.281 6.188 96.313 6.252 ;
			RECT	96.449 6.188 96.481 6.252 ;
			RECT	96.617 6.188 96.649 6.252 ;
			RECT	96.785 6.188 96.817 6.252 ;
			RECT	96.953 6.188 96.985 6.252 ;
			RECT	97.121 6.188 97.153 6.252 ;
			RECT	97.289 6.188 97.321 6.252 ;
			RECT	97.457 6.188 97.489 6.252 ;
			RECT	97.625 6.188 97.657 6.252 ;
			RECT	97.793 6.188 97.825 6.252 ;
			RECT	97.961 6.188 97.993 6.252 ;
			RECT	98.129 6.188 98.161 6.252 ;
			RECT	98.297 6.188 98.329 6.252 ;
			RECT	98.465 6.188 98.497 6.252 ;
			RECT	98.633 6.188 98.665 6.252 ;
			RECT	98.801 6.188 98.833 6.252 ;
			RECT	98.969 6.188 99.001 6.252 ;
			RECT	99.137 6.188 99.169 6.252 ;
			RECT	99.305 6.188 99.337 6.252 ;
			RECT	99.473 6.188 99.505 6.252 ;
			RECT	99.641 6.188 99.673 6.252 ;
			RECT	99.809 6.188 99.841 6.252 ;
			RECT	99.977 6.188 100.009 6.252 ;
			RECT	100.145 6.188 100.177 6.252 ;
			RECT	100.313 6.188 100.345 6.252 ;
			RECT	100.481 6.188 100.513 6.252 ;
			RECT	100.649 6.188 100.681 6.252 ;
			RECT	100.817 6.188 100.849 6.252 ;
			RECT	100.985 6.188 101.017 6.252 ;
			RECT	101.153 6.188 101.185 6.252 ;
			RECT	101.321 6.188 101.353 6.252 ;
			RECT	101.489 6.188 101.521 6.252 ;
			RECT	101.657 6.188 101.689 6.252 ;
			RECT	101.825 6.188 101.857 6.252 ;
			RECT	101.993 6.188 102.025 6.252 ;
			RECT	102.123 6.204 102.155 6.236 ;
			RECT	102.245 6.209 102.277 6.241 ;
			RECT	102.375 6.188 102.407 6.252 ;
			RECT	103.795 6.188 103.827 6.252 ;
			RECT	103.925 6.209 103.957 6.241 ;
			RECT	104.047 6.204 104.079 6.236 ;
			RECT	104.177 6.188 104.209 6.252 ;
			RECT	104.345 6.188 104.377 6.252 ;
			RECT	104.513 6.188 104.545 6.252 ;
			RECT	104.681 6.188 104.713 6.252 ;
			RECT	104.849 6.188 104.881 6.252 ;
			RECT	105.017 6.188 105.049 6.252 ;
			RECT	105.185 6.188 105.217 6.252 ;
			RECT	105.353 6.188 105.385 6.252 ;
			RECT	105.521 6.188 105.553 6.252 ;
			RECT	105.689 6.188 105.721 6.252 ;
			RECT	105.857 6.188 105.889 6.252 ;
			RECT	106.025 6.188 106.057 6.252 ;
			RECT	106.193 6.188 106.225 6.252 ;
			RECT	106.361 6.188 106.393 6.252 ;
			RECT	106.529 6.188 106.561 6.252 ;
			RECT	106.697 6.188 106.729 6.252 ;
			RECT	106.865 6.188 106.897 6.252 ;
			RECT	107.033 6.188 107.065 6.252 ;
			RECT	107.201 6.188 107.233 6.252 ;
			RECT	107.369 6.188 107.401 6.252 ;
			RECT	107.537 6.188 107.569 6.252 ;
			RECT	107.705 6.188 107.737 6.252 ;
			RECT	107.873 6.188 107.905 6.252 ;
			RECT	108.041 6.188 108.073 6.252 ;
			RECT	108.209 6.188 108.241 6.252 ;
			RECT	108.377 6.188 108.409 6.252 ;
			RECT	108.545 6.188 108.577 6.252 ;
			RECT	108.713 6.188 108.745 6.252 ;
			RECT	108.881 6.188 108.913 6.252 ;
			RECT	109.049 6.188 109.081 6.252 ;
			RECT	109.217 6.188 109.249 6.252 ;
			RECT	109.385 6.188 109.417 6.252 ;
			RECT	109.553 6.188 109.585 6.252 ;
			RECT	109.721 6.188 109.753 6.252 ;
			RECT	109.889 6.188 109.921 6.252 ;
			RECT	110.057 6.188 110.089 6.252 ;
			RECT	110.225 6.188 110.257 6.252 ;
			RECT	110.393 6.188 110.425 6.252 ;
			RECT	110.561 6.188 110.593 6.252 ;
			RECT	110.729 6.188 110.761 6.252 ;
			RECT	110.897 6.188 110.929 6.252 ;
			RECT	111.065 6.188 111.097 6.252 ;
			RECT	111.233 6.188 111.265 6.252 ;
			RECT	111.401 6.188 111.433 6.252 ;
			RECT	111.569 6.188 111.601 6.252 ;
			RECT	111.737 6.188 111.769 6.252 ;
			RECT	111.905 6.188 111.937 6.252 ;
			RECT	112.073 6.188 112.105 6.252 ;
			RECT	112.241 6.188 112.273 6.252 ;
			RECT	112.409 6.188 112.441 6.252 ;
			RECT	112.577 6.188 112.609 6.252 ;
			RECT	112.745 6.188 112.777 6.252 ;
			RECT	112.913 6.188 112.945 6.252 ;
			RECT	113.081 6.188 113.113 6.252 ;
			RECT	113.249 6.188 113.281 6.252 ;
			RECT	113.417 6.188 113.449 6.252 ;
			RECT	113.585 6.188 113.617 6.252 ;
			RECT	113.753 6.188 113.785 6.252 ;
			RECT	113.921 6.188 113.953 6.252 ;
			RECT	114.089 6.188 114.121 6.252 ;
			RECT	114.257 6.188 114.289 6.252 ;
			RECT	114.425 6.188 114.457 6.252 ;
			RECT	114.593 6.188 114.625 6.252 ;
			RECT	114.761 6.188 114.793 6.252 ;
			RECT	114.929 6.188 114.961 6.252 ;
			RECT	115.097 6.188 115.129 6.252 ;
			RECT	115.265 6.188 115.297 6.252 ;
			RECT	115.433 6.188 115.465 6.252 ;
			RECT	115.601 6.188 115.633 6.252 ;
			RECT	115.769 6.188 115.801 6.252 ;
			RECT	115.937 6.188 115.969 6.252 ;
			RECT	116.105 6.188 116.137 6.252 ;
			RECT	116.273 6.188 116.305 6.252 ;
			RECT	116.441 6.188 116.473 6.252 ;
			RECT	116.609 6.188 116.641 6.252 ;
			RECT	116.777 6.188 116.809 6.252 ;
			RECT	116.945 6.188 116.977 6.252 ;
			RECT	117.113 6.188 117.145 6.252 ;
			RECT	117.281 6.188 117.313 6.252 ;
			RECT	117.449 6.188 117.481 6.252 ;
			RECT	117.617 6.188 117.649 6.252 ;
			RECT	117.785 6.188 117.817 6.252 ;
			RECT	117.953 6.188 117.985 6.252 ;
			RECT	118.121 6.188 118.153 6.252 ;
			RECT	118.289 6.188 118.321 6.252 ;
			RECT	118.457 6.188 118.489 6.252 ;
			RECT	118.625 6.188 118.657 6.252 ;
			RECT	118.793 6.188 118.825 6.252 ;
			RECT	118.961 6.188 118.993 6.252 ;
			RECT	119.129 6.188 119.161 6.252 ;
			RECT	119.297 6.188 119.329 6.252 ;
			RECT	119.465 6.188 119.497 6.252 ;
			RECT	119.633 6.188 119.665 6.252 ;
			RECT	119.801 6.188 119.833 6.252 ;
			RECT	119.969 6.188 120.001 6.252 ;
			RECT	120.137 6.188 120.169 6.252 ;
			RECT	120.305 6.188 120.337 6.252 ;
			RECT	120.473 6.188 120.505 6.252 ;
			RECT	120.641 6.188 120.673 6.252 ;
			RECT	120.809 6.188 120.841 6.252 ;
			RECT	120.977 6.188 121.009 6.252 ;
			RECT	121.145 6.188 121.177 6.252 ;
			RECT	121.313 6.188 121.345 6.252 ;
			RECT	121.481 6.188 121.513 6.252 ;
			RECT	121.649 6.188 121.681 6.252 ;
			RECT	121.817 6.188 121.849 6.252 ;
			RECT	121.985 6.188 122.017 6.252 ;
			RECT	122.153 6.188 122.185 6.252 ;
			RECT	122.321 6.188 122.353 6.252 ;
			RECT	122.489 6.188 122.521 6.252 ;
			RECT	122.657 6.188 122.689 6.252 ;
			RECT	122.825 6.188 122.857 6.252 ;
			RECT	122.993 6.188 123.025 6.252 ;
			RECT	123.161 6.188 123.193 6.252 ;
			RECT	123.329 6.188 123.361 6.252 ;
			RECT	123.497 6.188 123.529 6.252 ;
			RECT	123.665 6.188 123.697 6.252 ;
			RECT	123.833 6.188 123.865 6.252 ;
			RECT	124.001 6.188 124.033 6.252 ;
			RECT	124.169 6.188 124.201 6.252 ;
			RECT	124.337 6.188 124.369 6.252 ;
			RECT	124.505 6.188 124.537 6.252 ;
			RECT	124.673 6.188 124.705 6.252 ;
			RECT	124.841 6.188 124.873 6.252 ;
			RECT	125.009 6.188 125.041 6.252 ;
			RECT	125.177 6.188 125.209 6.252 ;
			RECT	125.345 6.188 125.377 6.252 ;
			RECT	125.513 6.188 125.545 6.252 ;
			RECT	125.681 6.188 125.713 6.252 ;
			RECT	125.849 6.188 125.881 6.252 ;
			RECT	126.017 6.188 126.049 6.252 ;
			RECT	126.185 6.188 126.217 6.252 ;
			RECT	126.353 6.188 126.385 6.252 ;
			RECT	126.521 6.188 126.553 6.252 ;
			RECT	126.689 6.188 126.721 6.252 ;
			RECT	126.857 6.188 126.889 6.252 ;
			RECT	127.025 6.188 127.057 6.252 ;
			RECT	127.193 6.188 127.225 6.252 ;
			RECT	127.361 6.188 127.393 6.252 ;
			RECT	127.529 6.188 127.561 6.252 ;
			RECT	127.697 6.188 127.729 6.252 ;
			RECT	127.865 6.188 127.897 6.252 ;
			RECT	128.033 6.188 128.065 6.252 ;
			RECT	128.201 6.188 128.233 6.252 ;
			RECT	128.369 6.188 128.401 6.252 ;
			RECT	128.537 6.188 128.569 6.252 ;
			RECT	128.705 6.188 128.737 6.252 ;
			RECT	128.873 6.188 128.905 6.252 ;
			RECT	129.041 6.188 129.073 6.252 ;
			RECT	129.209 6.188 129.241 6.252 ;
			RECT	129.377 6.188 129.409 6.252 ;
			RECT	129.545 6.188 129.577 6.252 ;
			RECT	129.713 6.188 129.745 6.252 ;
			RECT	129.881 6.188 129.913 6.252 ;
			RECT	130.049 6.188 130.081 6.252 ;
			RECT	130.217 6.188 130.249 6.252 ;
			RECT	130.385 6.188 130.417 6.252 ;
			RECT	130.553 6.188 130.585 6.252 ;
			RECT	130.721 6.188 130.753 6.252 ;
			RECT	130.889 6.188 130.921 6.252 ;
			RECT	131.057 6.188 131.089 6.252 ;
			RECT	131.225 6.188 131.257 6.252 ;
			RECT	131.393 6.188 131.425 6.252 ;
			RECT	131.561 6.188 131.593 6.252 ;
			RECT	131.729 6.188 131.761 6.252 ;
			RECT	131.897 6.188 131.929 6.252 ;
			RECT	132.065 6.188 132.097 6.252 ;
			RECT	132.233 6.188 132.265 6.252 ;
			RECT	132.401 6.188 132.433 6.252 ;
			RECT	132.569 6.188 132.601 6.252 ;
			RECT	132.737 6.188 132.769 6.252 ;
			RECT	132.905 6.188 132.937 6.252 ;
			RECT	133.073 6.188 133.105 6.252 ;
			RECT	133.241 6.188 133.273 6.252 ;
			RECT	133.409 6.188 133.441 6.252 ;
			RECT	133.577 6.188 133.609 6.252 ;
			RECT	133.745 6.188 133.777 6.252 ;
			RECT	133.913 6.188 133.945 6.252 ;
			RECT	134.081 6.188 134.113 6.252 ;
			RECT	134.249 6.188 134.281 6.252 ;
			RECT	134.417 6.188 134.449 6.252 ;
			RECT	134.585 6.188 134.617 6.252 ;
			RECT	134.753 6.188 134.785 6.252 ;
			RECT	134.921 6.188 134.953 6.252 ;
			RECT	135.089 6.188 135.121 6.252 ;
			RECT	135.257 6.188 135.289 6.252 ;
			RECT	135.425 6.188 135.457 6.252 ;
			RECT	135.593 6.188 135.625 6.252 ;
			RECT	135.761 6.188 135.793 6.252 ;
			RECT	135.929 6.188 135.961 6.252 ;
			RECT	136.097 6.188 136.129 6.252 ;
			RECT	136.265 6.188 136.297 6.252 ;
			RECT	136.433 6.188 136.465 6.252 ;
			RECT	136.601 6.188 136.633 6.252 ;
			RECT	136.769 6.188 136.801 6.252 ;
			RECT	136.937 6.188 136.969 6.252 ;
			RECT	137.105 6.188 137.137 6.252 ;
			RECT	137.273 6.188 137.305 6.252 ;
			RECT	137.441 6.188 137.473 6.252 ;
			RECT	137.609 6.188 137.641 6.252 ;
			RECT	137.777 6.188 137.809 6.252 ;
			RECT	137.945 6.188 137.977 6.252 ;
			RECT	138.113 6.188 138.145 6.252 ;
			RECT	138.281 6.188 138.313 6.252 ;
			RECT	138.449 6.188 138.481 6.252 ;
			RECT	138.617 6.188 138.649 6.252 ;
			RECT	138.785 6.188 138.817 6.252 ;
			RECT	138.953 6.188 138.985 6.252 ;
			RECT	139.121 6.188 139.153 6.252 ;
			RECT	139.289 6.188 139.321 6.252 ;
			RECT	139.457 6.188 139.489 6.252 ;
			RECT	139.625 6.188 139.657 6.252 ;
			RECT	139.793 6.188 139.825 6.252 ;
			RECT	139.961 6.188 139.993 6.252 ;
			RECT	140.129 6.188 140.161 6.252 ;
			RECT	140.297 6.188 140.329 6.252 ;
			RECT	140.465 6.188 140.497 6.252 ;
			RECT	140.633 6.188 140.665 6.252 ;
			RECT	140.801 6.188 140.833 6.252 ;
			RECT	140.969 6.188 141.001 6.252 ;
			RECT	141.137 6.188 141.169 6.252 ;
			RECT	141.305 6.188 141.337 6.252 ;
			RECT	141.473 6.188 141.505 6.252 ;
			RECT	141.641 6.188 141.673 6.252 ;
			RECT	141.809 6.188 141.841 6.252 ;
			RECT	141.977 6.188 142.009 6.252 ;
			RECT	142.145 6.188 142.177 6.252 ;
			RECT	142.313 6.188 142.345 6.252 ;
			RECT	142.481 6.188 142.513 6.252 ;
			RECT	142.649 6.188 142.681 6.252 ;
			RECT	142.817 6.188 142.849 6.252 ;
			RECT	142.985 6.188 143.017 6.252 ;
			RECT	143.153 6.188 143.185 6.252 ;
			RECT	143.321 6.188 143.353 6.252 ;
			RECT	143.489 6.188 143.521 6.252 ;
			RECT	143.657 6.188 143.689 6.252 ;
			RECT	143.825 6.188 143.857 6.252 ;
			RECT	143.993 6.188 144.025 6.252 ;
			RECT	144.161 6.188 144.193 6.252 ;
			RECT	144.329 6.188 144.361 6.252 ;
			RECT	144.497 6.188 144.529 6.252 ;
			RECT	144.665 6.188 144.697 6.252 ;
			RECT	144.833 6.188 144.865 6.252 ;
			RECT	145.001 6.188 145.033 6.252 ;
			RECT	145.169 6.188 145.201 6.252 ;
			RECT	145.337 6.188 145.369 6.252 ;
			RECT	145.505 6.188 145.537 6.252 ;
			RECT	145.673 6.188 145.705 6.252 ;
			RECT	145.841 6.188 145.873 6.252 ;
			RECT	146.009 6.188 146.041 6.252 ;
			RECT	146.177 6.188 146.209 6.252 ;
			RECT	146.345 6.188 146.377 6.252 ;
			RECT	146.513 6.188 146.545 6.252 ;
			RECT	146.681 6.188 146.713 6.252 ;
			RECT	146.849 6.188 146.881 6.252 ;
			RECT	147.017 6.188 147.049 6.252 ;
			RECT	147.185 6.188 147.217 6.252 ;
			RECT	147.316 6.204 147.348 6.236 ;
			RECT	147.437 6.204 147.469 6.236 ;
			RECT	147.567 6.188 147.599 6.252 ;
			RECT	149.879 6.188 149.911 6.252 ;
			RECT	151.13 6.188 151.194 6.252 ;
			RECT	151.81 6.188 151.842 6.252 ;
			RECT	152.249 6.188 152.281 6.252 ;
			RECT	153.56 6.188 153.624 6.252 ;
			RECT	156.601 6.188 156.633 6.252 ;
			RECT	156.731 6.204 156.763 6.236 ;
			RECT	156.852 6.204 156.884 6.236 ;
			RECT	156.983 6.188 157.015 6.252 ;
			RECT	157.151 6.188 157.183 6.252 ;
			RECT	157.319 6.188 157.351 6.252 ;
			RECT	157.487 6.188 157.519 6.252 ;
			RECT	157.655 6.188 157.687 6.252 ;
			RECT	157.823 6.188 157.855 6.252 ;
			RECT	157.991 6.188 158.023 6.252 ;
			RECT	158.159 6.188 158.191 6.252 ;
			RECT	158.327 6.188 158.359 6.252 ;
			RECT	158.495 6.188 158.527 6.252 ;
			RECT	158.663 6.188 158.695 6.252 ;
			RECT	158.831 6.188 158.863 6.252 ;
			RECT	158.999 6.188 159.031 6.252 ;
			RECT	159.167 6.188 159.199 6.252 ;
			RECT	159.335 6.188 159.367 6.252 ;
			RECT	159.503 6.188 159.535 6.252 ;
			RECT	159.671 6.188 159.703 6.252 ;
			RECT	159.839 6.188 159.871 6.252 ;
			RECT	160.007 6.188 160.039 6.252 ;
			RECT	160.175 6.188 160.207 6.252 ;
			RECT	160.343 6.188 160.375 6.252 ;
			RECT	160.511 6.188 160.543 6.252 ;
			RECT	160.679 6.188 160.711 6.252 ;
			RECT	160.847 6.188 160.879 6.252 ;
			RECT	161.015 6.188 161.047 6.252 ;
			RECT	161.183 6.188 161.215 6.252 ;
			RECT	161.351 6.188 161.383 6.252 ;
			RECT	161.519 6.188 161.551 6.252 ;
			RECT	161.687 6.188 161.719 6.252 ;
			RECT	161.855 6.188 161.887 6.252 ;
			RECT	162.023 6.188 162.055 6.252 ;
			RECT	162.191 6.188 162.223 6.252 ;
			RECT	162.359 6.188 162.391 6.252 ;
			RECT	162.527 6.188 162.559 6.252 ;
			RECT	162.695 6.188 162.727 6.252 ;
			RECT	162.863 6.188 162.895 6.252 ;
			RECT	163.031 6.188 163.063 6.252 ;
			RECT	163.199 6.188 163.231 6.252 ;
			RECT	163.367 6.188 163.399 6.252 ;
			RECT	163.535 6.188 163.567 6.252 ;
			RECT	163.703 6.188 163.735 6.252 ;
			RECT	163.871 6.188 163.903 6.252 ;
			RECT	164.039 6.188 164.071 6.252 ;
			RECT	164.207 6.188 164.239 6.252 ;
			RECT	164.375 6.188 164.407 6.252 ;
			RECT	164.543 6.188 164.575 6.252 ;
			RECT	164.711 6.188 164.743 6.252 ;
			RECT	164.879 6.188 164.911 6.252 ;
			RECT	165.047 6.188 165.079 6.252 ;
			RECT	165.215 6.188 165.247 6.252 ;
			RECT	165.383 6.188 165.415 6.252 ;
			RECT	165.551 6.188 165.583 6.252 ;
			RECT	165.719 6.188 165.751 6.252 ;
			RECT	165.887 6.188 165.919 6.252 ;
			RECT	166.055 6.188 166.087 6.252 ;
			RECT	166.223 6.188 166.255 6.252 ;
			RECT	166.391 6.188 166.423 6.252 ;
			RECT	166.559 6.188 166.591 6.252 ;
			RECT	166.727 6.188 166.759 6.252 ;
			RECT	166.895 6.188 166.927 6.252 ;
			RECT	167.063 6.188 167.095 6.252 ;
			RECT	167.231 6.188 167.263 6.252 ;
			RECT	167.399 6.188 167.431 6.252 ;
			RECT	167.567 6.188 167.599 6.252 ;
			RECT	167.735 6.188 167.767 6.252 ;
			RECT	167.903 6.188 167.935 6.252 ;
			RECT	168.071 6.188 168.103 6.252 ;
			RECT	168.239 6.188 168.271 6.252 ;
			RECT	168.407 6.188 168.439 6.252 ;
			RECT	168.575 6.188 168.607 6.252 ;
			RECT	168.743 6.188 168.775 6.252 ;
			RECT	168.911 6.188 168.943 6.252 ;
			RECT	169.079 6.188 169.111 6.252 ;
			RECT	169.247 6.188 169.279 6.252 ;
			RECT	169.415 6.188 169.447 6.252 ;
			RECT	169.583 6.188 169.615 6.252 ;
			RECT	169.751 6.188 169.783 6.252 ;
			RECT	169.919 6.188 169.951 6.252 ;
			RECT	170.087 6.188 170.119 6.252 ;
			RECT	170.255 6.188 170.287 6.252 ;
			RECT	170.423 6.188 170.455 6.252 ;
			RECT	170.591 6.188 170.623 6.252 ;
			RECT	170.759 6.188 170.791 6.252 ;
			RECT	170.927 6.188 170.959 6.252 ;
			RECT	171.095 6.188 171.127 6.252 ;
			RECT	171.263 6.188 171.295 6.252 ;
			RECT	171.431 6.188 171.463 6.252 ;
			RECT	171.599 6.188 171.631 6.252 ;
			RECT	171.767 6.188 171.799 6.252 ;
			RECT	171.935 6.188 171.967 6.252 ;
			RECT	172.103 6.188 172.135 6.252 ;
			RECT	172.271 6.188 172.303 6.252 ;
			RECT	172.439 6.188 172.471 6.252 ;
			RECT	172.607 6.188 172.639 6.252 ;
			RECT	172.775 6.188 172.807 6.252 ;
			RECT	172.943 6.188 172.975 6.252 ;
			RECT	173.111 6.188 173.143 6.252 ;
			RECT	173.279 6.188 173.311 6.252 ;
			RECT	173.447 6.188 173.479 6.252 ;
			RECT	173.615 6.188 173.647 6.252 ;
			RECT	173.783 6.188 173.815 6.252 ;
			RECT	173.951 6.188 173.983 6.252 ;
			RECT	174.119 6.188 174.151 6.252 ;
			RECT	174.287 6.188 174.319 6.252 ;
			RECT	174.455 6.188 174.487 6.252 ;
			RECT	174.623 6.188 174.655 6.252 ;
			RECT	174.791 6.188 174.823 6.252 ;
			RECT	174.959 6.188 174.991 6.252 ;
			RECT	175.127 6.188 175.159 6.252 ;
			RECT	175.295 6.188 175.327 6.252 ;
			RECT	175.463 6.188 175.495 6.252 ;
			RECT	175.631 6.188 175.663 6.252 ;
			RECT	175.799 6.188 175.831 6.252 ;
			RECT	175.967 6.188 175.999 6.252 ;
			RECT	176.135 6.188 176.167 6.252 ;
			RECT	176.303 6.188 176.335 6.252 ;
			RECT	176.471 6.188 176.503 6.252 ;
			RECT	176.639 6.188 176.671 6.252 ;
			RECT	176.807 6.188 176.839 6.252 ;
			RECT	176.975 6.188 177.007 6.252 ;
			RECT	177.143 6.188 177.175 6.252 ;
			RECT	177.311 6.188 177.343 6.252 ;
			RECT	177.479 6.188 177.511 6.252 ;
			RECT	177.647 6.188 177.679 6.252 ;
			RECT	177.815 6.188 177.847 6.252 ;
			RECT	177.983 6.188 178.015 6.252 ;
			RECT	178.151 6.188 178.183 6.252 ;
			RECT	178.319 6.188 178.351 6.252 ;
			RECT	178.487 6.188 178.519 6.252 ;
			RECT	178.655 6.188 178.687 6.252 ;
			RECT	178.823 6.188 178.855 6.252 ;
			RECT	178.991 6.188 179.023 6.252 ;
			RECT	179.159 6.188 179.191 6.252 ;
			RECT	179.327 6.188 179.359 6.252 ;
			RECT	179.495 6.188 179.527 6.252 ;
			RECT	179.663 6.188 179.695 6.252 ;
			RECT	179.831 6.188 179.863 6.252 ;
			RECT	179.999 6.188 180.031 6.252 ;
			RECT	180.167 6.188 180.199 6.252 ;
			RECT	180.335 6.188 180.367 6.252 ;
			RECT	180.503 6.188 180.535 6.252 ;
			RECT	180.671 6.188 180.703 6.252 ;
			RECT	180.839 6.188 180.871 6.252 ;
			RECT	181.007 6.188 181.039 6.252 ;
			RECT	181.175 6.188 181.207 6.252 ;
			RECT	181.343 6.188 181.375 6.252 ;
			RECT	181.511 6.188 181.543 6.252 ;
			RECT	181.679 6.188 181.711 6.252 ;
			RECT	181.847 6.188 181.879 6.252 ;
			RECT	182.015 6.188 182.047 6.252 ;
			RECT	182.183 6.188 182.215 6.252 ;
			RECT	182.351 6.188 182.383 6.252 ;
			RECT	182.519 6.188 182.551 6.252 ;
			RECT	182.687 6.188 182.719 6.252 ;
			RECT	182.855 6.188 182.887 6.252 ;
			RECT	183.023 6.188 183.055 6.252 ;
			RECT	183.191 6.188 183.223 6.252 ;
			RECT	183.359 6.188 183.391 6.252 ;
			RECT	183.527 6.188 183.559 6.252 ;
			RECT	183.695 6.188 183.727 6.252 ;
			RECT	183.863 6.188 183.895 6.252 ;
			RECT	184.031 6.188 184.063 6.252 ;
			RECT	184.199 6.188 184.231 6.252 ;
			RECT	184.367 6.188 184.399 6.252 ;
			RECT	184.535 6.188 184.567 6.252 ;
			RECT	184.703 6.188 184.735 6.252 ;
			RECT	184.871 6.188 184.903 6.252 ;
			RECT	185.039 6.188 185.071 6.252 ;
			RECT	185.207 6.188 185.239 6.252 ;
			RECT	185.375 6.188 185.407 6.252 ;
			RECT	185.543 6.188 185.575 6.252 ;
			RECT	185.711 6.188 185.743 6.252 ;
			RECT	185.879 6.188 185.911 6.252 ;
			RECT	186.047 6.188 186.079 6.252 ;
			RECT	186.215 6.188 186.247 6.252 ;
			RECT	186.383 6.188 186.415 6.252 ;
			RECT	186.551 6.188 186.583 6.252 ;
			RECT	186.719 6.188 186.751 6.252 ;
			RECT	186.887 6.188 186.919 6.252 ;
			RECT	187.055 6.188 187.087 6.252 ;
			RECT	187.223 6.188 187.255 6.252 ;
			RECT	187.391 6.188 187.423 6.252 ;
			RECT	187.559 6.188 187.591 6.252 ;
			RECT	187.727 6.188 187.759 6.252 ;
			RECT	187.895 6.188 187.927 6.252 ;
			RECT	188.063 6.188 188.095 6.252 ;
			RECT	188.231 6.188 188.263 6.252 ;
			RECT	188.399 6.188 188.431 6.252 ;
			RECT	188.567 6.188 188.599 6.252 ;
			RECT	188.735 6.188 188.767 6.252 ;
			RECT	188.903 6.188 188.935 6.252 ;
			RECT	189.071 6.188 189.103 6.252 ;
			RECT	189.239 6.188 189.271 6.252 ;
			RECT	189.407 6.188 189.439 6.252 ;
			RECT	189.575 6.188 189.607 6.252 ;
			RECT	189.743 6.188 189.775 6.252 ;
			RECT	189.911 6.188 189.943 6.252 ;
			RECT	190.079 6.188 190.111 6.252 ;
			RECT	190.247 6.188 190.279 6.252 ;
			RECT	190.415 6.188 190.447 6.252 ;
			RECT	190.583 6.188 190.615 6.252 ;
			RECT	190.751 6.188 190.783 6.252 ;
			RECT	190.919 6.188 190.951 6.252 ;
			RECT	191.087 6.188 191.119 6.252 ;
			RECT	191.255 6.188 191.287 6.252 ;
			RECT	191.423 6.188 191.455 6.252 ;
			RECT	191.591 6.188 191.623 6.252 ;
			RECT	191.759 6.188 191.791 6.252 ;
			RECT	191.927 6.188 191.959 6.252 ;
			RECT	192.095 6.188 192.127 6.252 ;
			RECT	192.263 6.188 192.295 6.252 ;
			RECT	192.431 6.188 192.463 6.252 ;
			RECT	192.599 6.188 192.631 6.252 ;
			RECT	192.767 6.188 192.799 6.252 ;
			RECT	192.935 6.188 192.967 6.252 ;
			RECT	193.103 6.188 193.135 6.252 ;
			RECT	193.271 6.188 193.303 6.252 ;
			RECT	193.439 6.188 193.471 6.252 ;
			RECT	193.607 6.188 193.639 6.252 ;
			RECT	193.775 6.188 193.807 6.252 ;
			RECT	193.943 6.188 193.975 6.252 ;
			RECT	194.111 6.188 194.143 6.252 ;
			RECT	194.279 6.188 194.311 6.252 ;
			RECT	194.447 6.188 194.479 6.252 ;
			RECT	194.615 6.188 194.647 6.252 ;
			RECT	194.783 6.188 194.815 6.252 ;
			RECT	194.951 6.188 194.983 6.252 ;
			RECT	195.119 6.188 195.151 6.252 ;
			RECT	195.287 6.188 195.319 6.252 ;
			RECT	195.455 6.188 195.487 6.252 ;
			RECT	195.623 6.188 195.655 6.252 ;
			RECT	195.791 6.188 195.823 6.252 ;
			RECT	195.959 6.188 195.991 6.252 ;
			RECT	196.127 6.188 196.159 6.252 ;
			RECT	196.295 6.188 196.327 6.252 ;
			RECT	196.463 6.188 196.495 6.252 ;
			RECT	196.631 6.188 196.663 6.252 ;
			RECT	196.799 6.188 196.831 6.252 ;
			RECT	196.967 6.188 196.999 6.252 ;
			RECT	197.135 6.188 197.167 6.252 ;
			RECT	197.303 6.188 197.335 6.252 ;
			RECT	197.471 6.188 197.503 6.252 ;
			RECT	197.639 6.188 197.671 6.252 ;
			RECT	197.807 6.188 197.839 6.252 ;
			RECT	197.975 6.188 198.007 6.252 ;
			RECT	198.143 6.188 198.175 6.252 ;
			RECT	198.311 6.188 198.343 6.252 ;
			RECT	198.479 6.188 198.511 6.252 ;
			RECT	198.647 6.188 198.679 6.252 ;
			RECT	198.815 6.188 198.847 6.252 ;
			RECT	198.983 6.188 199.015 6.252 ;
			RECT	199.151 6.188 199.183 6.252 ;
			RECT	199.319 6.188 199.351 6.252 ;
			RECT	199.487 6.188 199.519 6.252 ;
			RECT	199.655 6.188 199.687 6.252 ;
			RECT	199.823 6.188 199.855 6.252 ;
			RECT	199.991 6.188 200.023 6.252 ;
			RECT	200.121 6.204 200.153 6.236 ;
			RECT	200.243 6.209 200.275 6.241 ;
			RECT	200.373 6.188 200.405 6.252 ;
			RECT	200.9 6.188 200.932 6.252 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 4.24 201.665 4.36 ;
			LAYER	J3 ;
			RECT	0.755 4.268 0.787 4.332 ;
			RECT	1.645 4.268 1.709 4.332 ;
			RECT	2.323 4.268 2.387 4.332 ;
			RECT	3.438 4.268 3.47 4.332 ;
			RECT	3.585 4.268 3.617 4.332 ;
			RECT	4.195 4.268 4.227 4.332 ;
			RECT	4.72 4.268 4.752 4.332 ;
			RECT	4.944 4.268 5.008 4.332 ;
			RECT	5.267 4.268 5.299 4.332 ;
			RECT	5.797 4.268 5.829 4.332 ;
			RECT	5.927 4.289 5.959 4.321 ;
			RECT	6.049 4.284 6.081 4.316 ;
			RECT	6.179 4.268 6.211 4.332 ;
			RECT	6.347 4.268 6.379 4.332 ;
			RECT	6.515 4.268 6.547 4.332 ;
			RECT	6.683 4.268 6.715 4.332 ;
			RECT	6.851 4.268 6.883 4.332 ;
			RECT	7.019 4.268 7.051 4.332 ;
			RECT	7.187 4.268 7.219 4.332 ;
			RECT	7.355 4.268 7.387 4.332 ;
			RECT	7.523 4.268 7.555 4.332 ;
			RECT	7.691 4.268 7.723 4.332 ;
			RECT	7.859 4.268 7.891 4.332 ;
			RECT	8.027 4.268 8.059 4.332 ;
			RECT	8.195 4.268 8.227 4.332 ;
			RECT	8.363 4.268 8.395 4.332 ;
			RECT	8.531 4.268 8.563 4.332 ;
			RECT	8.699 4.268 8.731 4.332 ;
			RECT	8.867 4.268 8.899 4.332 ;
			RECT	9.035 4.268 9.067 4.332 ;
			RECT	9.203 4.268 9.235 4.332 ;
			RECT	9.371 4.268 9.403 4.332 ;
			RECT	9.539 4.268 9.571 4.332 ;
			RECT	9.707 4.268 9.739 4.332 ;
			RECT	9.875 4.268 9.907 4.332 ;
			RECT	10.043 4.268 10.075 4.332 ;
			RECT	10.211 4.268 10.243 4.332 ;
			RECT	10.379 4.268 10.411 4.332 ;
			RECT	10.547 4.268 10.579 4.332 ;
			RECT	10.715 4.268 10.747 4.332 ;
			RECT	10.883 4.268 10.915 4.332 ;
			RECT	11.051 4.268 11.083 4.332 ;
			RECT	11.219 4.268 11.251 4.332 ;
			RECT	11.387 4.268 11.419 4.332 ;
			RECT	11.555 4.268 11.587 4.332 ;
			RECT	11.723 4.268 11.755 4.332 ;
			RECT	11.891 4.268 11.923 4.332 ;
			RECT	12.059 4.268 12.091 4.332 ;
			RECT	12.227 4.268 12.259 4.332 ;
			RECT	12.395 4.268 12.427 4.332 ;
			RECT	12.563 4.268 12.595 4.332 ;
			RECT	12.731 4.268 12.763 4.332 ;
			RECT	12.899 4.268 12.931 4.332 ;
			RECT	13.067 4.268 13.099 4.332 ;
			RECT	13.235 4.268 13.267 4.332 ;
			RECT	13.403 4.268 13.435 4.332 ;
			RECT	13.571 4.268 13.603 4.332 ;
			RECT	13.739 4.268 13.771 4.332 ;
			RECT	13.907 4.268 13.939 4.332 ;
			RECT	14.075 4.268 14.107 4.332 ;
			RECT	14.243 4.268 14.275 4.332 ;
			RECT	14.411 4.268 14.443 4.332 ;
			RECT	14.579 4.268 14.611 4.332 ;
			RECT	14.747 4.268 14.779 4.332 ;
			RECT	14.915 4.268 14.947 4.332 ;
			RECT	15.083 4.268 15.115 4.332 ;
			RECT	15.251 4.268 15.283 4.332 ;
			RECT	15.419 4.268 15.451 4.332 ;
			RECT	15.587 4.268 15.619 4.332 ;
			RECT	15.755 4.268 15.787 4.332 ;
			RECT	15.923 4.268 15.955 4.332 ;
			RECT	16.091 4.268 16.123 4.332 ;
			RECT	16.259 4.268 16.291 4.332 ;
			RECT	16.427 4.268 16.459 4.332 ;
			RECT	16.595 4.268 16.627 4.332 ;
			RECT	16.763 4.268 16.795 4.332 ;
			RECT	16.931 4.268 16.963 4.332 ;
			RECT	17.099 4.268 17.131 4.332 ;
			RECT	17.267 4.268 17.299 4.332 ;
			RECT	17.435 4.268 17.467 4.332 ;
			RECT	17.603 4.268 17.635 4.332 ;
			RECT	17.771 4.268 17.803 4.332 ;
			RECT	17.939 4.268 17.971 4.332 ;
			RECT	18.107 4.268 18.139 4.332 ;
			RECT	18.275 4.268 18.307 4.332 ;
			RECT	18.443 4.268 18.475 4.332 ;
			RECT	18.611 4.268 18.643 4.332 ;
			RECT	18.779 4.268 18.811 4.332 ;
			RECT	18.947 4.268 18.979 4.332 ;
			RECT	19.115 4.268 19.147 4.332 ;
			RECT	19.283 4.268 19.315 4.332 ;
			RECT	19.451 4.268 19.483 4.332 ;
			RECT	19.619 4.268 19.651 4.332 ;
			RECT	19.787 4.268 19.819 4.332 ;
			RECT	19.955 4.268 19.987 4.332 ;
			RECT	20.123 4.268 20.155 4.332 ;
			RECT	20.291 4.268 20.323 4.332 ;
			RECT	20.459 4.268 20.491 4.332 ;
			RECT	20.627 4.268 20.659 4.332 ;
			RECT	20.795 4.268 20.827 4.332 ;
			RECT	20.963 4.268 20.995 4.332 ;
			RECT	21.131 4.268 21.163 4.332 ;
			RECT	21.299 4.268 21.331 4.332 ;
			RECT	21.467 4.268 21.499 4.332 ;
			RECT	21.635 4.268 21.667 4.332 ;
			RECT	21.803 4.268 21.835 4.332 ;
			RECT	21.971 4.268 22.003 4.332 ;
			RECT	22.139 4.268 22.171 4.332 ;
			RECT	22.307 4.268 22.339 4.332 ;
			RECT	22.475 4.268 22.507 4.332 ;
			RECT	22.643 4.268 22.675 4.332 ;
			RECT	22.811 4.268 22.843 4.332 ;
			RECT	22.979 4.268 23.011 4.332 ;
			RECT	23.147 4.268 23.179 4.332 ;
			RECT	23.315 4.268 23.347 4.332 ;
			RECT	23.483 4.268 23.515 4.332 ;
			RECT	23.651 4.268 23.683 4.332 ;
			RECT	23.819 4.268 23.851 4.332 ;
			RECT	23.987 4.268 24.019 4.332 ;
			RECT	24.155 4.268 24.187 4.332 ;
			RECT	24.323 4.268 24.355 4.332 ;
			RECT	24.491 4.268 24.523 4.332 ;
			RECT	24.659 4.268 24.691 4.332 ;
			RECT	24.827 4.268 24.859 4.332 ;
			RECT	24.995 4.268 25.027 4.332 ;
			RECT	25.163 4.268 25.195 4.332 ;
			RECT	25.331 4.268 25.363 4.332 ;
			RECT	25.499 4.268 25.531 4.332 ;
			RECT	25.667 4.268 25.699 4.332 ;
			RECT	25.835 4.268 25.867 4.332 ;
			RECT	26.003 4.268 26.035 4.332 ;
			RECT	26.171 4.268 26.203 4.332 ;
			RECT	26.339 4.268 26.371 4.332 ;
			RECT	26.507 4.268 26.539 4.332 ;
			RECT	26.675 4.268 26.707 4.332 ;
			RECT	26.843 4.268 26.875 4.332 ;
			RECT	27.011 4.268 27.043 4.332 ;
			RECT	27.179 4.268 27.211 4.332 ;
			RECT	27.347 4.268 27.379 4.332 ;
			RECT	27.515 4.268 27.547 4.332 ;
			RECT	27.683 4.268 27.715 4.332 ;
			RECT	27.851 4.268 27.883 4.332 ;
			RECT	28.019 4.268 28.051 4.332 ;
			RECT	28.187 4.268 28.219 4.332 ;
			RECT	28.355 4.268 28.387 4.332 ;
			RECT	28.523 4.268 28.555 4.332 ;
			RECT	28.691 4.268 28.723 4.332 ;
			RECT	28.859 4.268 28.891 4.332 ;
			RECT	29.027 4.268 29.059 4.332 ;
			RECT	29.195 4.268 29.227 4.332 ;
			RECT	29.363 4.268 29.395 4.332 ;
			RECT	29.531 4.268 29.563 4.332 ;
			RECT	29.699 4.268 29.731 4.332 ;
			RECT	29.867 4.268 29.899 4.332 ;
			RECT	30.035 4.268 30.067 4.332 ;
			RECT	30.203 4.268 30.235 4.332 ;
			RECT	30.371 4.268 30.403 4.332 ;
			RECT	30.539 4.268 30.571 4.332 ;
			RECT	30.707 4.268 30.739 4.332 ;
			RECT	30.875 4.268 30.907 4.332 ;
			RECT	31.043 4.268 31.075 4.332 ;
			RECT	31.211 4.268 31.243 4.332 ;
			RECT	31.379 4.268 31.411 4.332 ;
			RECT	31.547 4.268 31.579 4.332 ;
			RECT	31.715 4.268 31.747 4.332 ;
			RECT	31.883 4.268 31.915 4.332 ;
			RECT	32.051 4.268 32.083 4.332 ;
			RECT	32.219 4.268 32.251 4.332 ;
			RECT	32.387 4.268 32.419 4.332 ;
			RECT	32.555 4.268 32.587 4.332 ;
			RECT	32.723 4.268 32.755 4.332 ;
			RECT	32.891 4.268 32.923 4.332 ;
			RECT	33.059 4.268 33.091 4.332 ;
			RECT	33.227 4.268 33.259 4.332 ;
			RECT	33.395 4.268 33.427 4.332 ;
			RECT	33.563 4.268 33.595 4.332 ;
			RECT	33.731 4.268 33.763 4.332 ;
			RECT	33.899 4.268 33.931 4.332 ;
			RECT	34.067 4.268 34.099 4.332 ;
			RECT	34.235 4.268 34.267 4.332 ;
			RECT	34.403 4.268 34.435 4.332 ;
			RECT	34.571 4.268 34.603 4.332 ;
			RECT	34.739 4.268 34.771 4.332 ;
			RECT	34.907 4.268 34.939 4.332 ;
			RECT	35.075 4.268 35.107 4.332 ;
			RECT	35.243 4.268 35.275 4.332 ;
			RECT	35.411 4.268 35.443 4.332 ;
			RECT	35.579 4.268 35.611 4.332 ;
			RECT	35.747 4.268 35.779 4.332 ;
			RECT	35.915 4.268 35.947 4.332 ;
			RECT	36.083 4.268 36.115 4.332 ;
			RECT	36.251 4.268 36.283 4.332 ;
			RECT	36.419 4.268 36.451 4.332 ;
			RECT	36.587 4.268 36.619 4.332 ;
			RECT	36.755 4.268 36.787 4.332 ;
			RECT	36.923 4.268 36.955 4.332 ;
			RECT	37.091 4.268 37.123 4.332 ;
			RECT	37.259 4.268 37.291 4.332 ;
			RECT	37.427 4.268 37.459 4.332 ;
			RECT	37.595 4.268 37.627 4.332 ;
			RECT	37.763 4.268 37.795 4.332 ;
			RECT	37.931 4.268 37.963 4.332 ;
			RECT	38.099 4.268 38.131 4.332 ;
			RECT	38.267 4.268 38.299 4.332 ;
			RECT	38.435 4.268 38.467 4.332 ;
			RECT	38.603 4.268 38.635 4.332 ;
			RECT	38.771 4.268 38.803 4.332 ;
			RECT	38.939 4.268 38.971 4.332 ;
			RECT	39.107 4.268 39.139 4.332 ;
			RECT	39.275 4.268 39.307 4.332 ;
			RECT	39.443 4.268 39.475 4.332 ;
			RECT	39.611 4.268 39.643 4.332 ;
			RECT	39.779 4.268 39.811 4.332 ;
			RECT	39.947 4.268 39.979 4.332 ;
			RECT	40.115 4.268 40.147 4.332 ;
			RECT	40.283 4.268 40.315 4.332 ;
			RECT	40.451 4.268 40.483 4.332 ;
			RECT	40.619 4.268 40.651 4.332 ;
			RECT	40.787 4.268 40.819 4.332 ;
			RECT	40.955 4.268 40.987 4.332 ;
			RECT	41.123 4.268 41.155 4.332 ;
			RECT	41.291 4.268 41.323 4.332 ;
			RECT	41.459 4.268 41.491 4.332 ;
			RECT	41.627 4.268 41.659 4.332 ;
			RECT	41.795 4.268 41.827 4.332 ;
			RECT	41.963 4.268 41.995 4.332 ;
			RECT	42.131 4.268 42.163 4.332 ;
			RECT	42.299 4.268 42.331 4.332 ;
			RECT	42.467 4.268 42.499 4.332 ;
			RECT	42.635 4.268 42.667 4.332 ;
			RECT	42.803 4.268 42.835 4.332 ;
			RECT	42.971 4.268 43.003 4.332 ;
			RECT	43.139 4.268 43.171 4.332 ;
			RECT	43.307 4.268 43.339 4.332 ;
			RECT	43.475 4.268 43.507 4.332 ;
			RECT	43.643 4.268 43.675 4.332 ;
			RECT	43.811 4.268 43.843 4.332 ;
			RECT	43.979 4.268 44.011 4.332 ;
			RECT	44.147 4.268 44.179 4.332 ;
			RECT	44.315 4.268 44.347 4.332 ;
			RECT	44.483 4.268 44.515 4.332 ;
			RECT	44.651 4.268 44.683 4.332 ;
			RECT	44.819 4.268 44.851 4.332 ;
			RECT	44.987 4.268 45.019 4.332 ;
			RECT	45.155 4.268 45.187 4.332 ;
			RECT	45.323 4.268 45.355 4.332 ;
			RECT	45.491 4.268 45.523 4.332 ;
			RECT	45.659 4.268 45.691 4.332 ;
			RECT	45.827 4.268 45.859 4.332 ;
			RECT	45.995 4.268 46.027 4.332 ;
			RECT	46.163 4.268 46.195 4.332 ;
			RECT	46.331 4.268 46.363 4.332 ;
			RECT	46.499 4.268 46.531 4.332 ;
			RECT	46.667 4.268 46.699 4.332 ;
			RECT	46.835 4.268 46.867 4.332 ;
			RECT	47.003 4.268 47.035 4.332 ;
			RECT	47.171 4.268 47.203 4.332 ;
			RECT	47.339 4.268 47.371 4.332 ;
			RECT	47.507 4.268 47.539 4.332 ;
			RECT	47.675 4.268 47.707 4.332 ;
			RECT	47.843 4.268 47.875 4.332 ;
			RECT	48.011 4.268 48.043 4.332 ;
			RECT	48.179 4.268 48.211 4.332 ;
			RECT	48.347 4.268 48.379 4.332 ;
			RECT	48.515 4.268 48.547 4.332 ;
			RECT	48.683 4.268 48.715 4.332 ;
			RECT	48.851 4.268 48.883 4.332 ;
			RECT	49.019 4.268 49.051 4.332 ;
			RECT	49.187 4.268 49.219 4.332 ;
			RECT	49.318 4.284 49.35 4.316 ;
			RECT	49.439 4.284 49.471 4.316 ;
			RECT	49.569 4.268 49.601 4.332 ;
			RECT	51.881 4.268 51.913 4.332 ;
			RECT	53.132 4.268 53.196 4.332 ;
			RECT	53.812 4.268 53.844 4.332 ;
			RECT	54.251 4.268 54.283 4.332 ;
			RECT	55.562 4.268 55.626 4.332 ;
			RECT	58.603 4.268 58.635 4.332 ;
			RECT	58.733 4.284 58.765 4.316 ;
			RECT	58.854 4.284 58.886 4.316 ;
			RECT	58.985 4.268 59.017 4.332 ;
			RECT	59.153 4.268 59.185 4.332 ;
			RECT	59.321 4.268 59.353 4.332 ;
			RECT	59.489 4.268 59.521 4.332 ;
			RECT	59.657 4.268 59.689 4.332 ;
			RECT	59.825 4.268 59.857 4.332 ;
			RECT	59.993 4.268 60.025 4.332 ;
			RECT	60.161 4.268 60.193 4.332 ;
			RECT	60.329 4.268 60.361 4.332 ;
			RECT	60.497 4.268 60.529 4.332 ;
			RECT	60.665 4.268 60.697 4.332 ;
			RECT	60.833 4.268 60.865 4.332 ;
			RECT	61.001 4.268 61.033 4.332 ;
			RECT	61.169 4.268 61.201 4.332 ;
			RECT	61.337 4.268 61.369 4.332 ;
			RECT	61.505 4.268 61.537 4.332 ;
			RECT	61.673 4.268 61.705 4.332 ;
			RECT	61.841 4.268 61.873 4.332 ;
			RECT	62.009 4.268 62.041 4.332 ;
			RECT	62.177 4.268 62.209 4.332 ;
			RECT	62.345 4.268 62.377 4.332 ;
			RECT	62.513 4.268 62.545 4.332 ;
			RECT	62.681 4.268 62.713 4.332 ;
			RECT	62.849 4.268 62.881 4.332 ;
			RECT	63.017 4.268 63.049 4.332 ;
			RECT	63.185 4.268 63.217 4.332 ;
			RECT	63.353 4.268 63.385 4.332 ;
			RECT	63.521 4.268 63.553 4.332 ;
			RECT	63.689 4.268 63.721 4.332 ;
			RECT	63.857 4.268 63.889 4.332 ;
			RECT	64.025 4.268 64.057 4.332 ;
			RECT	64.193 4.268 64.225 4.332 ;
			RECT	64.361 4.268 64.393 4.332 ;
			RECT	64.529 4.268 64.561 4.332 ;
			RECT	64.697 4.268 64.729 4.332 ;
			RECT	64.865 4.268 64.897 4.332 ;
			RECT	65.033 4.268 65.065 4.332 ;
			RECT	65.201 4.268 65.233 4.332 ;
			RECT	65.369 4.268 65.401 4.332 ;
			RECT	65.537 4.268 65.569 4.332 ;
			RECT	65.705 4.268 65.737 4.332 ;
			RECT	65.873 4.268 65.905 4.332 ;
			RECT	66.041 4.268 66.073 4.332 ;
			RECT	66.209 4.268 66.241 4.332 ;
			RECT	66.377 4.268 66.409 4.332 ;
			RECT	66.545 4.268 66.577 4.332 ;
			RECT	66.713 4.268 66.745 4.332 ;
			RECT	66.881 4.268 66.913 4.332 ;
			RECT	67.049 4.268 67.081 4.332 ;
			RECT	67.217 4.268 67.249 4.332 ;
			RECT	67.385 4.268 67.417 4.332 ;
			RECT	67.553 4.268 67.585 4.332 ;
			RECT	67.721 4.268 67.753 4.332 ;
			RECT	67.889 4.268 67.921 4.332 ;
			RECT	68.057 4.268 68.089 4.332 ;
			RECT	68.225 4.268 68.257 4.332 ;
			RECT	68.393 4.268 68.425 4.332 ;
			RECT	68.561 4.268 68.593 4.332 ;
			RECT	68.729 4.268 68.761 4.332 ;
			RECT	68.897 4.268 68.929 4.332 ;
			RECT	69.065 4.268 69.097 4.332 ;
			RECT	69.233 4.268 69.265 4.332 ;
			RECT	69.401 4.268 69.433 4.332 ;
			RECT	69.569 4.268 69.601 4.332 ;
			RECT	69.737 4.268 69.769 4.332 ;
			RECT	69.905 4.268 69.937 4.332 ;
			RECT	70.073 4.268 70.105 4.332 ;
			RECT	70.241 4.268 70.273 4.332 ;
			RECT	70.409 4.268 70.441 4.332 ;
			RECT	70.577 4.268 70.609 4.332 ;
			RECT	70.745 4.268 70.777 4.332 ;
			RECT	70.913 4.268 70.945 4.332 ;
			RECT	71.081 4.268 71.113 4.332 ;
			RECT	71.249 4.268 71.281 4.332 ;
			RECT	71.417 4.268 71.449 4.332 ;
			RECT	71.585 4.268 71.617 4.332 ;
			RECT	71.753 4.268 71.785 4.332 ;
			RECT	71.921 4.268 71.953 4.332 ;
			RECT	72.089 4.268 72.121 4.332 ;
			RECT	72.257 4.268 72.289 4.332 ;
			RECT	72.425 4.268 72.457 4.332 ;
			RECT	72.593 4.268 72.625 4.332 ;
			RECT	72.761 4.268 72.793 4.332 ;
			RECT	72.929 4.268 72.961 4.332 ;
			RECT	73.097 4.268 73.129 4.332 ;
			RECT	73.265 4.268 73.297 4.332 ;
			RECT	73.433 4.268 73.465 4.332 ;
			RECT	73.601 4.268 73.633 4.332 ;
			RECT	73.769 4.268 73.801 4.332 ;
			RECT	73.937 4.268 73.969 4.332 ;
			RECT	74.105 4.268 74.137 4.332 ;
			RECT	74.273 4.268 74.305 4.332 ;
			RECT	74.441 4.268 74.473 4.332 ;
			RECT	74.609 4.268 74.641 4.332 ;
			RECT	74.777 4.268 74.809 4.332 ;
			RECT	74.945 4.268 74.977 4.332 ;
			RECT	75.113 4.268 75.145 4.332 ;
			RECT	75.281 4.268 75.313 4.332 ;
			RECT	75.449 4.268 75.481 4.332 ;
			RECT	75.617 4.268 75.649 4.332 ;
			RECT	75.785 4.268 75.817 4.332 ;
			RECT	75.953 4.268 75.985 4.332 ;
			RECT	76.121 4.268 76.153 4.332 ;
			RECT	76.289 4.268 76.321 4.332 ;
			RECT	76.457 4.268 76.489 4.332 ;
			RECT	76.625 4.268 76.657 4.332 ;
			RECT	76.793 4.268 76.825 4.332 ;
			RECT	76.961 4.268 76.993 4.332 ;
			RECT	77.129 4.268 77.161 4.332 ;
			RECT	77.297 4.268 77.329 4.332 ;
			RECT	77.465 4.268 77.497 4.332 ;
			RECT	77.633 4.268 77.665 4.332 ;
			RECT	77.801 4.268 77.833 4.332 ;
			RECT	77.969 4.268 78.001 4.332 ;
			RECT	78.137 4.268 78.169 4.332 ;
			RECT	78.305 4.268 78.337 4.332 ;
			RECT	78.473 4.268 78.505 4.332 ;
			RECT	78.641 4.268 78.673 4.332 ;
			RECT	78.809 4.268 78.841 4.332 ;
			RECT	78.977 4.268 79.009 4.332 ;
			RECT	79.145 4.268 79.177 4.332 ;
			RECT	79.313 4.268 79.345 4.332 ;
			RECT	79.481 4.268 79.513 4.332 ;
			RECT	79.649 4.268 79.681 4.332 ;
			RECT	79.817 4.268 79.849 4.332 ;
			RECT	79.985 4.268 80.017 4.332 ;
			RECT	80.153 4.268 80.185 4.332 ;
			RECT	80.321 4.268 80.353 4.332 ;
			RECT	80.489 4.268 80.521 4.332 ;
			RECT	80.657 4.268 80.689 4.332 ;
			RECT	80.825 4.268 80.857 4.332 ;
			RECT	80.993 4.268 81.025 4.332 ;
			RECT	81.161 4.268 81.193 4.332 ;
			RECT	81.329 4.268 81.361 4.332 ;
			RECT	81.497 4.268 81.529 4.332 ;
			RECT	81.665 4.268 81.697 4.332 ;
			RECT	81.833 4.268 81.865 4.332 ;
			RECT	82.001 4.268 82.033 4.332 ;
			RECT	82.169 4.268 82.201 4.332 ;
			RECT	82.337 4.268 82.369 4.332 ;
			RECT	82.505 4.268 82.537 4.332 ;
			RECT	82.673 4.268 82.705 4.332 ;
			RECT	82.841 4.268 82.873 4.332 ;
			RECT	83.009 4.268 83.041 4.332 ;
			RECT	83.177 4.268 83.209 4.332 ;
			RECT	83.345 4.268 83.377 4.332 ;
			RECT	83.513 4.268 83.545 4.332 ;
			RECT	83.681 4.268 83.713 4.332 ;
			RECT	83.849 4.268 83.881 4.332 ;
			RECT	84.017 4.268 84.049 4.332 ;
			RECT	84.185 4.268 84.217 4.332 ;
			RECT	84.353 4.268 84.385 4.332 ;
			RECT	84.521 4.268 84.553 4.332 ;
			RECT	84.689 4.268 84.721 4.332 ;
			RECT	84.857 4.268 84.889 4.332 ;
			RECT	85.025 4.268 85.057 4.332 ;
			RECT	85.193 4.268 85.225 4.332 ;
			RECT	85.361 4.268 85.393 4.332 ;
			RECT	85.529 4.268 85.561 4.332 ;
			RECT	85.697 4.268 85.729 4.332 ;
			RECT	85.865 4.268 85.897 4.332 ;
			RECT	86.033 4.268 86.065 4.332 ;
			RECT	86.201 4.268 86.233 4.332 ;
			RECT	86.369 4.268 86.401 4.332 ;
			RECT	86.537 4.268 86.569 4.332 ;
			RECT	86.705 4.268 86.737 4.332 ;
			RECT	86.873 4.268 86.905 4.332 ;
			RECT	87.041 4.268 87.073 4.332 ;
			RECT	87.209 4.268 87.241 4.332 ;
			RECT	87.377 4.268 87.409 4.332 ;
			RECT	87.545 4.268 87.577 4.332 ;
			RECT	87.713 4.268 87.745 4.332 ;
			RECT	87.881 4.268 87.913 4.332 ;
			RECT	88.049 4.268 88.081 4.332 ;
			RECT	88.217 4.268 88.249 4.332 ;
			RECT	88.385 4.268 88.417 4.332 ;
			RECT	88.553 4.268 88.585 4.332 ;
			RECT	88.721 4.268 88.753 4.332 ;
			RECT	88.889 4.268 88.921 4.332 ;
			RECT	89.057 4.268 89.089 4.332 ;
			RECT	89.225 4.268 89.257 4.332 ;
			RECT	89.393 4.268 89.425 4.332 ;
			RECT	89.561 4.268 89.593 4.332 ;
			RECT	89.729 4.268 89.761 4.332 ;
			RECT	89.897 4.268 89.929 4.332 ;
			RECT	90.065 4.268 90.097 4.332 ;
			RECT	90.233 4.268 90.265 4.332 ;
			RECT	90.401 4.268 90.433 4.332 ;
			RECT	90.569 4.268 90.601 4.332 ;
			RECT	90.737 4.268 90.769 4.332 ;
			RECT	90.905 4.268 90.937 4.332 ;
			RECT	91.073 4.268 91.105 4.332 ;
			RECT	91.241 4.268 91.273 4.332 ;
			RECT	91.409 4.268 91.441 4.332 ;
			RECT	91.577 4.268 91.609 4.332 ;
			RECT	91.745 4.268 91.777 4.332 ;
			RECT	91.913 4.268 91.945 4.332 ;
			RECT	92.081 4.268 92.113 4.332 ;
			RECT	92.249 4.268 92.281 4.332 ;
			RECT	92.417 4.268 92.449 4.332 ;
			RECT	92.585 4.268 92.617 4.332 ;
			RECT	92.753 4.268 92.785 4.332 ;
			RECT	92.921 4.268 92.953 4.332 ;
			RECT	93.089 4.268 93.121 4.332 ;
			RECT	93.257 4.268 93.289 4.332 ;
			RECT	93.425 4.268 93.457 4.332 ;
			RECT	93.593 4.268 93.625 4.332 ;
			RECT	93.761 4.268 93.793 4.332 ;
			RECT	93.929 4.268 93.961 4.332 ;
			RECT	94.097 4.268 94.129 4.332 ;
			RECT	94.265 4.268 94.297 4.332 ;
			RECT	94.433 4.268 94.465 4.332 ;
			RECT	94.601 4.268 94.633 4.332 ;
			RECT	94.769 4.268 94.801 4.332 ;
			RECT	94.937 4.268 94.969 4.332 ;
			RECT	95.105 4.268 95.137 4.332 ;
			RECT	95.273 4.268 95.305 4.332 ;
			RECT	95.441 4.268 95.473 4.332 ;
			RECT	95.609 4.268 95.641 4.332 ;
			RECT	95.777 4.268 95.809 4.332 ;
			RECT	95.945 4.268 95.977 4.332 ;
			RECT	96.113 4.268 96.145 4.332 ;
			RECT	96.281 4.268 96.313 4.332 ;
			RECT	96.449 4.268 96.481 4.332 ;
			RECT	96.617 4.268 96.649 4.332 ;
			RECT	96.785 4.268 96.817 4.332 ;
			RECT	96.953 4.268 96.985 4.332 ;
			RECT	97.121 4.268 97.153 4.332 ;
			RECT	97.289 4.268 97.321 4.332 ;
			RECT	97.457 4.268 97.489 4.332 ;
			RECT	97.625 4.268 97.657 4.332 ;
			RECT	97.793 4.268 97.825 4.332 ;
			RECT	97.961 4.268 97.993 4.332 ;
			RECT	98.129 4.268 98.161 4.332 ;
			RECT	98.297 4.268 98.329 4.332 ;
			RECT	98.465 4.268 98.497 4.332 ;
			RECT	98.633 4.268 98.665 4.332 ;
			RECT	98.801 4.268 98.833 4.332 ;
			RECT	98.969 4.268 99.001 4.332 ;
			RECT	99.137 4.268 99.169 4.332 ;
			RECT	99.305 4.268 99.337 4.332 ;
			RECT	99.473 4.268 99.505 4.332 ;
			RECT	99.641 4.268 99.673 4.332 ;
			RECT	99.809 4.268 99.841 4.332 ;
			RECT	99.977 4.268 100.009 4.332 ;
			RECT	100.145 4.268 100.177 4.332 ;
			RECT	100.313 4.268 100.345 4.332 ;
			RECT	100.481 4.268 100.513 4.332 ;
			RECT	100.649 4.268 100.681 4.332 ;
			RECT	100.817 4.268 100.849 4.332 ;
			RECT	100.985 4.268 101.017 4.332 ;
			RECT	101.153 4.268 101.185 4.332 ;
			RECT	101.321 4.268 101.353 4.332 ;
			RECT	101.489 4.268 101.521 4.332 ;
			RECT	101.657 4.268 101.689 4.332 ;
			RECT	101.825 4.268 101.857 4.332 ;
			RECT	101.993 4.268 102.025 4.332 ;
			RECT	102.123 4.284 102.155 4.316 ;
			RECT	102.245 4.289 102.277 4.321 ;
			RECT	102.375 4.268 102.407 4.332 ;
			RECT	103.795 4.268 103.827 4.332 ;
			RECT	103.925 4.289 103.957 4.321 ;
			RECT	104.047 4.284 104.079 4.316 ;
			RECT	104.177 4.268 104.209 4.332 ;
			RECT	104.345 4.268 104.377 4.332 ;
			RECT	104.513 4.268 104.545 4.332 ;
			RECT	104.681 4.268 104.713 4.332 ;
			RECT	104.849 4.268 104.881 4.332 ;
			RECT	105.017 4.268 105.049 4.332 ;
			RECT	105.185 4.268 105.217 4.332 ;
			RECT	105.353 4.268 105.385 4.332 ;
			RECT	105.521 4.268 105.553 4.332 ;
			RECT	105.689 4.268 105.721 4.332 ;
			RECT	105.857 4.268 105.889 4.332 ;
			RECT	106.025 4.268 106.057 4.332 ;
			RECT	106.193 4.268 106.225 4.332 ;
			RECT	106.361 4.268 106.393 4.332 ;
			RECT	106.529 4.268 106.561 4.332 ;
			RECT	106.697 4.268 106.729 4.332 ;
			RECT	106.865 4.268 106.897 4.332 ;
			RECT	107.033 4.268 107.065 4.332 ;
			RECT	107.201 4.268 107.233 4.332 ;
			RECT	107.369 4.268 107.401 4.332 ;
			RECT	107.537 4.268 107.569 4.332 ;
			RECT	107.705 4.268 107.737 4.332 ;
			RECT	107.873 4.268 107.905 4.332 ;
			RECT	108.041 4.268 108.073 4.332 ;
			RECT	108.209 4.268 108.241 4.332 ;
			RECT	108.377 4.268 108.409 4.332 ;
			RECT	108.545 4.268 108.577 4.332 ;
			RECT	108.713 4.268 108.745 4.332 ;
			RECT	108.881 4.268 108.913 4.332 ;
			RECT	109.049 4.268 109.081 4.332 ;
			RECT	109.217 4.268 109.249 4.332 ;
			RECT	109.385 4.268 109.417 4.332 ;
			RECT	109.553 4.268 109.585 4.332 ;
			RECT	109.721 4.268 109.753 4.332 ;
			RECT	109.889 4.268 109.921 4.332 ;
			RECT	110.057 4.268 110.089 4.332 ;
			RECT	110.225 4.268 110.257 4.332 ;
			RECT	110.393 4.268 110.425 4.332 ;
			RECT	110.561 4.268 110.593 4.332 ;
			RECT	110.729 4.268 110.761 4.332 ;
			RECT	110.897 4.268 110.929 4.332 ;
			RECT	111.065 4.268 111.097 4.332 ;
			RECT	111.233 4.268 111.265 4.332 ;
			RECT	111.401 4.268 111.433 4.332 ;
			RECT	111.569 4.268 111.601 4.332 ;
			RECT	111.737 4.268 111.769 4.332 ;
			RECT	111.905 4.268 111.937 4.332 ;
			RECT	112.073 4.268 112.105 4.332 ;
			RECT	112.241 4.268 112.273 4.332 ;
			RECT	112.409 4.268 112.441 4.332 ;
			RECT	112.577 4.268 112.609 4.332 ;
			RECT	112.745 4.268 112.777 4.332 ;
			RECT	112.913 4.268 112.945 4.332 ;
			RECT	113.081 4.268 113.113 4.332 ;
			RECT	113.249 4.268 113.281 4.332 ;
			RECT	113.417 4.268 113.449 4.332 ;
			RECT	113.585 4.268 113.617 4.332 ;
			RECT	113.753 4.268 113.785 4.332 ;
			RECT	113.921 4.268 113.953 4.332 ;
			RECT	114.089 4.268 114.121 4.332 ;
			RECT	114.257 4.268 114.289 4.332 ;
			RECT	114.425 4.268 114.457 4.332 ;
			RECT	114.593 4.268 114.625 4.332 ;
			RECT	114.761 4.268 114.793 4.332 ;
			RECT	114.929 4.268 114.961 4.332 ;
			RECT	115.097 4.268 115.129 4.332 ;
			RECT	115.265 4.268 115.297 4.332 ;
			RECT	115.433 4.268 115.465 4.332 ;
			RECT	115.601 4.268 115.633 4.332 ;
			RECT	115.769 4.268 115.801 4.332 ;
			RECT	115.937 4.268 115.969 4.332 ;
			RECT	116.105 4.268 116.137 4.332 ;
			RECT	116.273 4.268 116.305 4.332 ;
			RECT	116.441 4.268 116.473 4.332 ;
			RECT	116.609 4.268 116.641 4.332 ;
			RECT	116.777 4.268 116.809 4.332 ;
			RECT	116.945 4.268 116.977 4.332 ;
			RECT	117.113 4.268 117.145 4.332 ;
			RECT	117.281 4.268 117.313 4.332 ;
			RECT	117.449 4.268 117.481 4.332 ;
			RECT	117.617 4.268 117.649 4.332 ;
			RECT	117.785 4.268 117.817 4.332 ;
			RECT	117.953 4.268 117.985 4.332 ;
			RECT	118.121 4.268 118.153 4.332 ;
			RECT	118.289 4.268 118.321 4.332 ;
			RECT	118.457 4.268 118.489 4.332 ;
			RECT	118.625 4.268 118.657 4.332 ;
			RECT	118.793 4.268 118.825 4.332 ;
			RECT	118.961 4.268 118.993 4.332 ;
			RECT	119.129 4.268 119.161 4.332 ;
			RECT	119.297 4.268 119.329 4.332 ;
			RECT	119.465 4.268 119.497 4.332 ;
			RECT	119.633 4.268 119.665 4.332 ;
			RECT	119.801 4.268 119.833 4.332 ;
			RECT	119.969 4.268 120.001 4.332 ;
			RECT	120.137 4.268 120.169 4.332 ;
			RECT	120.305 4.268 120.337 4.332 ;
			RECT	120.473 4.268 120.505 4.332 ;
			RECT	120.641 4.268 120.673 4.332 ;
			RECT	120.809 4.268 120.841 4.332 ;
			RECT	120.977 4.268 121.009 4.332 ;
			RECT	121.145 4.268 121.177 4.332 ;
			RECT	121.313 4.268 121.345 4.332 ;
			RECT	121.481 4.268 121.513 4.332 ;
			RECT	121.649 4.268 121.681 4.332 ;
			RECT	121.817 4.268 121.849 4.332 ;
			RECT	121.985 4.268 122.017 4.332 ;
			RECT	122.153 4.268 122.185 4.332 ;
			RECT	122.321 4.268 122.353 4.332 ;
			RECT	122.489 4.268 122.521 4.332 ;
			RECT	122.657 4.268 122.689 4.332 ;
			RECT	122.825 4.268 122.857 4.332 ;
			RECT	122.993 4.268 123.025 4.332 ;
			RECT	123.161 4.268 123.193 4.332 ;
			RECT	123.329 4.268 123.361 4.332 ;
			RECT	123.497 4.268 123.529 4.332 ;
			RECT	123.665 4.268 123.697 4.332 ;
			RECT	123.833 4.268 123.865 4.332 ;
			RECT	124.001 4.268 124.033 4.332 ;
			RECT	124.169 4.268 124.201 4.332 ;
			RECT	124.337 4.268 124.369 4.332 ;
			RECT	124.505 4.268 124.537 4.332 ;
			RECT	124.673 4.268 124.705 4.332 ;
			RECT	124.841 4.268 124.873 4.332 ;
			RECT	125.009 4.268 125.041 4.332 ;
			RECT	125.177 4.268 125.209 4.332 ;
			RECT	125.345 4.268 125.377 4.332 ;
			RECT	125.513 4.268 125.545 4.332 ;
			RECT	125.681 4.268 125.713 4.332 ;
			RECT	125.849 4.268 125.881 4.332 ;
			RECT	126.017 4.268 126.049 4.332 ;
			RECT	126.185 4.268 126.217 4.332 ;
			RECT	126.353 4.268 126.385 4.332 ;
			RECT	126.521 4.268 126.553 4.332 ;
			RECT	126.689 4.268 126.721 4.332 ;
			RECT	126.857 4.268 126.889 4.332 ;
			RECT	127.025 4.268 127.057 4.332 ;
			RECT	127.193 4.268 127.225 4.332 ;
			RECT	127.361 4.268 127.393 4.332 ;
			RECT	127.529 4.268 127.561 4.332 ;
			RECT	127.697 4.268 127.729 4.332 ;
			RECT	127.865 4.268 127.897 4.332 ;
			RECT	128.033 4.268 128.065 4.332 ;
			RECT	128.201 4.268 128.233 4.332 ;
			RECT	128.369 4.268 128.401 4.332 ;
			RECT	128.537 4.268 128.569 4.332 ;
			RECT	128.705 4.268 128.737 4.332 ;
			RECT	128.873 4.268 128.905 4.332 ;
			RECT	129.041 4.268 129.073 4.332 ;
			RECT	129.209 4.268 129.241 4.332 ;
			RECT	129.377 4.268 129.409 4.332 ;
			RECT	129.545 4.268 129.577 4.332 ;
			RECT	129.713 4.268 129.745 4.332 ;
			RECT	129.881 4.268 129.913 4.332 ;
			RECT	130.049 4.268 130.081 4.332 ;
			RECT	130.217 4.268 130.249 4.332 ;
			RECT	130.385 4.268 130.417 4.332 ;
			RECT	130.553 4.268 130.585 4.332 ;
			RECT	130.721 4.268 130.753 4.332 ;
			RECT	130.889 4.268 130.921 4.332 ;
			RECT	131.057 4.268 131.089 4.332 ;
			RECT	131.225 4.268 131.257 4.332 ;
			RECT	131.393 4.268 131.425 4.332 ;
			RECT	131.561 4.268 131.593 4.332 ;
			RECT	131.729 4.268 131.761 4.332 ;
			RECT	131.897 4.268 131.929 4.332 ;
			RECT	132.065 4.268 132.097 4.332 ;
			RECT	132.233 4.268 132.265 4.332 ;
			RECT	132.401 4.268 132.433 4.332 ;
			RECT	132.569 4.268 132.601 4.332 ;
			RECT	132.737 4.268 132.769 4.332 ;
			RECT	132.905 4.268 132.937 4.332 ;
			RECT	133.073 4.268 133.105 4.332 ;
			RECT	133.241 4.268 133.273 4.332 ;
			RECT	133.409 4.268 133.441 4.332 ;
			RECT	133.577 4.268 133.609 4.332 ;
			RECT	133.745 4.268 133.777 4.332 ;
			RECT	133.913 4.268 133.945 4.332 ;
			RECT	134.081 4.268 134.113 4.332 ;
			RECT	134.249 4.268 134.281 4.332 ;
			RECT	134.417 4.268 134.449 4.332 ;
			RECT	134.585 4.268 134.617 4.332 ;
			RECT	134.753 4.268 134.785 4.332 ;
			RECT	134.921 4.268 134.953 4.332 ;
			RECT	135.089 4.268 135.121 4.332 ;
			RECT	135.257 4.268 135.289 4.332 ;
			RECT	135.425 4.268 135.457 4.332 ;
			RECT	135.593 4.268 135.625 4.332 ;
			RECT	135.761 4.268 135.793 4.332 ;
			RECT	135.929 4.268 135.961 4.332 ;
			RECT	136.097 4.268 136.129 4.332 ;
			RECT	136.265 4.268 136.297 4.332 ;
			RECT	136.433 4.268 136.465 4.332 ;
			RECT	136.601 4.268 136.633 4.332 ;
			RECT	136.769 4.268 136.801 4.332 ;
			RECT	136.937 4.268 136.969 4.332 ;
			RECT	137.105 4.268 137.137 4.332 ;
			RECT	137.273 4.268 137.305 4.332 ;
			RECT	137.441 4.268 137.473 4.332 ;
			RECT	137.609 4.268 137.641 4.332 ;
			RECT	137.777 4.268 137.809 4.332 ;
			RECT	137.945 4.268 137.977 4.332 ;
			RECT	138.113 4.268 138.145 4.332 ;
			RECT	138.281 4.268 138.313 4.332 ;
			RECT	138.449 4.268 138.481 4.332 ;
			RECT	138.617 4.268 138.649 4.332 ;
			RECT	138.785 4.268 138.817 4.332 ;
			RECT	138.953 4.268 138.985 4.332 ;
			RECT	139.121 4.268 139.153 4.332 ;
			RECT	139.289 4.268 139.321 4.332 ;
			RECT	139.457 4.268 139.489 4.332 ;
			RECT	139.625 4.268 139.657 4.332 ;
			RECT	139.793 4.268 139.825 4.332 ;
			RECT	139.961 4.268 139.993 4.332 ;
			RECT	140.129 4.268 140.161 4.332 ;
			RECT	140.297 4.268 140.329 4.332 ;
			RECT	140.465 4.268 140.497 4.332 ;
			RECT	140.633 4.268 140.665 4.332 ;
			RECT	140.801 4.268 140.833 4.332 ;
			RECT	140.969 4.268 141.001 4.332 ;
			RECT	141.137 4.268 141.169 4.332 ;
			RECT	141.305 4.268 141.337 4.332 ;
			RECT	141.473 4.268 141.505 4.332 ;
			RECT	141.641 4.268 141.673 4.332 ;
			RECT	141.809 4.268 141.841 4.332 ;
			RECT	141.977 4.268 142.009 4.332 ;
			RECT	142.145 4.268 142.177 4.332 ;
			RECT	142.313 4.268 142.345 4.332 ;
			RECT	142.481 4.268 142.513 4.332 ;
			RECT	142.649 4.268 142.681 4.332 ;
			RECT	142.817 4.268 142.849 4.332 ;
			RECT	142.985 4.268 143.017 4.332 ;
			RECT	143.153 4.268 143.185 4.332 ;
			RECT	143.321 4.268 143.353 4.332 ;
			RECT	143.489 4.268 143.521 4.332 ;
			RECT	143.657 4.268 143.689 4.332 ;
			RECT	143.825 4.268 143.857 4.332 ;
			RECT	143.993 4.268 144.025 4.332 ;
			RECT	144.161 4.268 144.193 4.332 ;
			RECT	144.329 4.268 144.361 4.332 ;
			RECT	144.497 4.268 144.529 4.332 ;
			RECT	144.665 4.268 144.697 4.332 ;
			RECT	144.833 4.268 144.865 4.332 ;
			RECT	145.001 4.268 145.033 4.332 ;
			RECT	145.169 4.268 145.201 4.332 ;
			RECT	145.337 4.268 145.369 4.332 ;
			RECT	145.505 4.268 145.537 4.332 ;
			RECT	145.673 4.268 145.705 4.332 ;
			RECT	145.841 4.268 145.873 4.332 ;
			RECT	146.009 4.268 146.041 4.332 ;
			RECT	146.177 4.268 146.209 4.332 ;
			RECT	146.345 4.268 146.377 4.332 ;
			RECT	146.513 4.268 146.545 4.332 ;
			RECT	146.681 4.268 146.713 4.332 ;
			RECT	146.849 4.268 146.881 4.332 ;
			RECT	147.017 4.268 147.049 4.332 ;
			RECT	147.185 4.268 147.217 4.332 ;
			RECT	147.316 4.284 147.348 4.316 ;
			RECT	147.437 4.284 147.469 4.316 ;
			RECT	147.567 4.268 147.599 4.332 ;
			RECT	149.879 4.268 149.911 4.332 ;
			RECT	151.13 4.268 151.194 4.332 ;
			RECT	151.81 4.268 151.842 4.332 ;
			RECT	152.249 4.268 152.281 4.332 ;
			RECT	153.56 4.268 153.624 4.332 ;
			RECT	156.601 4.268 156.633 4.332 ;
			RECT	156.731 4.284 156.763 4.316 ;
			RECT	156.852 4.284 156.884 4.316 ;
			RECT	156.983 4.268 157.015 4.332 ;
			RECT	157.151 4.268 157.183 4.332 ;
			RECT	157.319 4.268 157.351 4.332 ;
			RECT	157.487 4.268 157.519 4.332 ;
			RECT	157.655 4.268 157.687 4.332 ;
			RECT	157.823 4.268 157.855 4.332 ;
			RECT	157.991 4.268 158.023 4.332 ;
			RECT	158.159 4.268 158.191 4.332 ;
			RECT	158.327 4.268 158.359 4.332 ;
			RECT	158.495 4.268 158.527 4.332 ;
			RECT	158.663 4.268 158.695 4.332 ;
			RECT	158.831 4.268 158.863 4.332 ;
			RECT	158.999 4.268 159.031 4.332 ;
			RECT	159.167 4.268 159.199 4.332 ;
			RECT	159.335 4.268 159.367 4.332 ;
			RECT	159.503 4.268 159.535 4.332 ;
			RECT	159.671 4.268 159.703 4.332 ;
			RECT	159.839 4.268 159.871 4.332 ;
			RECT	160.007 4.268 160.039 4.332 ;
			RECT	160.175 4.268 160.207 4.332 ;
			RECT	160.343 4.268 160.375 4.332 ;
			RECT	160.511 4.268 160.543 4.332 ;
			RECT	160.679 4.268 160.711 4.332 ;
			RECT	160.847 4.268 160.879 4.332 ;
			RECT	161.015 4.268 161.047 4.332 ;
			RECT	161.183 4.268 161.215 4.332 ;
			RECT	161.351 4.268 161.383 4.332 ;
			RECT	161.519 4.268 161.551 4.332 ;
			RECT	161.687 4.268 161.719 4.332 ;
			RECT	161.855 4.268 161.887 4.332 ;
			RECT	162.023 4.268 162.055 4.332 ;
			RECT	162.191 4.268 162.223 4.332 ;
			RECT	162.359 4.268 162.391 4.332 ;
			RECT	162.527 4.268 162.559 4.332 ;
			RECT	162.695 4.268 162.727 4.332 ;
			RECT	162.863 4.268 162.895 4.332 ;
			RECT	163.031 4.268 163.063 4.332 ;
			RECT	163.199 4.268 163.231 4.332 ;
			RECT	163.367 4.268 163.399 4.332 ;
			RECT	163.535 4.268 163.567 4.332 ;
			RECT	163.703 4.268 163.735 4.332 ;
			RECT	163.871 4.268 163.903 4.332 ;
			RECT	164.039 4.268 164.071 4.332 ;
			RECT	164.207 4.268 164.239 4.332 ;
			RECT	164.375 4.268 164.407 4.332 ;
			RECT	164.543 4.268 164.575 4.332 ;
			RECT	164.711 4.268 164.743 4.332 ;
			RECT	164.879 4.268 164.911 4.332 ;
			RECT	165.047 4.268 165.079 4.332 ;
			RECT	165.215 4.268 165.247 4.332 ;
			RECT	165.383 4.268 165.415 4.332 ;
			RECT	165.551 4.268 165.583 4.332 ;
			RECT	165.719 4.268 165.751 4.332 ;
			RECT	165.887 4.268 165.919 4.332 ;
			RECT	166.055 4.268 166.087 4.332 ;
			RECT	166.223 4.268 166.255 4.332 ;
			RECT	166.391 4.268 166.423 4.332 ;
			RECT	166.559 4.268 166.591 4.332 ;
			RECT	166.727 4.268 166.759 4.332 ;
			RECT	166.895 4.268 166.927 4.332 ;
			RECT	167.063 4.268 167.095 4.332 ;
			RECT	167.231 4.268 167.263 4.332 ;
			RECT	167.399 4.268 167.431 4.332 ;
			RECT	167.567 4.268 167.599 4.332 ;
			RECT	167.735 4.268 167.767 4.332 ;
			RECT	167.903 4.268 167.935 4.332 ;
			RECT	168.071 4.268 168.103 4.332 ;
			RECT	168.239 4.268 168.271 4.332 ;
			RECT	168.407 4.268 168.439 4.332 ;
			RECT	168.575 4.268 168.607 4.332 ;
			RECT	168.743 4.268 168.775 4.332 ;
			RECT	168.911 4.268 168.943 4.332 ;
			RECT	169.079 4.268 169.111 4.332 ;
			RECT	169.247 4.268 169.279 4.332 ;
			RECT	169.415 4.268 169.447 4.332 ;
			RECT	169.583 4.268 169.615 4.332 ;
			RECT	169.751 4.268 169.783 4.332 ;
			RECT	169.919 4.268 169.951 4.332 ;
			RECT	170.087 4.268 170.119 4.332 ;
			RECT	170.255 4.268 170.287 4.332 ;
			RECT	170.423 4.268 170.455 4.332 ;
			RECT	170.591 4.268 170.623 4.332 ;
			RECT	170.759 4.268 170.791 4.332 ;
			RECT	170.927 4.268 170.959 4.332 ;
			RECT	171.095 4.268 171.127 4.332 ;
			RECT	171.263 4.268 171.295 4.332 ;
			RECT	171.431 4.268 171.463 4.332 ;
			RECT	171.599 4.268 171.631 4.332 ;
			RECT	171.767 4.268 171.799 4.332 ;
			RECT	171.935 4.268 171.967 4.332 ;
			RECT	172.103 4.268 172.135 4.332 ;
			RECT	172.271 4.268 172.303 4.332 ;
			RECT	172.439 4.268 172.471 4.332 ;
			RECT	172.607 4.268 172.639 4.332 ;
			RECT	172.775 4.268 172.807 4.332 ;
			RECT	172.943 4.268 172.975 4.332 ;
			RECT	173.111 4.268 173.143 4.332 ;
			RECT	173.279 4.268 173.311 4.332 ;
			RECT	173.447 4.268 173.479 4.332 ;
			RECT	173.615 4.268 173.647 4.332 ;
			RECT	173.783 4.268 173.815 4.332 ;
			RECT	173.951 4.268 173.983 4.332 ;
			RECT	174.119 4.268 174.151 4.332 ;
			RECT	174.287 4.268 174.319 4.332 ;
			RECT	174.455 4.268 174.487 4.332 ;
			RECT	174.623 4.268 174.655 4.332 ;
			RECT	174.791 4.268 174.823 4.332 ;
			RECT	174.959 4.268 174.991 4.332 ;
			RECT	175.127 4.268 175.159 4.332 ;
			RECT	175.295 4.268 175.327 4.332 ;
			RECT	175.463 4.268 175.495 4.332 ;
			RECT	175.631 4.268 175.663 4.332 ;
			RECT	175.799 4.268 175.831 4.332 ;
			RECT	175.967 4.268 175.999 4.332 ;
			RECT	176.135 4.268 176.167 4.332 ;
			RECT	176.303 4.268 176.335 4.332 ;
			RECT	176.471 4.268 176.503 4.332 ;
			RECT	176.639 4.268 176.671 4.332 ;
			RECT	176.807 4.268 176.839 4.332 ;
			RECT	176.975 4.268 177.007 4.332 ;
			RECT	177.143 4.268 177.175 4.332 ;
			RECT	177.311 4.268 177.343 4.332 ;
			RECT	177.479 4.268 177.511 4.332 ;
			RECT	177.647 4.268 177.679 4.332 ;
			RECT	177.815 4.268 177.847 4.332 ;
			RECT	177.983 4.268 178.015 4.332 ;
			RECT	178.151 4.268 178.183 4.332 ;
			RECT	178.319 4.268 178.351 4.332 ;
			RECT	178.487 4.268 178.519 4.332 ;
			RECT	178.655 4.268 178.687 4.332 ;
			RECT	178.823 4.268 178.855 4.332 ;
			RECT	178.991 4.268 179.023 4.332 ;
			RECT	179.159 4.268 179.191 4.332 ;
			RECT	179.327 4.268 179.359 4.332 ;
			RECT	179.495 4.268 179.527 4.332 ;
			RECT	179.663 4.268 179.695 4.332 ;
			RECT	179.831 4.268 179.863 4.332 ;
			RECT	179.999 4.268 180.031 4.332 ;
			RECT	180.167 4.268 180.199 4.332 ;
			RECT	180.335 4.268 180.367 4.332 ;
			RECT	180.503 4.268 180.535 4.332 ;
			RECT	180.671 4.268 180.703 4.332 ;
			RECT	180.839 4.268 180.871 4.332 ;
			RECT	181.007 4.268 181.039 4.332 ;
			RECT	181.175 4.268 181.207 4.332 ;
			RECT	181.343 4.268 181.375 4.332 ;
			RECT	181.511 4.268 181.543 4.332 ;
			RECT	181.679 4.268 181.711 4.332 ;
			RECT	181.847 4.268 181.879 4.332 ;
			RECT	182.015 4.268 182.047 4.332 ;
			RECT	182.183 4.268 182.215 4.332 ;
			RECT	182.351 4.268 182.383 4.332 ;
			RECT	182.519 4.268 182.551 4.332 ;
			RECT	182.687 4.268 182.719 4.332 ;
			RECT	182.855 4.268 182.887 4.332 ;
			RECT	183.023 4.268 183.055 4.332 ;
			RECT	183.191 4.268 183.223 4.332 ;
			RECT	183.359 4.268 183.391 4.332 ;
			RECT	183.527 4.268 183.559 4.332 ;
			RECT	183.695 4.268 183.727 4.332 ;
			RECT	183.863 4.268 183.895 4.332 ;
			RECT	184.031 4.268 184.063 4.332 ;
			RECT	184.199 4.268 184.231 4.332 ;
			RECT	184.367 4.268 184.399 4.332 ;
			RECT	184.535 4.268 184.567 4.332 ;
			RECT	184.703 4.268 184.735 4.332 ;
			RECT	184.871 4.268 184.903 4.332 ;
			RECT	185.039 4.268 185.071 4.332 ;
			RECT	185.207 4.268 185.239 4.332 ;
			RECT	185.375 4.268 185.407 4.332 ;
			RECT	185.543 4.268 185.575 4.332 ;
			RECT	185.711 4.268 185.743 4.332 ;
			RECT	185.879 4.268 185.911 4.332 ;
			RECT	186.047 4.268 186.079 4.332 ;
			RECT	186.215 4.268 186.247 4.332 ;
			RECT	186.383 4.268 186.415 4.332 ;
			RECT	186.551 4.268 186.583 4.332 ;
			RECT	186.719 4.268 186.751 4.332 ;
			RECT	186.887 4.268 186.919 4.332 ;
			RECT	187.055 4.268 187.087 4.332 ;
			RECT	187.223 4.268 187.255 4.332 ;
			RECT	187.391 4.268 187.423 4.332 ;
			RECT	187.559 4.268 187.591 4.332 ;
			RECT	187.727 4.268 187.759 4.332 ;
			RECT	187.895 4.268 187.927 4.332 ;
			RECT	188.063 4.268 188.095 4.332 ;
			RECT	188.231 4.268 188.263 4.332 ;
			RECT	188.399 4.268 188.431 4.332 ;
			RECT	188.567 4.268 188.599 4.332 ;
			RECT	188.735 4.268 188.767 4.332 ;
			RECT	188.903 4.268 188.935 4.332 ;
			RECT	189.071 4.268 189.103 4.332 ;
			RECT	189.239 4.268 189.271 4.332 ;
			RECT	189.407 4.268 189.439 4.332 ;
			RECT	189.575 4.268 189.607 4.332 ;
			RECT	189.743 4.268 189.775 4.332 ;
			RECT	189.911 4.268 189.943 4.332 ;
			RECT	190.079 4.268 190.111 4.332 ;
			RECT	190.247 4.268 190.279 4.332 ;
			RECT	190.415 4.268 190.447 4.332 ;
			RECT	190.583 4.268 190.615 4.332 ;
			RECT	190.751 4.268 190.783 4.332 ;
			RECT	190.919 4.268 190.951 4.332 ;
			RECT	191.087 4.268 191.119 4.332 ;
			RECT	191.255 4.268 191.287 4.332 ;
			RECT	191.423 4.268 191.455 4.332 ;
			RECT	191.591 4.268 191.623 4.332 ;
			RECT	191.759 4.268 191.791 4.332 ;
			RECT	191.927 4.268 191.959 4.332 ;
			RECT	192.095 4.268 192.127 4.332 ;
			RECT	192.263 4.268 192.295 4.332 ;
			RECT	192.431 4.268 192.463 4.332 ;
			RECT	192.599 4.268 192.631 4.332 ;
			RECT	192.767 4.268 192.799 4.332 ;
			RECT	192.935 4.268 192.967 4.332 ;
			RECT	193.103 4.268 193.135 4.332 ;
			RECT	193.271 4.268 193.303 4.332 ;
			RECT	193.439 4.268 193.471 4.332 ;
			RECT	193.607 4.268 193.639 4.332 ;
			RECT	193.775 4.268 193.807 4.332 ;
			RECT	193.943 4.268 193.975 4.332 ;
			RECT	194.111 4.268 194.143 4.332 ;
			RECT	194.279 4.268 194.311 4.332 ;
			RECT	194.447 4.268 194.479 4.332 ;
			RECT	194.615 4.268 194.647 4.332 ;
			RECT	194.783 4.268 194.815 4.332 ;
			RECT	194.951 4.268 194.983 4.332 ;
			RECT	195.119 4.268 195.151 4.332 ;
			RECT	195.287 4.268 195.319 4.332 ;
			RECT	195.455 4.268 195.487 4.332 ;
			RECT	195.623 4.268 195.655 4.332 ;
			RECT	195.791 4.268 195.823 4.332 ;
			RECT	195.959 4.268 195.991 4.332 ;
			RECT	196.127 4.268 196.159 4.332 ;
			RECT	196.295 4.268 196.327 4.332 ;
			RECT	196.463 4.268 196.495 4.332 ;
			RECT	196.631 4.268 196.663 4.332 ;
			RECT	196.799 4.268 196.831 4.332 ;
			RECT	196.967 4.268 196.999 4.332 ;
			RECT	197.135 4.268 197.167 4.332 ;
			RECT	197.303 4.268 197.335 4.332 ;
			RECT	197.471 4.268 197.503 4.332 ;
			RECT	197.639 4.268 197.671 4.332 ;
			RECT	197.807 4.268 197.839 4.332 ;
			RECT	197.975 4.268 198.007 4.332 ;
			RECT	198.143 4.268 198.175 4.332 ;
			RECT	198.311 4.268 198.343 4.332 ;
			RECT	198.479 4.268 198.511 4.332 ;
			RECT	198.647 4.268 198.679 4.332 ;
			RECT	198.815 4.268 198.847 4.332 ;
			RECT	198.983 4.268 199.015 4.332 ;
			RECT	199.151 4.268 199.183 4.332 ;
			RECT	199.319 4.268 199.351 4.332 ;
			RECT	199.487 4.268 199.519 4.332 ;
			RECT	199.655 4.268 199.687 4.332 ;
			RECT	199.823 4.268 199.855 4.332 ;
			RECT	199.991 4.268 200.023 4.332 ;
			RECT	200.121 4.284 200.153 4.316 ;
			RECT	200.243 4.289 200.275 4.321 ;
			RECT	200.373 4.268 200.405 4.332 ;
			RECT	200.9 4.268 200.932 4.332 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 2.32 201.665 2.44 ;
			LAYER	J3 ;
			RECT	0.755 2.348 0.787 2.412 ;
			RECT	1.645 2.348 1.709 2.412 ;
			RECT	2.323 2.348 2.387 2.412 ;
			RECT	3.438 2.348 3.47 2.412 ;
			RECT	3.585 2.348 3.617 2.412 ;
			RECT	4.195 2.348 4.227 2.412 ;
			RECT	4.72 2.348 4.752 2.412 ;
			RECT	4.944 2.348 5.008 2.412 ;
			RECT	5.267 2.348 5.299 2.412 ;
			RECT	5.797 2.348 5.829 2.412 ;
			RECT	5.927 2.369 5.959 2.401 ;
			RECT	6.049 2.364 6.081 2.396 ;
			RECT	6.179 2.348 6.211 2.412 ;
			RECT	6.347 2.348 6.379 2.412 ;
			RECT	6.515 2.348 6.547 2.412 ;
			RECT	6.683 2.348 6.715 2.412 ;
			RECT	6.851 2.348 6.883 2.412 ;
			RECT	7.019 2.348 7.051 2.412 ;
			RECT	7.187 2.348 7.219 2.412 ;
			RECT	7.355 2.348 7.387 2.412 ;
			RECT	7.523 2.348 7.555 2.412 ;
			RECT	7.691 2.348 7.723 2.412 ;
			RECT	7.859 2.348 7.891 2.412 ;
			RECT	8.027 2.348 8.059 2.412 ;
			RECT	8.195 2.348 8.227 2.412 ;
			RECT	8.363 2.348 8.395 2.412 ;
			RECT	8.531 2.348 8.563 2.412 ;
			RECT	8.699 2.348 8.731 2.412 ;
			RECT	8.867 2.348 8.899 2.412 ;
			RECT	9.035 2.348 9.067 2.412 ;
			RECT	9.203 2.348 9.235 2.412 ;
			RECT	9.371 2.348 9.403 2.412 ;
			RECT	9.539 2.348 9.571 2.412 ;
			RECT	9.707 2.348 9.739 2.412 ;
			RECT	9.875 2.348 9.907 2.412 ;
			RECT	10.043 2.348 10.075 2.412 ;
			RECT	10.211 2.348 10.243 2.412 ;
			RECT	10.379 2.348 10.411 2.412 ;
			RECT	10.547 2.348 10.579 2.412 ;
			RECT	10.715 2.348 10.747 2.412 ;
			RECT	10.883 2.348 10.915 2.412 ;
			RECT	11.051 2.348 11.083 2.412 ;
			RECT	11.219 2.348 11.251 2.412 ;
			RECT	11.387 2.348 11.419 2.412 ;
			RECT	11.555 2.348 11.587 2.412 ;
			RECT	11.723 2.348 11.755 2.412 ;
			RECT	11.891 2.348 11.923 2.412 ;
			RECT	12.059 2.348 12.091 2.412 ;
			RECT	12.227 2.348 12.259 2.412 ;
			RECT	12.395 2.348 12.427 2.412 ;
			RECT	12.563 2.348 12.595 2.412 ;
			RECT	12.731 2.348 12.763 2.412 ;
			RECT	12.899 2.348 12.931 2.412 ;
			RECT	13.067 2.348 13.099 2.412 ;
			RECT	13.235 2.348 13.267 2.412 ;
			RECT	13.403 2.348 13.435 2.412 ;
			RECT	13.571 2.348 13.603 2.412 ;
			RECT	13.739 2.348 13.771 2.412 ;
			RECT	13.907 2.348 13.939 2.412 ;
			RECT	14.075 2.348 14.107 2.412 ;
			RECT	14.243 2.348 14.275 2.412 ;
			RECT	14.411 2.348 14.443 2.412 ;
			RECT	14.579 2.348 14.611 2.412 ;
			RECT	14.747 2.348 14.779 2.412 ;
			RECT	14.915 2.348 14.947 2.412 ;
			RECT	15.083 2.348 15.115 2.412 ;
			RECT	15.251 2.348 15.283 2.412 ;
			RECT	15.419 2.348 15.451 2.412 ;
			RECT	15.587 2.348 15.619 2.412 ;
			RECT	15.755 2.348 15.787 2.412 ;
			RECT	15.923 2.348 15.955 2.412 ;
			RECT	16.091 2.348 16.123 2.412 ;
			RECT	16.259 2.348 16.291 2.412 ;
			RECT	16.427 2.348 16.459 2.412 ;
			RECT	16.595 2.348 16.627 2.412 ;
			RECT	16.763 2.348 16.795 2.412 ;
			RECT	16.931 2.348 16.963 2.412 ;
			RECT	17.099 2.348 17.131 2.412 ;
			RECT	17.267 2.348 17.299 2.412 ;
			RECT	17.435 2.348 17.467 2.412 ;
			RECT	17.603 2.348 17.635 2.412 ;
			RECT	17.771 2.348 17.803 2.412 ;
			RECT	17.939 2.348 17.971 2.412 ;
			RECT	18.107 2.348 18.139 2.412 ;
			RECT	18.275 2.348 18.307 2.412 ;
			RECT	18.443 2.348 18.475 2.412 ;
			RECT	18.611 2.348 18.643 2.412 ;
			RECT	18.779 2.348 18.811 2.412 ;
			RECT	18.947 2.348 18.979 2.412 ;
			RECT	19.115 2.348 19.147 2.412 ;
			RECT	19.283 2.348 19.315 2.412 ;
			RECT	19.451 2.348 19.483 2.412 ;
			RECT	19.619 2.348 19.651 2.412 ;
			RECT	19.787 2.348 19.819 2.412 ;
			RECT	19.955 2.348 19.987 2.412 ;
			RECT	20.123 2.348 20.155 2.412 ;
			RECT	20.291 2.348 20.323 2.412 ;
			RECT	20.459 2.348 20.491 2.412 ;
			RECT	20.627 2.348 20.659 2.412 ;
			RECT	20.795 2.348 20.827 2.412 ;
			RECT	20.963 2.348 20.995 2.412 ;
			RECT	21.131 2.348 21.163 2.412 ;
			RECT	21.299 2.348 21.331 2.412 ;
			RECT	21.467 2.348 21.499 2.412 ;
			RECT	21.635 2.348 21.667 2.412 ;
			RECT	21.803 2.348 21.835 2.412 ;
			RECT	21.971 2.348 22.003 2.412 ;
			RECT	22.139 2.348 22.171 2.412 ;
			RECT	22.307 2.348 22.339 2.412 ;
			RECT	22.475 2.348 22.507 2.412 ;
			RECT	22.643 2.348 22.675 2.412 ;
			RECT	22.811 2.348 22.843 2.412 ;
			RECT	22.979 2.348 23.011 2.412 ;
			RECT	23.147 2.348 23.179 2.412 ;
			RECT	23.315 2.348 23.347 2.412 ;
			RECT	23.483 2.348 23.515 2.412 ;
			RECT	23.651 2.348 23.683 2.412 ;
			RECT	23.819 2.348 23.851 2.412 ;
			RECT	23.987 2.348 24.019 2.412 ;
			RECT	24.155 2.348 24.187 2.412 ;
			RECT	24.323 2.348 24.355 2.412 ;
			RECT	24.491 2.348 24.523 2.412 ;
			RECT	24.659 2.348 24.691 2.412 ;
			RECT	24.827 2.348 24.859 2.412 ;
			RECT	24.995 2.348 25.027 2.412 ;
			RECT	25.163 2.348 25.195 2.412 ;
			RECT	25.331 2.348 25.363 2.412 ;
			RECT	25.499 2.348 25.531 2.412 ;
			RECT	25.667 2.348 25.699 2.412 ;
			RECT	25.835 2.348 25.867 2.412 ;
			RECT	26.003 2.348 26.035 2.412 ;
			RECT	26.171 2.348 26.203 2.412 ;
			RECT	26.339 2.348 26.371 2.412 ;
			RECT	26.507 2.348 26.539 2.412 ;
			RECT	26.675 2.348 26.707 2.412 ;
			RECT	26.843 2.348 26.875 2.412 ;
			RECT	27.011 2.348 27.043 2.412 ;
			RECT	27.179 2.348 27.211 2.412 ;
			RECT	27.347 2.348 27.379 2.412 ;
			RECT	27.515 2.348 27.547 2.412 ;
			RECT	27.683 2.348 27.715 2.412 ;
			RECT	27.851 2.348 27.883 2.412 ;
			RECT	28.019 2.348 28.051 2.412 ;
			RECT	28.187 2.348 28.219 2.412 ;
			RECT	28.355 2.348 28.387 2.412 ;
			RECT	28.523 2.348 28.555 2.412 ;
			RECT	28.691 2.348 28.723 2.412 ;
			RECT	28.859 2.348 28.891 2.412 ;
			RECT	29.027 2.348 29.059 2.412 ;
			RECT	29.195 2.348 29.227 2.412 ;
			RECT	29.363 2.348 29.395 2.412 ;
			RECT	29.531 2.348 29.563 2.412 ;
			RECT	29.699 2.348 29.731 2.412 ;
			RECT	29.867 2.348 29.899 2.412 ;
			RECT	30.035 2.348 30.067 2.412 ;
			RECT	30.203 2.348 30.235 2.412 ;
			RECT	30.371 2.348 30.403 2.412 ;
			RECT	30.539 2.348 30.571 2.412 ;
			RECT	30.707 2.348 30.739 2.412 ;
			RECT	30.875 2.348 30.907 2.412 ;
			RECT	31.043 2.348 31.075 2.412 ;
			RECT	31.211 2.348 31.243 2.412 ;
			RECT	31.379 2.348 31.411 2.412 ;
			RECT	31.547 2.348 31.579 2.412 ;
			RECT	31.715 2.348 31.747 2.412 ;
			RECT	31.883 2.348 31.915 2.412 ;
			RECT	32.051 2.348 32.083 2.412 ;
			RECT	32.219 2.348 32.251 2.412 ;
			RECT	32.387 2.348 32.419 2.412 ;
			RECT	32.555 2.348 32.587 2.412 ;
			RECT	32.723 2.348 32.755 2.412 ;
			RECT	32.891 2.348 32.923 2.412 ;
			RECT	33.059 2.348 33.091 2.412 ;
			RECT	33.227 2.348 33.259 2.412 ;
			RECT	33.395 2.348 33.427 2.412 ;
			RECT	33.563 2.348 33.595 2.412 ;
			RECT	33.731 2.348 33.763 2.412 ;
			RECT	33.899 2.348 33.931 2.412 ;
			RECT	34.067 2.348 34.099 2.412 ;
			RECT	34.235 2.348 34.267 2.412 ;
			RECT	34.403 2.348 34.435 2.412 ;
			RECT	34.571 2.348 34.603 2.412 ;
			RECT	34.739 2.348 34.771 2.412 ;
			RECT	34.907 2.348 34.939 2.412 ;
			RECT	35.075 2.348 35.107 2.412 ;
			RECT	35.243 2.348 35.275 2.412 ;
			RECT	35.411 2.348 35.443 2.412 ;
			RECT	35.579 2.348 35.611 2.412 ;
			RECT	35.747 2.348 35.779 2.412 ;
			RECT	35.915 2.348 35.947 2.412 ;
			RECT	36.083 2.348 36.115 2.412 ;
			RECT	36.251 2.348 36.283 2.412 ;
			RECT	36.419 2.348 36.451 2.412 ;
			RECT	36.587 2.348 36.619 2.412 ;
			RECT	36.755 2.348 36.787 2.412 ;
			RECT	36.923 2.348 36.955 2.412 ;
			RECT	37.091 2.348 37.123 2.412 ;
			RECT	37.259 2.348 37.291 2.412 ;
			RECT	37.427 2.348 37.459 2.412 ;
			RECT	37.595 2.348 37.627 2.412 ;
			RECT	37.763 2.348 37.795 2.412 ;
			RECT	37.931 2.348 37.963 2.412 ;
			RECT	38.099 2.348 38.131 2.412 ;
			RECT	38.267 2.348 38.299 2.412 ;
			RECT	38.435 2.348 38.467 2.412 ;
			RECT	38.603 2.348 38.635 2.412 ;
			RECT	38.771 2.348 38.803 2.412 ;
			RECT	38.939 2.348 38.971 2.412 ;
			RECT	39.107 2.348 39.139 2.412 ;
			RECT	39.275 2.348 39.307 2.412 ;
			RECT	39.443 2.348 39.475 2.412 ;
			RECT	39.611 2.348 39.643 2.412 ;
			RECT	39.779 2.348 39.811 2.412 ;
			RECT	39.947 2.348 39.979 2.412 ;
			RECT	40.115 2.348 40.147 2.412 ;
			RECT	40.283 2.348 40.315 2.412 ;
			RECT	40.451 2.348 40.483 2.412 ;
			RECT	40.619 2.348 40.651 2.412 ;
			RECT	40.787 2.348 40.819 2.412 ;
			RECT	40.955 2.348 40.987 2.412 ;
			RECT	41.123 2.348 41.155 2.412 ;
			RECT	41.291 2.348 41.323 2.412 ;
			RECT	41.459 2.348 41.491 2.412 ;
			RECT	41.627 2.348 41.659 2.412 ;
			RECT	41.795 2.348 41.827 2.412 ;
			RECT	41.963 2.348 41.995 2.412 ;
			RECT	42.131 2.348 42.163 2.412 ;
			RECT	42.299 2.348 42.331 2.412 ;
			RECT	42.467 2.348 42.499 2.412 ;
			RECT	42.635 2.348 42.667 2.412 ;
			RECT	42.803 2.348 42.835 2.412 ;
			RECT	42.971 2.348 43.003 2.412 ;
			RECT	43.139 2.348 43.171 2.412 ;
			RECT	43.307 2.348 43.339 2.412 ;
			RECT	43.475 2.348 43.507 2.412 ;
			RECT	43.643 2.348 43.675 2.412 ;
			RECT	43.811 2.348 43.843 2.412 ;
			RECT	43.979 2.348 44.011 2.412 ;
			RECT	44.147 2.348 44.179 2.412 ;
			RECT	44.315 2.348 44.347 2.412 ;
			RECT	44.483 2.348 44.515 2.412 ;
			RECT	44.651 2.348 44.683 2.412 ;
			RECT	44.819 2.348 44.851 2.412 ;
			RECT	44.987 2.348 45.019 2.412 ;
			RECT	45.155 2.348 45.187 2.412 ;
			RECT	45.323 2.348 45.355 2.412 ;
			RECT	45.491 2.348 45.523 2.412 ;
			RECT	45.659 2.348 45.691 2.412 ;
			RECT	45.827 2.348 45.859 2.412 ;
			RECT	45.995 2.348 46.027 2.412 ;
			RECT	46.163 2.348 46.195 2.412 ;
			RECT	46.331 2.348 46.363 2.412 ;
			RECT	46.499 2.348 46.531 2.412 ;
			RECT	46.667 2.348 46.699 2.412 ;
			RECT	46.835 2.348 46.867 2.412 ;
			RECT	47.003 2.348 47.035 2.412 ;
			RECT	47.171 2.348 47.203 2.412 ;
			RECT	47.339 2.348 47.371 2.412 ;
			RECT	47.507 2.348 47.539 2.412 ;
			RECT	47.675 2.348 47.707 2.412 ;
			RECT	47.843 2.348 47.875 2.412 ;
			RECT	48.011 2.348 48.043 2.412 ;
			RECT	48.179 2.348 48.211 2.412 ;
			RECT	48.347 2.348 48.379 2.412 ;
			RECT	48.515 2.348 48.547 2.412 ;
			RECT	48.683 2.348 48.715 2.412 ;
			RECT	48.851 2.348 48.883 2.412 ;
			RECT	49.019 2.348 49.051 2.412 ;
			RECT	49.187 2.348 49.219 2.412 ;
			RECT	49.318 2.364 49.35 2.396 ;
			RECT	49.439 2.364 49.471 2.396 ;
			RECT	49.569 2.348 49.601 2.412 ;
			RECT	51.881 2.348 51.913 2.412 ;
			RECT	53.132 2.348 53.196 2.412 ;
			RECT	53.812 2.348 53.844 2.412 ;
			RECT	54.251 2.348 54.283 2.412 ;
			RECT	55.562 2.348 55.626 2.412 ;
			RECT	58.603 2.348 58.635 2.412 ;
			RECT	58.733 2.364 58.765 2.396 ;
			RECT	58.854 2.364 58.886 2.396 ;
			RECT	58.985 2.348 59.017 2.412 ;
			RECT	59.153 2.348 59.185 2.412 ;
			RECT	59.321 2.348 59.353 2.412 ;
			RECT	59.489 2.348 59.521 2.412 ;
			RECT	59.657 2.348 59.689 2.412 ;
			RECT	59.825 2.348 59.857 2.412 ;
			RECT	59.993 2.348 60.025 2.412 ;
			RECT	60.161 2.348 60.193 2.412 ;
			RECT	60.329 2.348 60.361 2.412 ;
			RECT	60.497 2.348 60.529 2.412 ;
			RECT	60.665 2.348 60.697 2.412 ;
			RECT	60.833 2.348 60.865 2.412 ;
			RECT	61.001 2.348 61.033 2.412 ;
			RECT	61.169 2.348 61.201 2.412 ;
			RECT	61.337 2.348 61.369 2.412 ;
			RECT	61.505 2.348 61.537 2.412 ;
			RECT	61.673 2.348 61.705 2.412 ;
			RECT	61.841 2.348 61.873 2.412 ;
			RECT	62.009 2.348 62.041 2.412 ;
			RECT	62.177 2.348 62.209 2.412 ;
			RECT	62.345 2.348 62.377 2.412 ;
			RECT	62.513 2.348 62.545 2.412 ;
			RECT	62.681 2.348 62.713 2.412 ;
			RECT	62.849 2.348 62.881 2.412 ;
			RECT	63.017 2.348 63.049 2.412 ;
			RECT	63.185 2.348 63.217 2.412 ;
			RECT	63.353 2.348 63.385 2.412 ;
			RECT	63.521 2.348 63.553 2.412 ;
			RECT	63.689 2.348 63.721 2.412 ;
			RECT	63.857 2.348 63.889 2.412 ;
			RECT	64.025 2.348 64.057 2.412 ;
			RECT	64.193 2.348 64.225 2.412 ;
			RECT	64.361 2.348 64.393 2.412 ;
			RECT	64.529 2.348 64.561 2.412 ;
			RECT	64.697 2.348 64.729 2.412 ;
			RECT	64.865 2.348 64.897 2.412 ;
			RECT	65.033 2.348 65.065 2.412 ;
			RECT	65.201 2.348 65.233 2.412 ;
			RECT	65.369 2.348 65.401 2.412 ;
			RECT	65.537 2.348 65.569 2.412 ;
			RECT	65.705 2.348 65.737 2.412 ;
			RECT	65.873 2.348 65.905 2.412 ;
			RECT	66.041 2.348 66.073 2.412 ;
			RECT	66.209 2.348 66.241 2.412 ;
			RECT	66.377 2.348 66.409 2.412 ;
			RECT	66.545 2.348 66.577 2.412 ;
			RECT	66.713 2.348 66.745 2.412 ;
			RECT	66.881 2.348 66.913 2.412 ;
			RECT	67.049 2.348 67.081 2.412 ;
			RECT	67.217 2.348 67.249 2.412 ;
			RECT	67.385 2.348 67.417 2.412 ;
			RECT	67.553 2.348 67.585 2.412 ;
			RECT	67.721 2.348 67.753 2.412 ;
			RECT	67.889 2.348 67.921 2.412 ;
			RECT	68.057 2.348 68.089 2.412 ;
			RECT	68.225 2.348 68.257 2.412 ;
			RECT	68.393 2.348 68.425 2.412 ;
			RECT	68.561 2.348 68.593 2.412 ;
			RECT	68.729 2.348 68.761 2.412 ;
			RECT	68.897 2.348 68.929 2.412 ;
			RECT	69.065 2.348 69.097 2.412 ;
			RECT	69.233 2.348 69.265 2.412 ;
			RECT	69.401 2.348 69.433 2.412 ;
			RECT	69.569 2.348 69.601 2.412 ;
			RECT	69.737 2.348 69.769 2.412 ;
			RECT	69.905 2.348 69.937 2.412 ;
			RECT	70.073 2.348 70.105 2.412 ;
			RECT	70.241 2.348 70.273 2.412 ;
			RECT	70.409 2.348 70.441 2.412 ;
			RECT	70.577 2.348 70.609 2.412 ;
			RECT	70.745 2.348 70.777 2.412 ;
			RECT	70.913 2.348 70.945 2.412 ;
			RECT	71.081 2.348 71.113 2.412 ;
			RECT	71.249 2.348 71.281 2.412 ;
			RECT	71.417 2.348 71.449 2.412 ;
			RECT	71.585 2.348 71.617 2.412 ;
			RECT	71.753 2.348 71.785 2.412 ;
			RECT	71.921 2.348 71.953 2.412 ;
			RECT	72.089 2.348 72.121 2.412 ;
			RECT	72.257 2.348 72.289 2.412 ;
			RECT	72.425 2.348 72.457 2.412 ;
			RECT	72.593 2.348 72.625 2.412 ;
			RECT	72.761 2.348 72.793 2.412 ;
			RECT	72.929 2.348 72.961 2.412 ;
			RECT	73.097 2.348 73.129 2.412 ;
			RECT	73.265 2.348 73.297 2.412 ;
			RECT	73.433 2.348 73.465 2.412 ;
			RECT	73.601 2.348 73.633 2.412 ;
			RECT	73.769 2.348 73.801 2.412 ;
			RECT	73.937 2.348 73.969 2.412 ;
			RECT	74.105 2.348 74.137 2.412 ;
			RECT	74.273 2.348 74.305 2.412 ;
			RECT	74.441 2.348 74.473 2.412 ;
			RECT	74.609 2.348 74.641 2.412 ;
			RECT	74.777 2.348 74.809 2.412 ;
			RECT	74.945 2.348 74.977 2.412 ;
			RECT	75.113 2.348 75.145 2.412 ;
			RECT	75.281 2.348 75.313 2.412 ;
			RECT	75.449 2.348 75.481 2.412 ;
			RECT	75.617 2.348 75.649 2.412 ;
			RECT	75.785 2.348 75.817 2.412 ;
			RECT	75.953 2.348 75.985 2.412 ;
			RECT	76.121 2.348 76.153 2.412 ;
			RECT	76.289 2.348 76.321 2.412 ;
			RECT	76.457 2.348 76.489 2.412 ;
			RECT	76.625 2.348 76.657 2.412 ;
			RECT	76.793 2.348 76.825 2.412 ;
			RECT	76.961 2.348 76.993 2.412 ;
			RECT	77.129 2.348 77.161 2.412 ;
			RECT	77.297 2.348 77.329 2.412 ;
			RECT	77.465 2.348 77.497 2.412 ;
			RECT	77.633 2.348 77.665 2.412 ;
			RECT	77.801 2.348 77.833 2.412 ;
			RECT	77.969 2.348 78.001 2.412 ;
			RECT	78.137 2.348 78.169 2.412 ;
			RECT	78.305 2.348 78.337 2.412 ;
			RECT	78.473 2.348 78.505 2.412 ;
			RECT	78.641 2.348 78.673 2.412 ;
			RECT	78.809 2.348 78.841 2.412 ;
			RECT	78.977 2.348 79.009 2.412 ;
			RECT	79.145 2.348 79.177 2.412 ;
			RECT	79.313 2.348 79.345 2.412 ;
			RECT	79.481 2.348 79.513 2.412 ;
			RECT	79.649 2.348 79.681 2.412 ;
			RECT	79.817 2.348 79.849 2.412 ;
			RECT	79.985 2.348 80.017 2.412 ;
			RECT	80.153 2.348 80.185 2.412 ;
			RECT	80.321 2.348 80.353 2.412 ;
			RECT	80.489 2.348 80.521 2.412 ;
			RECT	80.657 2.348 80.689 2.412 ;
			RECT	80.825 2.348 80.857 2.412 ;
			RECT	80.993 2.348 81.025 2.412 ;
			RECT	81.161 2.348 81.193 2.412 ;
			RECT	81.329 2.348 81.361 2.412 ;
			RECT	81.497 2.348 81.529 2.412 ;
			RECT	81.665 2.348 81.697 2.412 ;
			RECT	81.833 2.348 81.865 2.412 ;
			RECT	82.001 2.348 82.033 2.412 ;
			RECT	82.169 2.348 82.201 2.412 ;
			RECT	82.337 2.348 82.369 2.412 ;
			RECT	82.505 2.348 82.537 2.412 ;
			RECT	82.673 2.348 82.705 2.412 ;
			RECT	82.841 2.348 82.873 2.412 ;
			RECT	83.009 2.348 83.041 2.412 ;
			RECT	83.177 2.348 83.209 2.412 ;
			RECT	83.345 2.348 83.377 2.412 ;
			RECT	83.513 2.348 83.545 2.412 ;
			RECT	83.681 2.348 83.713 2.412 ;
			RECT	83.849 2.348 83.881 2.412 ;
			RECT	84.017 2.348 84.049 2.412 ;
			RECT	84.185 2.348 84.217 2.412 ;
			RECT	84.353 2.348 84.385 2.412 ;
			RECT	84.521 2.348 84.553 2.412 ;
			RECT	84.689 2.348 84.721 2.412 ;
			RECT	84.857 2.348 84.889 2.412 ;
			RECT	85.025 2.348 85.057 2.412 ;
			RECT	85.193 2.348 85.225 2.412 ;
			RECT	85.361 2.348 85.393 2.412 ;
			RECT	85.529 2.348 85.561 2.412 ;
			RECT	85.697 2.348 85.729 2.412 ;
			RECT	85.865 2.348 85.897 2.412 ;
			RECT	86.033 2.348 86.065 2.412 ;
			RECT	86.201 2.348 86.233 2.412 ;
			RECT	86.369 2.348 86.401 2.412 ;
			RECT	86.537 2.348 86.569 2.412 ;
			RECT	86.705 2.348 86.737 2.412 ;
			RECT	86.873 2.348 86.905 2.412 ;
			RECT	87.041 2.348 87.073 2.412 ;
			RECT	87.209 2.348 87.241 2.412 ;
			RECT	87.377 2.348 87.409 2.412 ;
			RECT	87.545 2.348 87.577 2.412 ;
			RECT	87.713 2.348 87.745 2.412 ;
			RECT	87.881 2.348 87.913 2.412 ;
			RECT	88.049 2.348 88.081 2.412 ;
			RECT	88.217 2.348 88.249 2.412 ;
			RECT	88.385 2.348 88.417 2.412 ;
			RECT	88.553 2.348 88.585 2.412 ;
			RECT	88.721 2.348 88.753 2.412 ;
			RECT	88.889 2.348 88.921 2.412 ;
			RECT	89.057 2.348 89.089 2.412 ;
			RECT	89.225 2.348 89.257 2.412 ;
			RECT	89.393 2.348 89.425 2.412 ;
			RECT	89.561 2.348 89.593 2.412 ;
			RECT	89.729 2.348 89.761 2.412 ;
			RECT	89.897 2.348 89.929 2.412 ;
			RECT	90.065 2.348 90.097 2.412 ;
			RECT	90.233 2.348 90.265 2.412 ;
			RECT	90.401 2.348 90.433 2.412 ;
			RECT	90.569 2.348 90.601 2.412 ;
			RECT	90.737 2.348 90.769 2.412 ;
			RECT	90.905 2.348 90.937 2.412 ;
			RECT	91.073 2.348 91.105 2.412 ;
			RECT	91.241 2.348 91.273 2.412 ;
			RECT	91.409 2.348 91.441 2.412 ;
			RECT	91.577 2.348 91.609 2.412 ;
			RECT	91.745 2.348 91.777 2.412 ;
			RECT	91.913 2.348 91.945 2.412 ;
			RECT	92.081 2.348 92.113 2.412 ;
			RECT	92.249 2.348 92.281 2.412 ;
			RECT	92.417 2.348 92.449 2.412 ;
			RECT	92.585 2.348 92.617 2.412 ;
			RECT	92.753 2.348 92.785 2.412 ;
			RECT	92.921 2.348 92.953 2.412 ;
			RECT	93.089 2.348 93.121 2.412 ;
			RECT	93.257 2.348 93.289 2.412 ;
			RECT	93.425 2.348 93.457 2.412 ;
			RECT	93.593 2.348 93.625 2.412 ;
			RECT	93.761 2.348 93.793 2.412 ;
			RECT	93.929 2.348 93.961 2.412 ;
			RECT	94.097 2.348 94.129 2.412 ;
			RECT	94.265 2.348 94.297 2.412 ;
			RECT	94.433 2.348 94.465 2.412 ;
			RECT	94.601 2.348 94.633 2.412 ;
			RECT	94.769 2.348 94.801 2.412 ;
			RECT	94.937 2.348 94.969 2.412 ;
			RECT	95.105 2.348 95.137 2.412 ;
			RECT	95.273 2.348 95.305 2.412 ;
			RECT	95.441 2.348 95.473 2.412 ;
			RECT	95.609 2.348 95.641 2.412 ;
			RECT	95.777 2.348 95.809 2.412 ;
			RECT	95.945 2.348 95.977 2.412 ;
			RECT	96.113 2.348 96.145 2.412 ;
			RECT	96.281 2.348 96.313 2.412 ;
			RECT	96.449 2.348 96.481 2.412 ;
			RECT	96.617 2.348 96.649 2.412 ;
			RECT	96.785 2.348 96.817 2.412 ;
			RECT	96.953 2.348 96.985 2.412 ;
			RECT	97.121 2.348 97.153 2.412 ;
			RECT	97.289 2.348 97.321 2.412 ;
			RECT	97.457 2.348 97.489 2.412 ;
			RECT	97.625 2.348 97.657 2.412 ;
			RECT	97.793 2.348 97.825 2.412 ;
			RECT	97.961 2.348 97.993 2.412 ;
			RECT	98.129 2.348 98.161 2.412 ;
			RECT	98.297 2.348 98.329 2.412 ;
			RECT	98.465 2.348 98.497 2.412 ;
			RECT	98.633 2.348 98.665 2.412 ;
			RECT	98.801 2.348 98.833 2.412 ;
			RECT	98.969 2.348 99.001 2.412 ;
			RECT	99.137 2.348 99.169 2.412 ;
			RECT	99.305 2.348 99.337 2.412 ;
			RECT	99.473 2.348 99.505 2.412 ;
			RECT	99.641 2.348 99.673 2.412 ;
			RECT	99.809 2.348 99.841 2.412 ;
			RECT	99.977 2.348 100.009 2.412 ;
			RECT	100.145 2.348 100.177 2.412 ;
			RECT	100.313 2.348 100.345 2.412 ;
			RECT	100.481 2.348 100.513 2.412 ;
			RECT	100.649 2.348 100.681 2.412 ;
			RECT	100.817 2.348 100.849 2.412 ;
			RECT	100.985 2.348 101.017 2.412 ;
			RECT	101.153 2.348 101.185 2.412 ;
			RECT	101.321 2.348 101.353 2.412 ;
			RECT	101.489 2.348 101.521 2.412 ;
			RECT	101.657 2.348 101.689 2.412 ;
			RECT	101.825 2.348 101.857 2.412 ;
			RECT	101.993 2.348 102.025 2.412 ;
			RECT	102.123 2.364 102.155 2.396 ;
			RECT	102.245 2.369 102.277 2.401 ;
			RECT	102.375 2.348 102.407 2.412 ;
			RECT	103.795 2.348 103.827 2.412 ;
			RECT	103.925 2.369 103.957 2.401 ;
			RECT	104.047 2.364 104.079 2.396 ;
			RECT	104.177 2.348 104.209 2.412 ;
			RECT	104.345 2.348 104.377 2.412 ;
			RECT	104.513 2.348 104.545 2.412 ;
			RECT	104.681 2.348 104.713 2.412 ;
			RECT	104.849 2.348 104.881 2.412 ;
			RECT	105.017 2.348 105.049 2.412 ;
			RECT	105.185 2.348 105.217 2.412 ;
			RECT	105.353 2.348 105.385 2.412 ;
			RECT	105.521 2.348 105.553 2.412 ;
			RECT	105.689 2.348 105.721 2.412 ;
			RECT	105.857 2.348 105.889 2.412 ;
			RECT	106.025 2.348 106.057 2.412 ;
			RECT	106.193 2.348 106.225 2.412 ;
			RECT	106.361 2.348 106.393 2.412 ;
			RECT	106.529 2.348 106.561 2.412 ;
			RECT	106.697 2.348 106.729 2.412 ;
			RECT	106.865 2.348 106.897 2.412 ;
			RECT	107.033 2.348 107.065 2.412 ;
			RECT	107.201 2.348 107.233 2.412 ;
			RECT	107.369 2.348 107.401 2.412 ;
			RECT	107.537 2.348 107.569 2.412 ;
			RECT	107.705 2.348 107.737 2.412 ;
			RECT	107.873 2.348 107.905 2.412 ;
			RECT	108.041 2.348 108.073 2.412 ;
			RECT	108.209 2.348 108.241 2.412 ;
			RECT	108.377 2.348 108.409 2.412 ;
			RECT	108.545 2.348 108.577 2.412 ;
			RECT	108.713 2.348 108.745 2.412 ;
			RECT	108.881 2.348 108.913 2.412 ;
			RECT	109.049 2.348 109.081 2.412 ;
			RECT	109.217 2.348 109.249 2.412 ;
			RECT	109.385 2.348 109.417 2.412 ;
			RECT	109.553 2.348 109.585 2.412 ;
			RECT	109.721 2.348 109.753 2.412 ;
			RECT	109.889 2.348 109.921 2.412 ;
			RECT	110.057 2.348 110.089 2.412 ;
			RECT	110.225 2.348 110.257 2.412 ;
			RECT	110.393 2.348 110.425 2.412 ;
			RECT	110.561 2.348 110.593 2.412 ;
			RECT	110.729 2.348 110.761 2.412 ;
			RECT	110.897 2.348 110.929 2.412 ;
			RECT	111.065 2.348 111.097 2.412 ;
			RECT	111.233 2.348 111.265 2.412 ;
			RECT	111.401 2.348 111.433 2.412 ;
			RECT	111.569 2.348 111.601 2.412 ;
			RECT	111.737 2.348 111.769 2.412 ;
			RECT	111.905 2.348 111.937 2.412 ;
			RECT	112.073 2.348 112.105 2.412 ;
			RECT	112.241 2.348 112.273 2.412 ;
			RECT	112.409 2.348 112.441 2.412 ;
			RECT	112.577 2.348 112.609 2.412 ;
			RECT	112.745 2.348 112.777 2.412 ;
			RECT	112.913 2.348 112.945 2.412 ;
			RECT	113.081 2.348 113.113 2.412 ;
			RECT	113.249 2.348 113.281 2.412 ;
			RECT	113.417 2.348 113.449 2.412 ;
			RECT	113.585 2.348 113.617 2.412 ;
			RECT	113.753 2.348 113.785 2.412 ;
			RECT	113.921 2.348 113.953 2.412 ;
			RECT	114.089 2.348 114.121 2.412 ;
			RECT	114.257 2.348 114.289 2.412 ;
			RECT	114.425 2.348 114.457 2.412 ;
			RECT	114.593 2.348 114.625 2.412 ;
			RECT	114.761 2.348 114.793 2.412 ;
			RECT	114.929 2.348 114.961 2.412 ;
			RECT	115.097 2.348 115.129 2.412 ;
			RECT	115.265 2.348 115.297 2.412 ;
			RECT	115.433 2.348 115.465 2.412 ;
			RECT	115.601 2.348 115.633 2.412 ;
			RECT	115.769 2.348 115.801 2.412 ;
			RECT	115.937 2.348 115.969 2.412 ;
			RECT	116.105 2.348 116.137 2.412 ;
			RECT	116.273 2.348 116.305 2.412 ;
			RECT	116.441 2.348 116.473 2.412 ;
			RECT	116.609 2.348 116.641 2.412 ;
			RECT	116.777 2.348 116.809 2.412 ;
			RECT	116.945 2.348 116.977 2.412 ;
			RECT	117.113 2.348 117.145 2.412 ;
			RECT	117.281 2.348 117.313 2.412 ;
			RECT	117.449 2.348 117.481 2.412 ;
			RECT	117.617 2.348 117.649 2.412 ;
			RECT	117.785 2.348 117.817 2.412 ;
			RECT	117.953 2.348 117.985 2.412 ;
			RECT	118.121 2.348 118.153 2.412 ;
			RECT	118.289 2.348 118.321 2.412 ;
			RECT	118.457 2.348 118.489 2.412 ;
			RECT	118.625 2.348 118.657 2.412 ;
			RECT	118.793 2.348 118.825 2.412 ;
			RECT	118.961 2.348 118.993 2.412 ;
			RECT	119.129 2.348 119.161 2.412 ;
			RECT	119.297 2.348 119.329 2.412 ;
			RECT	119.465 2.348 119.497 2.412 ;
			RECT	119.633 2.348 119.665 2.412 ;
			RECT	119.801 2.348 119.833 2.412 ;
			RECT	119.969 2.348 120.001 2.412 ;
			RECT	120.137 2.348 120.169 2.412 ;
			RECT	120.305 2.348 120.337 2.412 ;
			RECT	120.473 2.348 120.505 2.412 ;
			RECT	120.641 2.348 120.673 2.412 ;
			RECT	120.809 2.348 120.841 2.412 ;
			RECT	120.977 2.348 121.009 2.412 ;
			RECT	121.145 2.348 121.177 2.412 ;
			RECT	121.313 2.348 121.345 2.412 ;
			RECT	121.481 2.348 121.513 2.412 ;
			RECT	121.649 2.348 121.681 2.412 ;
			RECT	121.817 2.348 121.849 2.412 ;
			RECT	121.985 2.348 122.017 2.412 ;
			RECT	122.153 2.348 122.185 2.412 ;
			RECT	122.321 2.348 122.353 2.412 ;
			RECT	122.489 2.348 122.521 2.412 ;
			RECT	122.657 2.348 122.689 2.412 ;
			RECT	122.825 2.348 122.857 2.412 ;
			RECT	122.993 2.348 123.025 2.412 ;
			RECT	123.161 2.348 123.193 2.412 ;
			RECT	123.329 2.348 123.361 2.412 ;
			RECT	123.497 2.348 123.529 2.412 ;
			RECT	123.665 2.348 123.697 2.412 ;
			RECT	123.833 2.348 123.865 2.412 ;
			RECT	124.001 2.348 124.033 2.412 ;
			RECT	124.169 2.348 124.201 2.412 ;
			RECT	124.337 2.348 124.369 2.412 ;
			RECT	124.505 2.348 124.537 2.412 ;
			RECT	124.673 2.348 124.705 2.412 ;
			RECT	124.841 2.348 124.873 2.412 ;
			RECT	125.009 2.348 125.041 2.412 ;
			RECT	125.177 2.348 125.209 2.412 ;
			RECT	125.345 2.348 125.377 2.412 ;
			RECT	125.513 2.348 125.545 2.412 ;
			RECT	125.681 2.348 125.713 2.412 ;
			RECT	125.849 2.348 125.881 2.412 ;
			RECT	126.017 2.348 126.049 2.412 ;
			RECT	126.185 2.348 126.217 2.412 ;
			RECT	126.353 2.348 126.385 2.412 ;
			RECT	126.521 2.348 126.553 2.412 ;
			RECT	126.689 2.348 126.721 2.412 ;
			RECT	126.857 2.348 126.889 2.412 ;
			RECT	127.025 2.348 127.057 2.412 ;
			RECT	127.193 2.348 127.225 2.412 ;
			RECT	127.361 2.348 127.393 2.412 ;
			RECT	127.529 2.348 127.561 2.412 ;
			RECT	127.697 2.348 127.729 2.412 ;
			RECT	127.865 2.348 127.897 2.412 ;
			RECT	128.033 2.348 128.065 2.412 ;
			RECT	128.201 2.348 128.233 2.412 ;
			RECT	128.369 2.348 128.401 2.412 ;
			RECT	128.537 2.348 128.569 2.412 ;
			RECT	128.705 2.348 128.737 2.412 ;
			RECT	128.873 2.348 128.905 2.412 ;
			RECT	129.041 2.348 129.073 2.412 ;
			RECT	129.209 2.348 129.241 2.412 ;
			RECT	129.377 2.348 129.409 2.412 ;
			RECT	129.545 2.348 129.577 2.412 ;
			RECT	129.713 2.348 129.745 2.412 ;
			RECT	129.881 2.348 129.913 2.412 ;
			RECT	130.049 2.348 130.081 2.412 ;
			RECT	130.217 2.348 130.249 2.412 ;
			RECT	130.385 2.348 130.417 2.412 ;
			RECT	130.553 2.348 130.585 2.412 ;
			RECT	130.721 2.348 130.753 2.412 ;
			RECT	130.889 2.348 130.921 2.412 ;
			RECT	131.057 2.348 131.089 2.412 ;
			RECT	131.225 2.348 131.257 2.412 ;
			RECT	131.393 2.348 131.425 2.412 ;
			RECT	131.561 2.348 131.593 2.412 ;
			RECT	131.729 2.348 131.761 2.412 ;
			RECT	131.897 2.348 131.929 2.412 ;
			RECT	132.065 2.348 132.097 2.412 ;
			RECT	132.233 2.348 132.265 2.412 ;
			RECT	132.401 2.348 132.433 2.412 ;
			RECT	132.569 2.348 132.601 2.412 ;
			RECT	132.737 2.348 132.769 2.412 ;
			RECT	132.905 2.348 132.937 2.412 ;
			RECT	133.073 2.348 133.105 2.412 ;
			RECT	133.241 2.348 133.273 2.412 ;
			RECT	133.409 2.348 133.441 2.412 ;
			RECT	133.577 2.348 133.609 2.412 ;
			RECT	133.745 2.348 133.777 2.412 ;
			RECT	133.913 2.348 133.945 2.412 ;
			RECT	134.081 2.348 134.113 2.412 ;
			RECT	134.249 2.348 134.281 2.412 ;
			RECT	134.417 2.348 134.449 2.412 ;
			RECT	134.585 2.348 134.617 2.412 ;
			RECT	134.753 2.348 134.785 2.412 ;
			RECT	134.921 2.348 134.953 2.412 ;
			RECT	135.089 2.348 135.121 2.412 ;
			RECT	135.257 2.348 135.289 2.412 ;
			RECT	135.425 2.348 135.457 2.412 ;
			RECT	135.593 2.348 135.625 2.412 ;
			RECT	135.761 2.348 135.793 2.412 ;
			RECT	135.929 2.348 135.961 2.412 ;
			RECT	136.097 2.348 136.129 2.412 ;
			RECT	136.265 2.348 136.297 2.412 ;
			RECT	136.433 2.348 136.465 2.412 ;
			RECT	136.601 2.348 136.633 2.412 ;
			RECT	136.769 2.348 136.801 2.412 ;
			RECT	136.937 2.348 136.969 2.412 ;
			RECT	137.105 2.348 137.137 2.412 ;
			RECT	137.273 2.348 137.305 2.412 ;
			RECT	137.441 2.348 137.473 2.412 ;
			RECT	137.609 2.348 137.641 2.412 ;
			RECT	137.777 2.348 137.809 2.412 ;
			RECT	137.945 2.348 137.977 2.412 ;
			RECT	138.113 2.348 138.145 2.412 ;
			RECT	138.281 2.348 138.313 2.412 ;
			RECT	138.449 2.348 138.481 2.412 ;
			RECT	138.617 2.348 138.649 2.412 ;
			RECT	138.785 2.348 138.817 2.412 ;
			RECT	138.953 2.348 138.985 2.412 ;
			RECT	139.121 2.348 139.153 2.412 ;
			RECT	139.289 2.348 139.321 2.412 ;
			RECT	139.457 2.348 139.489 2.412 ;
			RECT	139.625 2.348 139.657 2.412 ;
			RECT	139.793 2.348 139.825 2.412 ;
			RECT	139.961 2.348 139.993 2.412 ;
			RECT	140.129 2.348 140.161 2.412 ;
			RECT	140.297 2.348 140.329 2.412 ;
			RECT	140.465 2.348 140.497 2.412 ;
			RECT	140.633 2.348 140.665 2.412 ;
			RECT	140.801 2.348 140.833 2.412 ;
			RECT	140.969 2.348 141.001 2.412 ;
			RECT	141.137 2.348 141.169 2.412 ;
			RECT	141.305 2.348 141.337 2.412 ;
			RECT	141.473 2.348 141.505 2.412 ;
			RECT	141.641 2.348 141.673 2.412 ;
			RECT	141.809 2.348 141.841 2.412 ;
			RECT	141.977 2.348 142.009 2.412 ;
			RECT	142.145 2.348 142.177 2.412 ;
			RECT	142.313 2.348 142.345 2.412 ;
			RECT	142.481 2.348 142.513 2.412 ;
			RECT	142.649 2.348 142.681 2.412 ;
			RECT	142.817 2.348 142.849 2.412 ;
			RECT	142.985 2.348 143.017 2.412 ;
			RECT	143.153 2.348 143.185 2.412 ;
			RECT	143.321 2.348 143.353 2.412 ;
			RECT	143.489 2.348 143.521 2.412 ;
			RECT	143.657 2.348 143.689 2.412 ;
			RECT	143.825 2.348 143.857 2.412 ;
			RECT	143.993 2.348 144.025 2.412 ;
			RECT	144.161 2.348 144.193 2.412 ;
			RECT	144.329 2.348 144.361 2.412 ;
			RECT	144.497 2.348 144.529 2.412 ;
			RECT	144.665 2.348 144.697 2.412 ;
			RECT	144.833 2.348 144.865 2.412 ;
			RECT	145.001 2.348 145.033 2.412 ;
			RECT	145.169 2.348 145.201 2.412 ;
			RECT	145.337 2.348 145.369 2.412 ;
			RECT	145.505 2.348 145.537 2.412 ;
			RECT	145.673 2.348 145.705 2.412 ;
			RECT	145.841 2.348 145.873 2.412 ;
			RECT	146.009 2.348 146.041 2.412 ;
			RECT	146.177 2.348 146.209 2.412 ;
			RECT	146.345 2.348 146.377 2.412 ;
			RECT	146.513 2.348 146.545 2.412 ;
			RECT	146.681 2.348 146.713 2.412 ;
			RECT	146.849 2.348 146.881 2.412 ;
			RECT	147.017 2.348 147.049 2.412 ;
			RECT	147.185 2.348 147.217 2.412 ;
			RECT	147.316 2.364 147.348 2.396 ;
			RECT	147.437 2.364 147.469 2.396 ;
			RECT	147.567 2.348 147.599 2.412 ;
			RECT	149.879 2.348 149.911 2.412 ;
			RECT	151.13 2.348 151.194 2.412 ;
			RECT	151.81 2.348 151.842 2.412 ;
			RECT	152.249 2.348 152.281 2.412 ;
			RECT	153.56 2.348 153.624 2.412 ;
			RECT	156.601 2.348 156.633 2.412 ;
			RECT	156.731 2.364 156.763 2.396 ;
			RECT	156.852 2.364 156.884 2.396 ;
			RECT	156.983 2.348 157.015 2.412 ;
			RECT	157.151 2.348 157.183 2.412 ;
			RECT	157.319 2.348 157.351 2.412 ;
			RECT	157.487 2.348 157.519 2.412 ;
			RECT	157.655 2.348 157.687 2.412 ;
			RECT	157.823 2.348 157.855 2.412 ;
			RECT	157.991 2.348 158.023 2.412 ;
			RECT	158.159 2.348 158.191 2.412 ;
			RECT	158.327 2.348 158.359 2.412 ;
			RECT	158.495 2.348 158.527 2.412 ;
			RECT	158.663 2.348 158.695 2.412 ;
			RECT	158.831 2.348 158.863 2.412 ;
			RECT	158.999 2.348 159.031 2.412 ;
			RECT	159.167 2.348 159.199 2.412 ;
			RECT	159.335 2.348 159.367 2.412 ;
			RECT	159.503 2.348 159.535 2.412 ;
			RECT	159.671 2.348 159.703 2.412 ;
			RECT	159.839 2.348 159.871 2.412 ;
			RECT	160.007 2.348 160.039 2.412 ;
			RECT	160.175 2.348 160.207 2.412 ;
			RECT	160.343 2.348 160.375 2.412 ;
			RECT	160.511 2.348 160.543 2.412 ;
			RECT	160.679 2.348 160.711 2.412 ;
			RECT	160.847 2.348 160.879 2.412 ;
			RECT	161.015 2.348 161.047 2.412 ;
			RECT	161.183 2.348 161.215 2.412 ;
			RECT	161.351 2.348 161.383 2.412 ;
			RECT	161.519 2.348 161.551 2.412 ;
			RECT	161.687 2.348 161.719 2.412 ;
			RECT	161.855 2.348 161.887 2.412 ;
			RECT	162.023 2.348 162.055 2.412 ;
			RECT	162.191 2.348 162.223 2.412 ;
			RECT	162.359 2.348 162.391 2.412 ;
			RECT	162.527 2.348 162.559 2.412 ;
			RECT	162.695 2.348 162.727 2.412 ;
			RECT	162.863 2.348 162.895 2.412 ;
			RECT	163.031 2.348 163.063 2.412 ;
			RECT	163.199 2.348 163.231 2.412 ;
			RECT	163.367 2.348 163.399 2.412 ;
			RECT	163.535 2.348 163.567 2.412 ;
			RECT	163.703 2.348 163.735 2.412 ;
			RECT	163.871 2.348 163.903 2.412 ;
			RECT	164.039 2.348 164.071 2.412 ;
			RECT	164.207 2.348 164.239 2.412 ;
			RECT	164.375 2.348 164.407 2.412 ;
			RECT	164.543 2.348 164.575 2.412 ;
			RECT	164.711 2.348 164.743 2.412 ;
			RECT	164.879 2.348 164.911 2.412 ;
			RECT	165.047 2.348 165.079 2.412 ;
			RECT	165.215 2.348 165.247 2.412 ;
			RECT	165.383 2.348 165.415 2.412 ;
			RECT	165.551 2.348 165.583 2.412 ;
			RECT	165.719 2.348 165.751 2.412 ;
			RECT	165.887 2.348 165.919 2.412 ;
			RECT	166.055 2.348 166.087 2.412 ;
			RECT	166.223 2.348 166.255 2.412 ;
			RECT	166.391 2.348 166.423 2.412 ;
			RECT	166.559 2.348 166.591 2.412 ;
			RECT	166.727 2.348 166.759 2.412 ;
			RECT	166.895 2.348 166.927 2.412 ;
			RECT	167.063 2.348 167.095 2.412 ;
			RECT	167.231 2.348 167.263 2.412 ;
			RECT	167.399 2.348 167.431 2.412 ;
			RECT	167.567 2.348 167.599 2.412 ;
			RECT	167.735 2.348 167.767 2.412 ;
			RECT	167.903 2.348 167.935 2.412 ;
			RECT	168.071 2.348 168.103 2.412 ;
			RECT	168.239 2.348 168.271 2.412 ;
			RECT	168.407 2.348 168.439 2.412 ;
			RECT	168.575 2.348 168.607 2.412 ;
			RECT	168.743 2.348 168.775 2.412 ;
			RECT	168.911 2.348 168.943 2.412 ;
			RECT	169.079 2.348 169.111 2.412 ;
			RECT	169.247 2.348 169.279 2.412 ;
			RECT	169.415 2.348 169.447 2.412 ;
			RECT	169.583 2.348 169.615 2.412 ;
			RECT	169.751 2.348 169.783 2.412 ;
			RECT	169.919 2.348 169.951 2.412 ;
			RECT	170.087 2.348 170.119 2.412 ;
			RECT	170.255 2.348 170.287 2.412 ;
			RECT	170.423 2.348 170.455 2.412 ;
			RECT	170.591 2.348 170.623 2.412 ;
			RECT	170.759 2.348 170.791 2.412 ;
			RECT	170.927 2.348 170.959 2.412 ;
			RECT	171.095 2.348 171.127 2.412 ;
			RECT	171.263 2.348 171.295 2.412 ;
			RECT	171.431 2.348 171.463 2.412 ;
			RECT	171.599 2.348 171.631 2.412 ;
			RECT	171.767 2.348 171.799 2.412 ;
			RECT	171.935 2.348 171.967 2.412 ;
			RECT	172.103 2.348 172.135 2.412 ;
			RECT	172.271 2.348 172.303 2.412 ;
			RECT	172.439 2.348 172.471 2.412 ;
			RECT	172.607 2.348 172.639 2.412 ;
			RECT	172.775 2.348 172.807 2.412 ;
			RECT	172.943 2.348 172.975 2.412 ;
			RECT	173.111 2.348 173.143 2.412 ;
			RECT	173.279 2.348 173.311 2.412 ;
			RECT	173.447 2.348 173.479 2.412 ;
			RECT	173.615 2.348 173.647 2.412 ;
			RECT	173.783 2.348 173.815 2.412 ;
			RECT	173.951 2.348 173.983 2.412 ;
			RECT	174.119 2.348 174.151 2.412 ;
			RECT	174.287 2.348 174.319 2.412 ;
			RECT	174.455 2.348 174.487 2.412 ;
			RECT	174.623 2.348 174.655 2.412 ;
			RECT	174.791 2.348 174.823 2.412 ;
			RECT	174.959 2.348 174.991 2.412 ;
			RECT	175.127 2.348 175.159 2.412 ;
			RECT	175.295 2.348 175.327 2.412 ;
			RECT	175.463 2.348 175.495 2.412 ;
			RECT	175.631 2.348 175.663 2.412 ;
			RECT	175.799 2.348 175.831 2.412 ;
			RECT	175.967 2.348 175.999 2.412 ;
			RECT	176.135 2.348 176.167 2.412 ;
			RECT	176.303 2.348 176.335 2.412 ;
			RECT	176.471 2.348 176.503 2.412 ;
			RECT	176.639 2.348 176.671 2.412 ;
			RECT	176.807 2.348 176.839 2.412 ;
			RECT	176.975 2.348 177.007 2.412 ;
			RECT	177.143 2.348 177.175 2.412 ;
			RECT	177.311 2.348 177.343 2.412 ;
			RECT	177.479 2.348 177.511 2.412 ;
			RECT	177.647 2.348 177.679 2.412 ;
			RECT	177.815 2.348 177.847 2.412 ;
			RECT	177.983 2.348 178.015 2.412 ;
			RECT	178.151 2.348 178.183 2.412 ;
			RECT	178.319 2.348 178.351 2.412 ;
			RECT	178.487 2.348 178.519 2.412 ;
			RECT	178.655 2.348 178.687 2.412 ;
			RECT	178.823 2.348 178.855 2.412 ;
			RECT	178.991 2.348 179.023 2.412 ;
			RECT	179.159 2.348 179.191 2.412 ;
			RECT	179.327 2.348 179.359 2.412 ;
			RECT	179.495 2.348 179.527 2.412 ;
			RECT	179.663 2.348 179.695 2.412 ;
			RECT	179.831 2.348 179.863 2.412 ;
			RECT	179.999 2.348 180.031 2.412 ;
			RECT	180.167 2.348 180.199 2.412 ;
			RECT	180.335 2.348 180.367 2.412 ;
			RECT	180.503 2.348 180.535 2.412 ;
			RECT	180.671 2.348 180.703 2.412 ;
			RECT	180.839 2.348 180.871 2.412 ;
			RECT	181.007 2.348 181.039 2.412 ;
			RECT	181.175 2.348 181.207 2.412 ;
			RECT	181.343 2.348 181.375 2.412 ;
			RECT	181.511 2.348 181.543 2.412 ;
			RECT	181.679 2.348 181.711 2.412 ;
			RECT	181.847 2.348 181.879 2.412 ;
			RECT	182.015 2.348 182.047 2.412 ;
			RECT	182.183 2.348 182.215 2.412 ;
			RECT	182.351 2.348 182.383 2.412 ;
			RECT	182.519 2.348 182.551 2.412 ;
			RECT	182.687 2.348 182.719 2.412 ;
			RECT	182.855 2.348 182.887 2.412 ;
			RECT	183.023 2.348 183.055 2.412 ;
			RECT	183.191 2.348 183.223 2.412 ;
			RECT	183.359 2.348 183.391 2.412 ;
			RECT	183.527 2.348 183.559 2.412 ;
			RECT	183.695 2.348 183.727 2.412 ;
			RECT	183.863 2.348 183.895 2.412 ;
			RECT	184.031 2.348 184.063 2.412 ;
			RECT	184.199 2.348 184.231 2.412 ;
			RECT	184.367 2.348 184.399 2.412 ;
			RECT	184.535 2.348 184.567 2.412 ;
			RECT	184.703 2.348 184.735 2.412 ;
			RECT	184.871 2.348 184.903 2.412 ;
			RECT	185.039 2.348 185.071 2.412 ;
			RECT	185.207 2.348 185.239 2.412 ;
			RECT	185.375 2.348 185.407 2.412 ;
			RECT	185.543 2.348 185.575 2.412 ;
			RECT	185.711 2.348 185.743 2.412 ;
			RECT	185.879 2.348 185.911 2.412 ;
			RECT	186.047 2.348 186.079 2.412 ;
			RECT	186.215 2.348 186.247 2.412 ;
			RECT	186.383 2.348 186.415 2.412 ;
			RECT	186.551 2.348 186.583 2.412 ;
			RECT	186.719 2.348 186.751 2.412 ;
			RECT	186.887 2.348 186.919 2.412 ;
			RECT	187.055 2.348 187.087 2.412 ;
			RECT	187.223 2.348 187.255 2.412 ;
			RECT	187.391 2.348 187.423 2.412 ;
			RECT	187.559 2.348 187.591 2.412 ;
			RECT	187.727 2.348 187.759 2.412 ;
			RECT	187.895 2.348 187.927 2.412 ;
			RECT	188.063 2.348 188.095 2.412 ;
			RECT	188.231 2.348 188.263 2.412 ;
			RECT	188.399 2.348 188.431 2.412 ;
			RECT	188.567 2.348 188.599 2.412 ;
			RECT	188.735 2.348 188.767 2.412 ;
			RECT	188.903 2.348 188.935 2.412 ;
			RECT	189.071 2.348 189.103 2.412 ;
			RECT	189.239 2.348 189.271 2.412 ;
			RECT	189.407 2.348 189.439 2.412 ;
			RECT	189.575 2.348 189.607 2.412 ;
			RECT	189.743 2.348 189.775 2.412 ;
			RECT	189.911 2.348 189.943 2.412 ;
			RECT	190.079 2.348 190.111 2.412 ;
			RECT	190.247 2.348 190.279 2.412 ;
			RECT	190.415 2.348 190.447 2.412 ;
			RECT	190.583 2.348 190.615 2.412 ;
			RECT	190.751 2.348 190.783 2.412 ;
			RECT	190.919 2.348 190.951 2.412 ;
			RECT	191.087 2.348 191.119 2.412 ;
			RECT	191.255 2.348 191.287 2.412 ;
			RECT	191.423 2.348 191.455 2.412 ;
			RECT	191.591 2.348 191.623 2.412 ;
			RECT	191.759 2.348 191.791 2.412 ;
			RECT	191.927 2.348 191.959 2.412 ;
			RECT	192.095 2.348 192.127 2.412 ;
			RECT	192.263 2.348 192.295 2.412 ;
			RECT	192.431 2.348 192.463 2.412 ;
			RECT	192.599 2.348 192.631 2.412 ;
			RECT	192.767 2.348 192.799 2.412 ;
			RECT	192.935 2.348 192.967 2.412 ;
			RECT	193.103 2.348 193.135 2.412 ;
			RECT	193.271 2.348 193.303 2.412 ;
			RECT	193.439 2.348 193.471 2.412 ;
			RECT	193.607 2.348 193.639 2.412 ;
			RECT	193.775 2.348 193.807 2.412 ;
			RECT	193.943 2.348 193.975 2.412 ;
			RECT	194.111 2.348 194.143 2.412 ;
			RECT	194.279 2.348 194.311 2.412 ;
			RECT	194.447 2.348 194.479 2.412 ;
			RECT	194.615 2.348 194.647 2.412 ;
			RECT	194.783 2.348 194.815 2.412 ;
			RECT	194.951 2.348 194.983 2.412 ;
			RECT	195.119 2.348 195.151 2.412 ;
			RECT	195.287 2.348 195.319 2.412 ;
			RECT	195.455 2.348 195.487 2.412 ;
			RECT	195.623 2.348 195.655 2.412 ;
			RECT	195.791 2.348 195.823 2.412 ;
			RECT	195.959 2.348 195.991 2.412 ;
			RECT	196.127 2.348 196.159 2.412 ;
			RECT	196.295 2.348 196.327 2.412 ;
			RECT	196.463 2.348 196.495 2.412 ;
			RECT	196.631 2.348 196.663 2.412 ;
			RECT	196.799 2.348 196.831 2.412 ;
			RECT	196.967 2.348 196.999 2.412 ;
			RECT	197.135 2.348 197.167 2.412 ;
			RECT	197.303 2.348 197.335 2.412 ;
			RECT	197.471 2.348 197.503 2.412 ;
			RECT	197.639 2.348 197.671 2.412 ;
			RECT	197.807 2.348 197.839 2.412 ;
			RECT	197.975 2.348 198.007 2.412 ;
			RECT	198.143 2.348 198.175 2.412 ;
			RECT	198.311 2.348 198.343 2.412 ;
			RECT	198.479 2.348 198.511 2.412 ;
			RECT	198.647 2.348 198.679 2.412 ;
			RECT	198.815 2.348 198.847 2.412 ;
			RECT	198.983 2.348 199.015 2.412 ;
			RECT	199.151 2.348 199.183 2.412 ;
			RECT	199.319 2.348 199.351 2.412 ;
			RECT	199.487 2.348 199.519 2.412 ;
			RECT	199.655 2.348 199.687 2.412 ;
			RECT	199.823 2.348 199.855 2.412 ;
			RECT	199.991 2.348 200.023 2.412 ;
			RECT	200.121 2.364 200.153 2.396 ;
			RECT	200.243 2.369 200.275 2.401 ;
			RECT	200.373 2.348 200.405 2.412 ;
			RECT	200.9 2.348 200.932 2.412 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 72.056 201.665 72.176 ;
			LAYER	J3 ;
			RECT	0.755 72.084 0.787 72.148 ;
			RECT	1.645 72.084 1.709 72.148 ;
			RECT	2.323 72.084 2.387 72.148 ;
			RECT	3.438 72.084 3.47 72.148 ;
			RECT	3.585 72.084 3.617 72.148 ;
			RECT	4.195 72.084 4.227 72.148 ;
			RECT	4.72 72.084 4.752 72.148 ;
			RECT	4.944 72.084 5.008 72.148 ;
			RECT	5.267 72.084 5.299 72.148 ;
			RECT	5.797 72.084 5.829 72.148 ;
			RECT	5.927 72.095 5.959 72.127 ;
			RECT	6.049 72.1 6.081 72.132 ;
			RECT	6.179 72.084 6.211 72.148 ;
			RECT	6.347 72.084 6.379 72.148 ;
			RECT	6.515 72.084 6.547 72.148 ;
			RECT	6.683 72.084 6.715 72.148 ;
			RECT	6.851 72.084 6.883 72.148 ;
			RECT	7.019 72.084 7.051 72.148 ;
			RECT	7.187 72.084 7.219 72.148 ;
			RECT	7.355 72.084 7.387 72.148 ;
			RECT	7.523 72.084 7.555 72.148 ;
			RECT	7.691 72.084 7.723 72.148 ;
			RECT	7.859 72.084 7.891 72.148 ;
			RECT	8.027 72.084 8.059 72.148 ;
			RECT	8.195 72.084 8.227 72.148 ;
			RECT	8.363 72.084 8.395 72.148 ;
			RECT	8.531 72.084 8.563 72.148 ;
			RECT	8.699 72.084 8.731 72.148 ;
			RECT	8.867 72.084 8.899 72.148 ;
			RECT	9.035 72.084 9.067 72.148 ;
			RECT	9.203 72.084 9.235 72.148 ;
			RECT	9.371 72.084 9.403 72.148 ;
			RECT	9.539 72.084 9.571 72.148 ;
			RECT	9.707 72.084 9.739 72.148 ;
			RECT	9.875 72.084 9.907 72.148 ;
			RECT	10.043 72.084 10.075 72.148 ;
			RECT	10.211 72.084 10.243 72.148 ;
			RECT	10.379 72.084 10.411 72.148 ;
			RECT	10.547 72.084 10.579 72.148 ;
			RECT	10.715 72.084 10.747 72.148 ;
			RECT	10.883 72.084 10.915 72.148 ;
			RECT	11.051 72.084 11.083 72.148 ;
			RECT	11.219 72.084 11.251 72.148 ;
			RECT	11.387 72.084 11.419 72.148 ;
			RECT	11.555 72.084 11.587 72.148 ;
			RECT	11.723 72.084 11.755 72.148 ;
			RECT	11.891 72.084 11.923 72.148 ;
			RECT	12.059 72.084 12.091 72.148 ;
			RECT	12.227 72.084 12.259 72.148 ;
			RECT	12.395 72.084 12.427 72.148 ;
			RECT	12.563 72.084 12.595 72.148 ;
			RECT	12.731 72.084 12.763 72.148 ;
			RECT	12.899 72.084 12.931 72.148 ;
			RECT	13.067 72.084 13.099 72.148 ;
			RECT	13.235 72.084 13.267 72.148 ;
			RECT	13.403 72.084 13.435 72.148 ;
			RECT	13.571 72.084 13.603 72.148 ;
			RECT	13.739 72.084 13.771 72.148 ;
			RECT	13.907 72.084 13.939 72.148 ;
			RECT	14.075 72.084 14.107 72.148 ;
			RECT	14.243 72.084 14.275 72.148 ;
			RECT	14.411 72.084 14.443 72.148 ;
			RECT	14.579 72.084 14.611 72.148 ;
			RECT	14.747 72.084 14.779 72.148 ;
			RECT	14.915 72.084 14.947 72.148 ;
			RECT	15.083 72.084 15.115 72.148 ;
			RECT	15.251 72.084 15.283 72.148 ;
			RECT	15.419 72.084 15.451 72.148 ;
			RECT	15.587 72.084 15.619 72.148 ;
			RECT	15.755 72.084 15.787 72.148 ;
			RECT	15.923 72.084 15.955 72.148 ;
			RECT	16.091 72.084 16.123 72.148 ;
			RECT	16.259 72.084 16.291 72.148 ;
			RECT	16.427 72.084 16.459 72.148 ;
			RECT	16.595 72.084 16.627 72.148 ;
			RECT	16.763 72.084 16.795 72.148 ;
			RECT	16.931 72.084 16.963 72.148 ;
			RECT	17.099 72.084 17.131 72.148 ;
			RECT	17.267 72.084 17.299 72.148 ;
			RECT	17.435 72.084 17.467 72.148 ;
			RECT	17.603 72.084 17.635 72.148 ;
			RECT	17.771 72.084 17.803 72.148 ;
			RECT	17.939 72.084 17.971 72.148 ;
			RECT	18.107 72.084 18.139 72.148 ;
			RECT	18.275 72.084 18.307 72.148 ;
			RECT	18.443 72.084 18.475 72.148 ;
			RECT	18.611 72.084 18.643 72.148 ;
			RECT	18.779 72.084 18.811 72.148 ;
			RECT	18.947 72.084 18.979 72.148 ;
			RECT	19.115 72.084 19.147 72.148 ;
			RECT	19.283 72.084 19.315 72.148 ;
			RECT	19.451 72.084 19.483 72.148 ;
			RECT	19.619 72.084 19.651 72.148 ;
			RECT	19.787 72.084 19.819 72.148 ;
			RECT	19.955 72.084 19.987 72.148 ;
			RECT	20.123 72.084 20.155 72.148 ;
			RECT	20.291 72.084 20.323 72.148 ;
			RECT	20.459 72.084 20.491 72.148 ;
			RECT	20.627 72.084 20.659 72.148 ;
			RECT	20.795 72.084 20.827 72.148 ;
			RECT	20.963 72.084 20.995 72.148 ;
			RECT	21.131 72.084 21.163 72.148 ;
			RECT	21.299 72.084 21.331 72.148 ;
			RECT	21.467 72.084 21.499 72.148 ;
			RECT	21.635 72.084 21.667 72.148 ;
			RECT	21.803 72.084 21.835 72.148 ;
			RECT	21.971 72.084 22.003 72.148 ;
			RECT	22.139 72.084 22.171 72.148 ;
			RECT	22.307 72.084 22.339 72.148 ;
			RECT	22.475 72.084 22.507 72.148 ;
			RECT	22.643 72.084 22.675 72.148 ;
			RECT	22.811 72.084 22.843 72.148 ;
			RECT	22.979 72.084 23.011 72.148 ;
			RECT	23.147 72.084 23.179 72.148 ;
			RECT	23.315 72.084 23.347 72.148 ;
			RECT	23.483 72.084 23.515 72.148 ;
			RECT	23.651 72.084 23.683 72.148 ;
			RECT	23.819 72.084 23.851 72.148 ;
			RECT	23.987 72.084 24.019 72.148 ;
			RECT	24.155 72.084 24.187 72.148 ;
			RECT	24.323 72.084 24.355 72.148 ;
			RECT	24.491 72.084 24.523 72.148 ;
			RECT	24.659 72.084 24.691 72.148 ;
			RECT	24.827 72.084 24.859 72.148 ;
			RECT	24.995 72.084 25.027 72.148 ;
			RECT	25.163 72.084 25.195 72.148 ;
			RECT	25.331 72.084 25.363 72.148 ;
			RECT	25.499 72.084 25.531 72.148 ;
			RECT	25.667 72.084 25.699 72.148 ;
			RECT	25.835 72.084 25.867 72.148 ;
			RECT	26.003 72.084 26.035 72.148 ;
			RECT	26.171 72.084 26.203 72.148 ;
			RECT	26.339 72.084 26.371 72.148 ;
			RECT	26.507 72.084 26.539 72.148 ;
			RECT	26.675 72.084 26.707 72.148 ;
			RECT	26.843 72.084 26.875 72.148 ;
			RECT	27.011 72.084 27.043 72.148 ;
			RECT	27.179 72.084 27.211 72.148 ;
			RECT	27.347 72.084 27.379 72.148 ;
			RECT	27.515 72.084 27.547 72.148 ;
			RECT	27.683 72.084 27.715 72.148 ;
			RECT	27.851 72.084 27.883 72.148 ;
			RECT	28.019 72.084 28.051 72.148 ;
			RECT	28.187 72.084 28.219 72.148 ;
			RECT	28.355 72.084 28.387 72.148 ;
			RECT	28.523 72.084 28.555 72.148 ;
			RECT	28.691 72.084 28.723 72.148 ;
			RECT	28.859 72.084 28.891 72.148 ;
			RECT	29.027 72.084 29.059 72.148 ;
			RECT	29.195 72.084 29.227 72.148 ;
			RECT	29.363 72.084 29.395 72.148 ;
			RECT	29.531 72.084 29.563 72.148 ;
			RECT	29.699 72.084 29.731 72.148 ;
			RECT	29.867 72.084 29.899 72.148 ;
			RECT	30.035 72.084 30.067 72.148 ;
			RECT	30.203 72.084 30.235 72.148 ;
			RECT	30.371 72.084 30.403 72.148 ;
			RECT	30.539 72.084 30.571 72.148 ;
			RECT	30.707 72.084 30.739 72.148 ;
			RECT	30.875 72.084 30.907 72.148 ;
			RECT	31.043 72.084 31.075 72.148 ;
			RECT	31.211 72.084 31.243 72.148 ;
			RECT	31.379 72.084 31.411 72.148 ;
			RECT	31.547 72.084 31.579 72.148 ;
			RECT	31.715 72.084 31.747 72.148 ;
			RECT	31.883 72.084 31.915 72.148 ;
			RECT	32.051 72.084 32.083 72.148 ;
			RECT	32.219 72.084 32.251 72.148 ;
			RECT	32.387 72.084 32.419 72.148 ;
			RECT	32.555 72.084 32.587 72.148 ;
			RECT	32.723 72.084 32.755 72.148 ;
			RECT	32.891 72.084 32.923 72.148 ;
			RECT	33.059 72.084 33.091 72.148 ;
			RECT	33.227 72.084 33.259 72.148 ;
			RECT	33.395 72.084 33.427 72.148 ;
			RECT	33.563 72.084 33.595 72.148 ;
			RECT	33.731 72.084 33.763 72.148 ;
			RECT	33.899 72.084 33.931 72.148 ;
			RECT	34.067 72.084 34.099 72.148 ;
			RECT	34.235 72.084 34.267 72.148 ;
			RECT	34.403 72.084 34.435 72.148 ;
			RECT	34.571 72.084 34.603 72.148 ;
			RECT	34.739 72.084 34.771 72.148 ;
			RECT	34.907 72.084 34.939 72.148 ;
			RECT	35.075 72.084 35.107 72.148 ;
			RECT	35.243 72.084 35.275 72.148 ;
			RECT	35.411 72.084 35.443 72.148 ;
			RECT	35.579 72.084 35.611 72.148 ;
			RECT	35.747 72.084 35.779 72.148 ;
			RECT	35.915 72.084 35.947 72.148 ;
			RECT	36.083 72.084 36.115 72.148 ;
			RECT	36.251 72.084 36.283 72.148 ;
			RECT	36.419 72.084 36.451 72.148 ;
			RECT	36.587 72.084 36.619 72.148 ;
			RECT	36.755 72.084 36.787 72.148 ;
			RECT	36.923 72.084 36.955 72.148 ;
			RECT	37.091 72.084 37.123 72.148 ;
			RECT	37.259 72.084 37.291 72.148 ;
			RECT	37.427 72.084 37.459 72.148 ;
			RECT	37.595 72.084 37.627 72.148 ;
			RECT	37.763 72.084 37.795 72.148 ;
			RECT	37.931 72.084 37.963 72.148 ;
			RECT	38.099 72.084 38.131 72.148 ;
			RECT	38.267 72.084 38.299 72.148 ;
			RECT	38.435 72.084 38.467 72.148 ;
			RECT	38.603 72.084 38.635 72.148 ;
			RECT	38.771 72.084 38.803 72.148 ;
			RECT	38.939 72.084 38.971 72.148 ;
			RECT	39.107 72.084 39.139 72.148 ;
			RECT	39.275 72.084 39.307 72.148 ;
			RECT	39.443 72.084 39.475 72.148 ;
			RECT	39.611 72.084 39.643 72.148 ;
			RECT	39.779 72.084 39.811 72.148 ;
			RECT	39.947 72.084 39.979 72.148 ;
			RECT	40.115 72.084 40.147 72.148 ;
			RECT	40.283 72.084 40.315 72.148 ;
			RECT	40.451 72.084 40.483 72.148 ;
			RECT	40.619 72.084 40.651 72.148 ;
			RECT	40.787 72.084 40.819 72.148 ;
			RECT	40.955 72.084 40.987 72.148 ;
			RECT	41.123 72.084 41.155 72.148 ;
			RECT	41.291 72.084 41.323 72.148 ;
			RECT	41.459 72.084 41.491 72.148 ;
			RECT	41.627 72.084 41.659 72.148 ;
			RECT	41.795 72.084 41.827 72.148 ;
			RECT	41.963 72.084 41.995 72.148 ;
			RECT	42.131 72.084 42.163 72.148 ;
			RECT	42.299 72.084 42.331 72.148 ;
			RECT	42.467 72.084 42.499 72.148 ;
			RECT	42.635 72.084 42.667 72.148 ;
			RECT	42.803 72.084 42.835 72.148 ;
			RECT	42.971 72.084 43.003 72.148 ;
			RECT	43.139 72.084 43.171 72.148 ;
			RECT	43.307 72.084 43.339 72.148 ;
			RECT	43.475 72.084 43.507 72.148 ;
			RECT	43.643 72.084 43.675 72.148 ;
			RECT	43.811 72.084 43.843 72.148 ;
			RECT	43.979 72.084 44.011 72.148 ;
			RECT	44.147 72.084 44.179 72.148 ;
			RECT	44.315 72.084 44.347 72.148 ;
			RECT	44.483 72.084 44.515 72.148 ;
			RECT	44.651 72.084 44.683 72.148 ;
			RECT	44.819 72.084 44.851 72.148 ;
			RECT	44.987 72.084 45.019 72.148 ;
			RECT	45.155 72.084 45.187 72.148 ;
			RECT	45.323 72.084 45.355 72.148 ;
			RECT	45.491 72.084 45.523 72.148 ;
			RECT	45.659 72.084 45.691 72.148 ;
			RECT	45.827 72.084 45.859 72.148 ;
			RECT	45.995 72.084 46.027 72.148 ;
			RECT	46.163 72.084 46.195 72.148 ;
			RECT	46.331 72.084 46.363 72.148 ;
			RECT	46.499 72.084 46.531 72.148 ;
			RECT	46.667 72.084 46.699 72.148 ;
			RECT	46.835 72.084 46.867 72.148 ;
			RECT	47.003 72.084 47.035 72.148 ;
			RECT	47.171 72.084 47.203 72.148 ;
			RECT	47.339 72.084 47.371 72.148 ;
			RECT	47.507 72.084 47.539 72.148 ;
			RECT	47.675 72.084 47.707 72.148 ;
			RECT	47.843 72.084 47.875 72.148 ;
			RECT	48.011 72.084 48.043 72.148 ;
			RECT	48.179 72.084 48.211 72.148 ;
			RECT	48.347 72.084 48.379 72.148 ;
			RECT	48.515 72.084 48.547 72.148 ;
			RECT	48.683 72.084 48.715 72.148 ;
			RECT	48.851 72.084 48.883 72.148 ;
			RECT	49.019 72.084 49.051 72.148 ;
			RECT	49.187 72.084 49.219 72.148 ;
			RECT	49.318 72.1 49.35 72.132 ;
			RECT	49.439 72.1 49.471 72.132 ;
			RECT	49.569 72.084 49.601 72.148 ;
			RECT	51.881 72.084 51.913 72.148 ;
			RECT	53.132 72.084 53.196 72.148 ;
			RECT	53.812 72.084 53.844 72.148 ;
			RECT	54.251 72.084 54.283 72.148 ;
			RECT	55.562 72.084 55.626 72.148 ;
			RECT	58.603 72.084 58.635 72.148 ;
			RECT	58.733 72.1 58.765 72.132 ;
			RECT	58.854 72.1 58.886 72.132 ;
			RECT	58.985 72.084 59.017 72.148 ;
			RECT	59.153 72.084 59.185 72.148 ;
			RECT	59.321 72.084 59.353 72.148 ;
			RECT	59.489 72.084 59.521 72.148 ;
			RECT	59.657 72.084 59.689 72.148 ;
			RECT	59.825 72.084 59.857 72.148 ;
			RECT	59.993 72.084 60.025 72.148 ;
			RECT	60.161 72.084 60.193 72.148 ;
			RECT	60.329 72.084 60.361 72.148 ;
			RECT	60.497 72.084 60.529 72.148 ;
			RECT	60.665 72.084 60.697 72.148 ;
			RECT	60.833 72.084 60.865 72.148 ;
			RECT	61.001 72.084 61.033 72.148 ;
			RECT	61.169 72.084 61.201 72.148 ;
			RECT	61.337 72.084 61.369 72.148 ;
			RECT	61.505 72.084 61.537 72.148 ;
			RECT	61.673 72.084 61.705 72.148 ;
			RECT	61.841 72.084 61.873 72.148 ;
			RECT	62.009 72.084 62.041 72.148 ;
			RECT	62.177 72.084 62.209 72.148 ;
			RECT	62.345 72.084 62.377 72.148 ;
			RECT	62.513 72.084 62.545 72.148 ;
			RECT	62.681 72.084 62.713 72.148 ;
			RECT	62.849 72.084 62.881 72.148 ;
			RECT	63.017 72.084 63.049 72.148 ;
			RECT	63.185 72.084 63.217 72.148 ;
			RECT	63.353 72.084 63.385 72.148 ;
			RECT	63.521 72.084 63.553 72.148 ;
			RECT	63.689 72.084 63.721 72.148 ;
			RECT	63.857 72.084 63.889 72.148 ;
			RECT	64.025 72.084 64.057 72.148 ;
			RECT	64.193 72.084 64.225 72.148 ;
			RECT	64.361 72.084 64.393 72.148 ;
			RECT	64.529 72.084 64.561 72.148 ;
			RECT	64.697 72.084 64.729 72.148 ;
			RECT	64.865 72.084 64.897 72.148 ;
			RECT	65.033 72.084 65.065 72.148 ;
			RECT	65.201 72.084 65.233 72.148 ;
			RECT	65.369 72.084 65.401 72.148 ;
			RECT	65.537 72.084 65.569 72.148 ;
			RECT	65.705 72.084 65.737 72.148 ;
			RECT	65.873 72.084 65.905 72.148 ;
			RECT	66.041 72.084 66.073 72.148 ;
			RECT	66.209 72.084 66.241 72.148 ;
			RECT	66.377 72.084 66.409 72.148 ;
			RECT	66.545 72.084 66.577 72.148 ;
			RECT	66.713 72.084 66.745 72.148 ;
			RECT	66.881 72.084 66.913 72.148 ;
			RECT	67.049 72.084 67.081 72.148 ;
			RECT	67.217 72.084 67.249 72.148 ;
			RECT	67.385 72.084 67.417 72.148 ;
			RECT	67.553 72.084 67.585 72.148 ;
			RECT	67.721 72.084 67.753 72.148 ;
			RECT	67.889 72.084 67.921 72.148 ;
			RECT	68.057 72.084 68.089 72.148 ;
			RECT	68.225 72.084 68.257 72.148 ;
			RECT	68.393 72.084 68.425 72.148 ;
			RECT	68.561 72.084 68.593 72.148 ;
			RECT	68.729 72.084 68.761 72.148 ;
			RECT	68.897 72.084 68.929 72.148 ;
			RECT	69.065 72.084 69.097 72.148 ;
			RECT	69.233 72.084 69.265 72.148 ;
			RECT	69.401 72.084 69.433 72.148 ;
			RECT	69.569 72.084 69.601 72.148 ;
			RECT	69.737 72.084 69.769 72.148 ;
			RECT	69.905 72.084 69.937 72.148 ;
			RECT	70.073 72.084 70.105 72.148 ;
			RECT	70.241 72.084 70.273 72.148 ;
			RECT	70.409 72.084 70.441 72.148 ;
			RECT	70.577 72.084 70.609 72.148 ;
			RECT	70.745 72.084 70.777 72.148 ;
			RECT	70.913 72.084 70.945 72.148 ;
			RECT	71.081 72.084 71.113 72.148 ;
			RECT	71.249 72.084 71.281 72.148 ;
			RECT	71.417 72.084 71.449 72.148 ;
			RECT	71.585 72.084 71.617 72.148 ;
			RECT	71.753 72.084 71.785 72.148 ;
			RECT	71.921 72.084 71.953 72.148 ;
			RECT	72.089 72.084 72.121 72.148 ;
			RECT	72.257 72.084 72.289 72.148 ;
			RECT	72.425 72.084 72.457 72.148 ;
			RECT	72.593 72.084 72.625 72.148 ;
			RECT	72.761 72.084 72.793 72.148 ;
			RECT	72.929 72.084 72.961 72.148 ;
			RECT	73.097 72.084 73.129 72.148 ;
			RECT	73.265 72.084 73.297 72.148 ;
			RECT	73.433 72.084 73.465 72.148 ;
			RECT	73.601 72.084 73.633 72.148 ;
			RECT	73.769 72.084 73.801 72.148 ;
			RECT	73.937 72.084 73.969 72.148 ;
			RECT	74.105 72.084 74.137 72.148 ;
			RECT	74.273 72.084 74.305 72.148 ;
			RECT	74.441 72.084 74.473 72.148 ;
			RECT	74.609 72.084 74.641 72.148 ;
			RECT	74.777 72.084 74.809 72.148 ;
			RECT	74.945 72.084 74.977 72.148 ;
			RECT	75.113 72.084 75.145 72.148 ;
			RECT	75.281 72.084 75.313 72.148 ;
			RECT	75.449 72.084 75.481 72.148 ;
			RECT	75.617 72.084 75.649 72.148 ;
			RECT	75.785 72.084 75.817 72.148 ;
			RECT	75.953 72.084 75.985 72.148 ;
			RECT	76.121 72.084 76.153 72.148 ;
			RECT	76.289 72.084 76.321 72.148 ;
			RECT	76.457 72.084 76.489 72.148 ;
			RECT	76.625 72.084 76.657 72.148 ;
			RECT	76.793 72.084 76.825 72.148 ;
			RECT	76.961 72.084 76.993 72.148 ;
			RECT	77.129 72.084 77.161 72.148 ;
			RECT	77.297 72.084 77.329 72.148 ;
			RECT	77.465 72.084 77.497 72.148 ;
			RECT	77.633 72.084 77.665 72.148 ;
			RECT	77.801 72.084 77.833 72.148 ;
			RECT	77.969 72.084 78.001 72.148 ;
			RECT	78.137 72.084 78.169 72.148 ;
			RECT	78.305 72.084 78.337 72.148 ;
			RECT	78.473 72.084 78.505 72.148 ;
			RECT	78.641 72.084 78.673 72.148 ;
			RECT	78.809 72.084 78.841 72.148 ;
			RECT	78.977 72.084 79.009 72.148 ;
			RECT	79.145 72.084 79.177 72.148 ;
			RECT	79.313 72.084 79.345 72.148 ;
			RECT	79.481 72.084 79.513 72.148 ;
			RECT	79.649 72.084 79.681 72.148 ;
			RECT	79.817 72.084 79.849 72.148 ;
			RECT	79.985 72.084 80.017 72.148 ;
			RECT	80.153 72.084 80.185 72.148 ;
			RECT	80.321 72.084 80.353 72.148 ;
			RECT	80.489 72.084 80.521 72.148 ;
			RECT	80.657 72.084 80.689 72.148 ;
			RECT	80.825 72.084 80.857 72.148 ;
			RECT	80.993 72.084 81.025 72.148 ;
			RECT	81.161 72.084 81.193 72.148 ;
			RECT	81.329 72.084 81.361 72.148 ;
			RECT	81.497 72.084 81.529 72.148 ;
			RECT	81.665 72.084 81.697 72.148 ;
			RECT	81.833 72.084 81.865 72.148 ;
			RECT	82.001 72.084 82.033 72.148 ;
			RECT	82.169 72.084 82.201 72.148 ;
			RECT	82.337 72.084 82.369 72.148 ;
			RECT	82.505 72.084 82.537 72.148 ;
			RECT	82.673 72.084 82.705 72.148 ;
			RECT	82.841 72.084 82.873 72.148 ;
			RECT	83.009 72.084 83.041 72.148 ;
			RECT	83.177 72.084 83.209 72.148 ;
			RECT	83.345 72.084 83.377 72.148 ;
			RECT	83.513 72.084 83.545 72.148 ;
			RECT	83.681 72.084 83.713 72.148 ;
			RECT	83.849 72.084 83.881 72.148 ;
			RECT	84.017 72.084 84.049 72.148 ;
			RECT	84.185 72.084 84.217 72.148 ;
			RECT	84.353 72.084 84.385 72.148 ;
			RECT	84.521 72.084 84.553 72.148 ;
			RECT	84.689 72.084 84.721 72.148 ;
			RECT	84.857 72.084 84.889 72.148 ;
			RECT	85.025 72.084 85.057 72.148 ;
			RECT	85.193 72.084 85.225 72.148 ;
			RECT	85.361 72.084 85.393 72.148 ;
			RECT	85.529 72.084 85.561 72.148 ;
			RECT	85.697 72.084 85.729 72.148 ;
			RECT	85.865 72.084 85.897 72.148 ;
			RECT	86.033 72.084 86.065 72.148 ;
			RECT	86.201 72.084 86.233 72.148 ;
			RECT	86.369 72.084 86.401 72.148 ;
			RECT	86.537 72.084 86.569 72.148 ;
			RECT	86.705 72.084 86.737 72.148 ;
			RECT	86.873 72.084 86.905 72.148 ;
			RECT	87.041 72.084 87.073 72.148 ;
			RECT	87.209 72.084 87.241 72.148 ;
			RECT	87.377 72.084 87.409 72.148 ;
			RECT	87.545 72.084 87.577 72.148 ;
			RECT	87.713 72.084 87.745 72.148 ;
			RECT	87.881 72.084 87.913 72.148 ;
			RECT	88.049 72.084 88.081 72.148 ;
			RECT	88.217 72.084 88.249 72.148 ;
			RECT	88.385 72.084 88.417 72.148 ;
			RECT	88.553 72.084 88.585 72.148 ;
			RECT	88.721 72.084 88.753 72.148 ;
			RECT	88.889 72.084 88.921 72.148 ;
			RECT	89.057 72.084 89.089 72.148 ;
			RECT	89.225 72.084 89.257 72.148 ;
			RECT	89.393 72.084 89.425 72.148 ;
			RECT	89.561 72.084 89.593 72.148 ;
			RECT	89.729 72.084 89.761 72.148 ;
			RECT	89.897 72.084 89.929 72.148 ;
			RECT	90.065 72.084 90.097 72.148 ;
			RECT	90.233 72.084 90.265 72.148 ;
			RECT	90.401 72.084 90.433 72.148 ;
			RECT	90.569 72.084 90.601 72.148 ;
			RECT	90.737 72.084 90.769 72.148 ;
			RECT	90.905 72.084 90.937 72.148 ;
			RECT	91.073 72.084 91.105 72.148 ;
			RECT	91.241 72.084 91.273 72.148 ;
			RECT	91.409 72.084 91.441 72.148 ;
			RECT	91.577 72.084 91.609 72.148 ;
			RECT	91.745 72.084 91.777 72.148 ;
			RECT	91.913 72.084 91.945 72.148 ;
			RECT	92.081 72.084 92.113 72.148 ;
			RECT	92.249 72.084 92.281 72.148 ;
			RECT	92.417 72.084 92.449 72.148 ;
			RECT	92.585 72.084 92.617 72.148 ;
			RECT	92.753 72.084 92.785 72.148 ;
			RECT	92.921 72.084 92.953 72.148 ;
			RECT	93.089 72.084 93.121 72.148 ;
			RECT	93.257 72.084 93.289 72.148 ;
			RECT	93.425 72.084 93.457 72.148 ;
			RECT	93.593 72.084 93.625 72.148 ;
			RECT	93.761 72.084 93.793 72.148 ;
			RECT	93.929 72.084 93.961 72.148 ;
			RECT	94.097 72.084 94.129 72.148 ;
			RECT	94.265 72.084 94.297 72.148 ;
			RECT	94.433 72.084 94.465 72.148 ;
			RECT	94.601 72.084 94.633 72.148 ;
			RECT	94.769 72.084 94.801 72.148 ;
			RECT	94.937 72.084 94.969 72.148 ;
			RECT	95.105 72.084 95.137 72.148 ;
			RECT	95.273 72.084 95.305 72.148 ;
			RECT	95.441 72.084 95.473 72.148 ;
			RECT	95.609 72.084 95.641 72.148 ;
			RECT	95.777 72.084 95.809 72.148 ;
			RECT	95.945 72.084 95.977 72.148 ;
			RECT	96.113 72.084 96.145 72.148 ;
			RECT	96.281 72.084 96.313 72.148 ;
			RECT	96.449 72.084 96.481 72.148 ;
			RECT	96.617 72.084 96.649 72.148 ;
			RECT	96.785 72.084 96.817 72.148 ;
			RECT	96.953 72.084 96.985 72.148 ;
			RECT	97.121 72.084 97.153 72.148 ;
			RECT	97.289 72.084 97.321 72.148 ;
			RECT	97.457 72.084 97.489 72.148 ;
			RECT	97.625 72.084 97.657 72.148 ;
			RECT	97.793 72.084 97.825 72.148 ;
			RECT	97.961 72.084 97.993 72.148 ;
			RECT	98.129 72.084 98.161 72.148 ;
			RECT	98.297 72.084 98.329 72.148 ;
			RECT	98.465 72.084 98.497 72.148 ;
			RECT	98.633 72.084 98.665 72.148 ;
			RECT	98.801 72.084 98.833 72.148 ;
			RECT	98.969 72.084 99.001 72.148 ;
			RECT	99.137 72.084 99.169 72.148 ;
			RECT	99.305 72.084 99.337 72.148 ;
			RECT	99.473 72.084 99.505 72.148 ;
			RECT	99.641 72.084 99.673 72.148 ;
			RECT	99.809 72.084 99.841 72.148 ;
			RECT	99.977 72.084 100.009 72.148 ;
			RECT	100.145 72.084 100.177 72.148 ;
			RECT	100.313 72.084 100.345 72.148 ;
			RECT	100.481 72.084 100.513 72.148 ;
			RECT	100.649 72.084 100.681 72.148 ;
			RECT	100.817 72.084 100.849 72.148 ;
			RECT	100.985 72.084 101.017 72.148 ;
			RECT	101.153 72.084 101.185 72.148 ;
			RECT	101.321 72.084 101.353 72.148 ;
			RECT	101.489 72.084 101.521 72.148 ;
			RECT	101.657 72.084 101.689 72.148 ;
			RECT	101.825 72.084 101.857 72.148 ;
			RECT	101.993 72.084 102.025 72.148 ;
			RECT	102.123 72.1 102.155 72.132 ;
			RECT	102.245 72.095 102.277 72.127 ;
			RECT	102.375 72.084 102.407 72.148 ;
			RECT	103.795 72.084 103.827 72.148 ;
			RECT	103.925 72.095 103.957 72.127 ;
			RECT	104.047 72.1 104.079 72.132 ;
			RECT	104.177 72.084 104.209 72.148 ;
			RECT	104.345 72.084 104.377 72.148 ;
			RECT	104.513 72.084 104.545 72.148 ;
			RECT	104.681 72.084 104.713 72.148 ;
			RECT	104.849 72.084 104.881 72.148 ;
			RECT	105.017 72.084 105.049 72.148 ;
			RECT	105.185 72.084 105.217 72.148 ;
			RECT	105.353 72.084 105.385 72.148 ;
			RECT	105.521 72.084 105.553 72.148 ;
			RECT	105.689 72.084 105.721 72.148 ;
			RECT	105.857 72.084 105.889 72.148 ;
			RECT	106.025 72.084 106.057 72.148 ;
			RECT	106.193 72.084 106.225 72.148 ;
			RECT	106.361 72.084 106.393 72.148 ;
			RECT	106.529 72.084 106.561 72.148 ;
			RECT	106.697 72.084 106.729 72.148 ;
			RECT	106.865 72.084 106.897 72.148 ;
			RECT	107.033 72.084 107.065 72.148 ;
			RECT	107.201 72.084 107.233 72.148 ;
			RECT	107.369 72.084 107.401 72.148 ;
			RECT	107.537 72.084 107.569 72.148 ;
			RECT	107.705 72.084 107.737 72.148 ;
			RECT	107.873 72.084 107.905 72.148 ;
			RECT	108.041 72.084 108.073 72.148 ;
			RECT	108.209 72.084 108.241 72.148 ;
			RECT	108.377 72.084 108.409 72.148 ;
			RECT	108.545 72.084 108.577 72.148 ;
			RECT	108.713 72.084 108.745 72.148 ;
			RECT	108.881 72.084 108.913 72.148 ;
			RECT	109.049 72.084 109.081 72.148 ;
			RECT	109.217 72.084 109.249 72.148 ;
			RECT	109.385 72.084 109.417 72.148 ;
			RECT	109.553 72.084 109.585 72.148 ;
			RECT	109.721 72.084 109.753 72.148 ;
			RECT	109.889 72.084 109.921 72.148 ;
			RECT	110.057 72.084 110.089 72.148 ;
			RECT	110.225 72.084 110.257 72.148 ;
			RECT	110.393 72.084 110.425 72.148 ;
			RECT	110.561 72.084 110.593 72.148 ;
			RECT	110.729 72.084 110.761 72.148 ;
			RECT	110.897 72.084 110.929 72.148 ;
			RECT	111.065 72.084 111.097 72.148 ;
			RECT	111.233 72.084 111.265 72.148 ;
			RECT	111.401 72.084 111.433 72.148 ;
			RECT	111.569 72.084 111.601 72.148 ;
			RECT	111.737 72.084 111.769 72.148 ;
			RECT	111.905 72.084 111.937 72.148 ;
			RECT	112.073 72.084 112.105 72.148 ;
			RECT	112.241 72.084 112.273 72.148 ;
			RECT	112.409 72.084 112.441 72.148 ;
			RECT	112.577 72.084 112.609 72.148 ;
			RECT	112.745 72.084 112.777 72.148 ;
			RECT	112.913 72.084 112.945 72.148 ;
			RECT	113.081 72.084 113.113 72.148 ;
			RECT	113.249 72.084 113.281 72.148 ;
			RECT	113.417 72.084 113.449 72.148 ;
			RECT	113.585 72.084 113.617 72.148 ;
			RECT	113.753 72.084 113.785 72.148 ;
			RECT	113.921 72.084 113.953 72.148 ;
			RECT	114.089 72.084 114.121 72.148 ;
			RECT	114.257 72.084 114.289 72.148 ;
			RECT	114.425 72.084 114.457 72.148 ;
			RECT	114.593 72.084 114.625 72.148 ;
			RECT	114.761 72.084 114.793 72.148 ;
			RECT	114.929 72.084 114.961 72.148 ;
			RECT	115.097 72.084 115.129 72.148 ;
			RECT	115.265 72.084 115.297 72.148 ;
			RECT	115.433 72.084 115.465 72.148 ;
			RECT	115.601 72.084 115.633 72.148 ;
			RECT	115.769 72.084 115.801 72.148 ;
			RECT	115.937 72.084 115.969 72.148 ;
			RECT	116.105 72.084 116.137 72.148 ;
			RECT	116.273 72.084 116.305 72.148 ;
			RECT	116.441 72.084 116.473 72.148 ;
			RECT	116.609 72.084 116.641 72.148 ;
			RECT	116.777 72.084 116.809 72.148 ;
			RECT	116.945 72.084 116.977 72.148 ;
			RECT	117.113 72.084 117.145 72.148 ;
			RECT	117.281 72.084 117.313 72.148 ;
			RECT	117.449 72.084 117.481 72.148 ;
			RECT	117.617 72.084 117.649 72.148 ;
			RECT	117.785 72.084 117.817 72.148 ;
			RECT	117.953 72.084 117.985 72.148 ;
			RECT	118.121 72.084 118.153 72.148 ;
			RECT	118.289 72.084 118.321 72.148 ;
			RECT	118.457 72.084 118.489 72.148 ;
			RECT	118.625 72.084 118.657 72.148 ;
			RECT	118.793 72.084 118.825 72.148 ;
			RECT	118.961 72.084 118.993 72.148 ;
			RECT	119.129 72.084 119.161 72.148 ;
			RECT	119.297 72.084 119.329 72.148 ;
			RECT	119.465 72.084 119.497 72.148 ;
			RECT	119.633 72.084 119.665 72.148 ;
			RECT	119.801 72.084 119.833 72.148 ;
			RECT	119.969 72.084 120.001 72.148 ;
			RECT	120.137 72.084 120.169 72.148 ;
			RECT	120.305 72.084 120.337 72.148 ;
			RECT	120.473 72.084 120.505 72.148 ;
			RECT	120.641 72.084 120.673 72.148 ;
			RECT	120.809 72.084 120.841 72.148 ;
			RECT	120.977 72.084 121.009 72.148 ;
			RECT	121.145 72.084 121.177 72.148 ;
			RECT	121.313 72.084 121.345 72.148 ;
			RECT	121.481 72.084 121.513 72.148 ;
			RECT	121.649 72.084 121.681 72.148 ;
			RECT	121.817 72.084 121.849 72.148 ;
			RECT	121.985 72.084 122.017 72.148 ;
			RECT	122.153 72.084 122.185 72.148 ;
			RECT	122.321 72.084 122.353 72.148 ;
			RECT	122.489 72.084 122.521 72.148 ;
			RECT	122.657 72.084 122.689 72.148 ;
			RECT	122.825 72.084 122.857 72.148 ;
			RECT	122.993 72.084 123.025 72.148 ;
			RECT	123.161 72.084 123.193 72.148 ;
			RECT	123.329 72.084 123.361 72.148 ;
			RECT	123.497 72.084 123.529 72.148 ;
			RECT	123.665 72.084 123.697 72.148 ;
			RECT	123.833 72.084 123.865 72.148 ;
			RECT	124.001 72.084 124.033 72.148 ;
			RECT	124.169 72.084 124.201 72.148 ;
			RECT	124.337 72.084 124.369 72.148 ;
			RECT	124.505 72.084 124.537 72.148 ;
			RECT	124.673 72.084 124.705 72.148 ;
			RECT	124.841 72.084 124.873 72.148 ;
			RECT	125.009 72.084 125.041 72.148 ;
			RECT	125.177 72.084 125.209 72.148 ;
			RECT	125.345 72.084 125.377 72.148 ;
			RECT	125.513 72.084 125.545 72.148 ;
			RECT	125.681 72.084 125.713 72.148 ;
			RECT	125.849 72.084 125.881 72.148 ;
			RECT	126.017 72.084 126.049 72.148 ;
			RECT	126.185 72.084 126.217 72.148 ;
			RECT	126.353 72.084 126.385 72.148 ;
			RECT	126.521 72.084 126.553 72.148 ;
			RECT	126.689 72.084 126.721 72.148 ;
			RECT	126.857 72.084 126.889 72.148 ;
			RECT	127.025 72.084 127.057 72.148 ;
			RECT	127.193 72.084 127.225 72.148 ;
			RECT	127.361 72.084 127.393 72.148 ;
			RECT	127.529 72.084 127.561 72.148 ;
			RECT	127.697 72.084 127.729 72.148 ;
			RECT	127.865 72.084 127.897 72.148 ;
			RECT	128.033 72.084 128.065 72.148 ;
			RECT	128.201 72.084 128.233 72.148 ;
			RECT	128.369 72.084 128.401 72.148 ;
			RECT	128.537 72.084 128.569 72.148 ;
			RECT	128.705 72.084 128.737 72.148 ;
			RECT	128.873 72.084 128.905 72.148 ;
			RECT	129.041 72.084 129.073 72.148 ;
			RECT	129.209 72.084 129.241 72.148 ;
			RECT	129.377 72.084 129.409 72.148 ;
			RECT	129.545 72.084 129.577 72.148 ;
			RECT	129.713 72.084 129.745 72.148 ;
			RECT	129.881 72.084 129.913 72.148 ;
			RECT	130.049 72.084 130.081 72.148 ;
			RECT	130.217 72.084 130.249 72.148 ;
			RECT	130.385 72.084 130.417 72.148 ;
			RECT	130.553 72.084 130.585 72.148 ;
			RECT	130.721 72.084 130.753 72.148 ;
			RECT	130.889 72.084 130.921 72.148 ;
			RECT	131.057 72.084 131.089 72.148 ;
			RECT	131.225 72.084 131.257 72.148 ;
			RECT	131.393 72.084 131.425 72.148 ;
			RECT	131.561 72.084 131.593 72.148 ;
			RECT	131.729 72.084 131.761 72.148 ;
			RECT	131.897 72.084 131.929 72.148 ;
			RECT	132.065 72.084 132.097 72.148 ;
			RECT	132.233 72.084 132.265 72.148 ;
			RECT	132.401 72.084 132.433 72.148 ;
			RECT	132.569 72.084 132.601 72.148 ;
			RECT	132.737 72.084 132.769 72.148 ;
			RECT	132.905 72.084 132.937 72.148 ;
			RECT	133.073 72.084 133.105 72.148 ;
			RECT	133.241 72.084 133.273 72.148 ;
			RECT	133.409 72.084 133.441 72.148 ;
			RECT	133.577 72.084 133.609 72.148 ;
			RECT	133.745 72.084 133.777 72.148 ;
			RECT	133.913 72.084 133.945 72.148 ;
			RECT	134.081 72.084 134.113 72.148 ;
			RECT	134.249 72.084 134.281 72.148 ;
			RECT	134.417 72.084 134.449 72.148 ;
			RECT	134.585 72.084 134.617 72.148 ;
			RECT	134.753 72.084 134.785 72.148 ;
			RECT	134.921 72.084 134.953 72.148 ;
			RECT	135.089 72.084 135.121 72.148 ;
			RECT	135.257 72.084 135.289 72.148 ;
			RECT	135.425 72.084 135.457 72.148 ;
			RECT	135.593 72.084 135.625 72.148 ;
			RECT	135.761 72.084 135.793 72.148 ;
			RECT	135.929 72.084 135.961 72.148 ;
			RECT	136.097 72.084 136.129 72.148 ;
			RECT	136.265 72.084 136.297 72.148 ;
			RECT	136.433 72.084 136.465 72.148 ;
			RECT	136.601 72.084 136.633 72.148 ;
			RECT	136.769 72.084 136.801 72.148 ;
			RECT	136.937 72.084 136.969 72.148 ;
			RECT	137.105 72.084 137.137 72.148 ;
			RECT	137.273 72.084 137.305 72.148 ;
			RECT	137.441 72.084 137.473 72.148 ;
			RECT	137.609 72.084 137.641 72.148 ;
			RECT	137.777 72.084 137.809 72.148 ;
			RECT	137.945 72.084 137.977 72.148 ;
			RECT	138.113 72.084 138.145 72.148 ;
			RECT	138.281 72.084 138.313 72.148 ;
			RECT	138.449 72.084 138.481 72.148 ;
			RECT	138.617 72.084 138.649 72.148 ;
			RECT	138.785 72.084 138.817 72.148 ;
			RECT	138.953 72.084 138.985 72.148 ;
			RECT	139.121 72.084 139.153 72.148 ;
			RECT	139.289 72.084 139.321 72.148 ;
			RECT	139.457 72.084 139.489 72.148 ;
			RECT	139.625 72.084 139.657 72.148 ;
			RECT	139.793 72.084 139.825 72.148 ;
			RECT	139.961 72.084 139.993 72.148 ;
			RECT	140.129 72.084 140.161 72.148 ;
			RECT	140.297 72.084 140.329 72.148 ;
			RECT	140.465 72.084 140.497 72.148 ;
			RECT	140.633 72.084 140.665 72.148 ;
			RECT	140.801 72.084 140.833 72.148 ;
			RECT	140.969 72.084 141.001 72.148 ;
			RECT	141.137 72.084 141.169 72.148 ;
			RECT	141.305 72.084 141.337 72.148 ;
			RECT	141.473 72.084 141.505 72.148 ;
			RECT	141.641 72.084 141.673 72.148 ;
			RECT	141.809 72.084 141.841 72.148 ;
			RECT	141.977 72.084 142.009 72.148 ;
			RECT	142.145 72.084 142.177 72.148 ;
			RECT	142.313 72.084 142.345 72.148 ;
			RECT	142.481 72.084 142.513 72.148 ;
			RECT	142.649 72.084 142.681 72.148 ;
			RECT	142.817 72.084 142.849 72.148 ;
			RECT	142.985 72.084 143.017 72.148 ;
			RECT	143.153 72.084 143.185 72.148 ;
			RECT	143.321 72.084 143.353 72.148 ;
			RECT	143.489 72.084 143.521 72.148 ;
			RECT	143.657 72.084 143.689 72.148 ;
			RECT	143.825 72.084 143.857 72.148 ;
			RECT	143.993 72.084 144.025 72.148 ;
			RECT	144.161 72.084 144.193 72.148 ;
			RECT	144.329 72.084 144.361 72.148 ;
			RECT	144.497 72.084 144.529 72.148 ;
			RECT	144.665 72.084 144.697 72.148 ;
			RECT	144.833 72.084 144.865 72.148 ;
			RECT	145.001 72.084 145.033 72.148 ;
			RECT	145.169 72.084 145.201 72.148 ;
			RECT	145.337 72.084 145.369 72.148 ;
			RECT	145.505 72.084 145.537 72.148 ;
			RECT	145.673 72.084 145.705 72.148 ;
			RECT	145.841 72.084 145.873 72.148 ;
			RECT	146.009 72.084 146.041 72.148 ;
			RECT	146.177 72.084 146.209 72.148 ;
			RECT	146.345 72.084 146.377 72.148 ;
			RECT	146.513 72.084 146.545 72.148 ;
			RECT	146.681 72.084 146.713 72.148 ;
			RECT	146.849 72.084 146.881 72.148 ;
			RECT	147.017 72.084 147.049 72.148 ;
			RECT	147.185 72.084 147.217 72.148 ;
			RECT	147.316 72.1 147.348 72.132 ;
			RECT	147.437 72.1 147.469 72.132 ;
			RECT	147.567 72.084 147.599 72.148 ;
			RECT	149.879 72.084 149.911 72.148 ;
			RECT	151.13 72.084 151.194 72.148 ;
			RECT	151.81 72.084 151.842 72.148 ;
			RECT	152.249 72.084 152.281 72.148 ;
			RECT	153.56 72.084 153.624 72.148 ;
			RECT	156.601 72.084 156.633 72.148 ;
			RECT	156.731 72.1 156.763 72.132 ;
			RECT	156.852 72.1 156.884 72.132 ;
			RECT	156.983 72.084 157.015 72.148 ;
			RECT	157.151 72.084 157.183 72.148 ;
			RECT	157.319 72.084 157.351 72.148 ;
			RECT	157.487 72.084 157.519 72.148 ;
			RECT	157.655 72.084 157.687 72.148 ;
			RECT	157.823 72.084 157.855 72.148 ;
			RECT	157.991 72.084 158.023 72.148 ;
			RECT	158.159 72.084 158.191 72.148 ;
			RECT	158.327 72.084 158.359 72.148 ;
			RECT	158.495 72.084 158.527 72.148 ;
			RECT	158.663 72.084 158.695 72.148 ;
			RECT	158.831 72.084 158.863 72.148 ;
			RECT	158.999 72.084 159.031 72.148 ;
			RECT	159.167 72.084 159.199 72.148 ;
			RECT	159.335 72.084 159.367 72.148 ;
			RECT	159.503 72.084 159.535 72.148 ;
			RECT	159.671 72.084 159.703 72.148 ;
			RECT	159.839 72.084 159.871 72.148 ;
			RECT	160.007 72.084 160.039 72.148 ;
			RECT	160.175 72.084 160.207 72.148 ;
			RECT	160.343 72.084 160.375 72.148 ;
			RECT	160.511 72.084 160.543 72.148 ;
			RECT	160.679 72.084 160.711 72.148 ;
			RECT	160.847 72.084 160.879 72.148 ;
			RECT	161.015 72.084 161.047 72.148 ;
			RECT	161.183 72.084 161.215 72.148 ;
			RECT	161.351 72.084 161.383 72.148 ;
			RECT	161.519 72.084 161.551 72.148 ;
			RECT	161.687 72.084 161.719 72.148 ;
			RECT	161.855 72.084 161.887 72.148 ;
			RECT	162.023 72.084 162.055 72.148 ;
			RECT	162.191 72.084 162.223 72.148 ;
			RECT	162.359 72.084 162.391 72.148 ;
			RECT	162.527 72.084 162.559 72.148 ;
			RECT	162.695 72.084 162.727 72.148 ;
			RECT	162.863 72.084 162.895 72.148 ;
			RECT	163.031 72.084 163.063 72.148 ;
			RECT	163.199 72.084 163.231 72.148 ;
			RECT	163.367 72.084 163.399 72.148 ;
			RECT	163.535 72.084 163.567 72.148 ;
			RECT	163.703 72.084 163.735 72.148 ;
			RECT	163.871 72.084 163.903 72.148 ;
			RECT	164.039 72.084 164.071 72.148 ;
			RECT	164.207 72.084 164.239 72.148 ;
			RECT	164.375 72.084 164.407 72.148 ;
			RECT	164.543 72.084 164.575 72.148 ;
			RECT	164.711 72.084 164.743 72.148 ;
			RECT	164.879 72.084 164.911 72.148 ;
			RECT	165.047 72.084 165.079 72.148 ;
			RECT	165.215 72.084 165.247 72.148 ;
			RECT	165.383 72.084 165.415 72.148 ;
			RECT	165.551 72.084 165.583 72.148 ;
			RECT	165.719 72.084 165.751 72.148 ;
			RECT	165.887 72.084 165.919 72.148 ;
			RECT	166.055 72.084 166.087 72.148 ;
			RECT	166.223 72.084 166.255 72.148 ;
			RECT	166.391 72.084 166.423 72.148 ;
			RECT	166.559 72.084 166.591 72.148 ;
			RECT	166.727 72.084 166.759 72.148 ;
			RECT	166.895 72.084 166.927 72.148 ;
			RECT	167.063 72.084 167.095 72.148 ;
			RECT	167.231 72.084 167.263 72.148 ;
			RECT	167.399 72.084 167.431 72.148 ;
			RECT	167.567 72.084 167.599 72.148 ;
			RECT	167.735 72.084 167.767 72.148 ;
			RECT	167.903 72.084 167.935 72.148 ;
			RECT	168.071 72.084 168.103 72.148 ;
			RECT	168.239 72.084 168.271 72.148 ;
			RECT	168.407 72.084 168.439 72.148 ;
			RECT	168.575 72.084 168.607 72.148 ;
			RECT	168.743 72.084 168.775 72.148 ;
			RECT	168.911 72.084 168.943 72.148 ;
			RECT	169.079 72.084 169.111 72.148 ;
			RECT	169.247 72.084 169.279 72.148 ;
			RECT	169.415 72.084 169.447 72.148 ;
			RECT	169.583 72.084 169.615 72.148 ;
			RECT	169.751 72.084 169.783 72.148 ;
			RECT	169.919 72.084 169.951 72.148 ;
			RECT	170.087 72.084 170.119 72.148 ;
			RECT	170.255 72.084 170.287 72.148 ;
			RECT	170.423 72.084 170.455 72.148 ;
			RECT	170.591 72.084 170.623 72.148 ;
			RECT	170.759 72.084 170.791 72.148 ;
			RECT	170.927 72.084 170.959 72.148 ;
			RECT	171.095 72.084 171.127 72.148 ;
			RECT	171.263 72.084 171.295 72.148 ;
			RECT	171.431 72.084 171.463 72.148 ;
			RECT	171.599 72.084 171.631 72.148 ;
			RECT	171.767 72.084 171.799 72.148 ;
			RECT	171.935 72.084 171.967 72.148 ;
			RECT	172.103 72.084 172.135 72.148 ;
			RECT	172.271 72.084 172.303 72.148 ;
			RECT	172.439 72.084 172.471 72.148 ;
			RECT	172.607 72.084 172.639 72.148 ;
			RECT	172.775 72.084 172.807 72.148 ;
			RECT	172.943 72.084 172.975 72.148 ;
			RECT	173.111 72.084 173.143 72.148 ;
			RECT	173.279 72.084 173.311 72.148 ;
			RECT	173.447 72.084 173.479 72.148 ;
			RECT	173.615 72.084 173.647 72.148 ;
			RECT	173.783 72.084 173.815 72.148 ;
			RECT	173.951 72.084 173.983 72.148 ;
			RECT	174.119 72.084 174.151 72.148 ;
			RECT	174.287 72.084 174.319 72.148 ;
			RECT	174.455 72.084 174.487 72.148 ;
			RECT	174.623 72.084 174.655 72.148 ;
			RECT	174.791 72.084 174.823 72.148 ;
			RECT	174.959 72.084 174.991 72.148 ;
			RECT	175.127 72.084 175.159 72.148 ;
			RECT	175.295 72.084 175.327 72.148 ;
			RECT	175.463 72.084 175.495 72.148 ;
			RECT	175.631 72.084 175.663 72.148 ;
			RECT	175.799 72.084 175.831 72.148 ;
			RECT	175.967 72.084 175.999 72.148 ;
			RECT	176.135 72.084 176.167 72.148 ;
			RECT	176.303 72.084 176.335 72.148 ;
			RECT	176.471 72.084 176.503 72.148 ;
			RECT	176.639 72.084 176.671 72.148 ;
			RECT	176.807 72.084 176.839 72.148 ;
			RECT	176.975 72.084 177.007 72.148 ;
			RECT	177.143 72.084 177.175 72.148 ;
			RECT	177.311 72.084 177.343 72.148 ;
			RECT	177.479 72.084 177.511 72.148 ;
			RECT	177.647 72.084 177.679 72.148 ;
			RECT	177.815 72.084 177.847 72.148 ;
			RECT	177.983 72.084 178.015 72.148 ;
			RECT	178.151 72.084 178.183 72.148 ;
			RECT	178.319 72.084 178.351 72.148 ;
			RECT	178.487 72.084 178.519 72.148 ;
			RECT	178.655 72.084 178.687 72.148 ;
			RECT	178.823 72.084 178.855 72.148 ;
			RECT	178.991 72.084 179.023 72.148 ;
			RECT	179.159 72.084 179.191 72.148 ;
			RECT	179.327 72.084 179.359 72.148 ;
			RECT	179.495 72.084 179.527 72.148 ;
			RECT	179.663 72.084 179.695 72.148 ;
			RECT	179.831 72.084 179.863 72.148 ;
			RECT	179.999 72.084 180.031 72.148 ;
			RECT	180.167 72.084 180.199 72.148 ;
			RECT	180.335 72.084 180.367 72.148 ;
			RECT	180.503 72.084 180.535 72.148 ;
			RECT	180.671 72.084 180.703 72.148 ;
			RECT	180.839 72.084 180.871 72.148 ;
			RECT	181.007 72.084 181.039 72.148 ;
			RECT	181.175 72.084 181.207 72.148 ;
			RECT	181.343 72.084 181.375 72.148 ;
			RECT	181.511 72.084 181.543 72.148 ;
			RECT	181.679 72.084 181.711 72.148 ;
			RECT	181.847 72.084 181.879 72.148 ;
			RECT	182.015 72.084 182.047 72.148 ;
			RECT	182.183 72.084 182.215 72.148 ;
			RECT	182.351 72.084 182.383 72.148 ;
			RECT	182.519 72.084 182.551 72.148 ;
			RECT	182.687 72.084 182.719 72.148 ;
			RECT	182.855 72.084 182.887 72.148 ;
			RECT	183.023 72.084 183.055 72.148 ;
			RECT	183.191 72.084 183.223 72.148 ;
			RECT	183.359 72.084 183.391 72.148 ;
			RECT	183.527 72.084 183.559 72.148 ;
			RECT	183.695 72.084 183.727 72.148 ;
			RECT	183.863 72.084 183.895 72.148 ;
			RECT	184.031 72.084 184.063 72.148 ;
			RECT	184.199 72.084 184.231 72.148 ;
			RECT	184.367 72.084 184.399 72.148 ;
			RECT	184.535 72.084 184.567 72.148 ;
			RECT	184.703 72.084 184.735 72.148 ;
			RECT	184.871 72.084 184.903 72.148 ;
			RECT	185.039 72.084 185.071 72.148 ;
			RECT	185.207 72.084 185.239 72.148 ;
			RECT	185.375 72.084 185.407 72.148 ;
			RECT	185.543 72.084 185.575 72.148 ;
			RECT	185.711 72.084 185.743 72.148 ;
			RECT	185.879 72.084 185.911 72.148 ;
			RECT	186.047 72.084 186.079 72.148 ;
			RECT	186.215 72.084 186.247 72.148 ;
			RECT	186.383 72.084 186.415 72.148 ;
			RECT	186.551 72.084 186.583 72.148 ;
			RECT	186.719 72.084 186.751 72.148 ;
			RECT	186.887 72.084 186.919 72.148 ;
			RECT	187.055 72.084 187.087 72.148 ;
			RECT	187.223 72.084 187.255 72.148 ;
			RECT	187.391 72.084 187.423 72.148 ;
			RECT	187.559 72.084 187.591 72.148 ;
			RECT	187.727 72.084 187.759 72.148 ;
			RECT	187.895 72.084 187.927 72.148 ;
			RECT	188.063 72.084 188.095 72.148 ;
			RECT	188.231 72.084 188.263 72.148 ;
			RECT	188.399 72.084 188.431 72.148 ;
			RECT	188.567 72.084 188.599 72.148 ;
			RECT	188.735 72.084 188.767 72.148 ;
			RECT	188.903 72.084 188.935 72.148 ;
			RECT	189.071 72.084 189.103 72.148 ;
			RECT	189.239 72.084 189.271 72.148 ;
			RECT	189.407 72.084 189.439 72.148 ;
			RECT	189.575 72.084 189.607 72.148 ;
			RECT	189.743 72.084 189.775 72.148 ;
			RECT	189.911 72.084 189.943 72.148 ;
			RECT	190.079 72.084 190.111 72.148 ;
			RECT	190.247 72.084 190.279 72.148 ;
			RECT	190.415 72.084 190.447 72.148 ;
			RECT	190.583 72.084 190.615 72.148 ;
			RECT	190.751 72.084 190.783 72.148 ;
			RECT	190.919 72.084 190.951 72.148 ;
			RECT	191.087 72.084 191.119 72.148 ;
			RECT	191.255 72.084 191.287 72.148 ;
			RECT	191.423 72.084 191.455 72.148 ;
			RECT	191.591 72.084 191.623 72.148 ;
			RECT	191.759 72.084 191.791 72.148 ;
			RECT	191.927 72.084 191.959 72.148 ;
			RECT	192.095 72.084 192.127 72.148 ;
			RECT	192.263 72.084 192.295 72.148 ;
			RECT	192.431 72.084 192.463 72.148 ;
			RECT	192.599 72.084 192.631 72.148 ;
			RECT	192.767 72.084 192.799 72.148 ;
			RECT	192.935 72.084 192.967 72.148 ;
			RECT	193.103 72.084 193.135 72.148 ;
			RECT	193.271 72.084 193.303 72.148 ;
			RECT	193.439 72.084 193.471 72.148 ;
			RECT	193.607 72.084 193.639 72.148 ;
			RECT	193.775 72.084 193.807 72.148 ;
			RECT	193.943 72.084 193.975 72.148 ;
			RECT	194.111 72.084 194.143 72.148 ;
			RECT	194.279 72.084 194.311 72.148 ;
			RECT	194.447 72.084 194.479 72.148 ;
			RECT	194.615 72.084 194.647 72.148 ;
			RECT	194.783 72.084 194.815 72.148 ;
			RECT	194.951 72.084 194.983 72.148 ;
			RECT	195.119 72.084 195.151 72.148 ;
			RECT	195.287 72.084 195.319 72.148 ;
			RECT	195.455 72.084 195.487 72.148 ;
			RECT	195.623 72.084 195.655 72.148 ;
			RECT	195.791 72.084 195.823 72.148 ;
			RECT	195.959 72.084 195.991 72.148 ;
			RECT	196.127 72.084 196.159 72.148 ;
			RECT	196.295 72.084 196.327 72.148 ;
			RECT	196.463 72.084 196.495 72.148 ;
			RECT	196.631 72.084 196.663 72.148 ;
			RECT	196.799 72.084 196.831 72.148 ;
			RECT	196.967 72.084 196.999 72.148 ;
			RECT	197.135 72.084 197.167 72.148 ;
			RECT	197.303 72.084 197.335 72.148 ;
			RECT	197.471 72.084 197.503 72.148 ;
			RECT	197.639 72.084 197.671 72.148 ;
			RECT	197.807 72.084 197.839 72.148 ;
			RECT	197.975 72.084 198.007 72.148 ;
			RECT	198.143 72.084 198.175 72.148 ;
			RECT	198.311 72.084 198.343 72.148 ;
			RECT	198.479 72.084 198.511 72.148 ;
			RECT	198.647 72.084 198.679 72.148 ;
			RECT	198.815 72.084 198.847 72.148 ;
			RECT	198.983 72.084 199.015 72.148 ;
			RECT	199.151 72.084 199.183 72.148 ;
			RECT	199.319 72.084 199.351 72.148 ;
			RECT	199.487 72.084 199.519 72.148 ;
			RECT	199.655 72.084 199.687 72.148 ;
			RECT	199.823 72.084 199.855 72.148 ;
			RECT	199.991 72.084 200.023 72.148 ;
			RECT	200.121 72.1 200.153 72.132 ;
			RECT	200.243 72.095 200.275 72.127 ;
			RECT	200.373 72.084 200.405 72.148 ;
			RECT	200.9 72.084 200.932 72.148 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 70.136 201.665 70.256 ;
			LAYER	J3 ;
			RECT	0.755 70.164 0.787 70.228 ;
			RECT	1.645 70.164 1.709 70.228 ;
			RECT	2.323 70.164 2.387 70.228 ;
			RECT	3.438 70.164 3.47 70.228 ;
			RECT	3.585 70.164 3.617 70.228 ;
			RECT	4.195 70.164 4.227 70.228 ;
			RECT	4.72 70.164 4.752 70.228 ;
			RECT	4.944 70.164 5.008 70.228 ;
			RECT	5.267 70.164 5.299 70.228 ;
			RECT	5.797 70.164 5.829 70.228 ;
			RECT	5.927 70.175 5.959 70.207 ;
			RECT	6.049 70.18 6.081 70.212 ;
			RECT	6.179 70.164 6.211 70.228 ;
			RECT	6.347 70.164 6.379 70.228 ;
			RECT	6.515 70.164 6.547 70.228 ;
			RECT	6.683 70.164 6.715 70.228 ;
			RECT	6.851 70.164 6.883 70.228 ;
			RECT	7.019 70.164 7.051 70.228 ;
			RECT	7.187 70.164 7.219 70.228 ;
			RECT	7.355 70.164 7.387 70.228 ;
			RECT	7.523 70.164 7.555 70.228 ;
			RECT	7.691 70.164 7.723 70.228 ;
			RECT	7.859 70.164 7.891 70.228 ;
			RECT	8.027 70.164 8.059 70.228 ;
			RECT	8.195 70.164 8.227 70.228 ;
			RECT	8.363 70.164 8.395 70.228 ;
			RECT	8.531 70.164 8.563 70.228 ;
			RECT	8.699 70.164 8.731 70.228 ;
			RECT	8.867 70.164 8.899 70.228 ;
			RECT	9.035 70.164 9.067 70.228 ;
			RECT	9.203 70.164 9.235 70.228 ;
			RECT	9.371 70.164 9.403 70.228 ;
			RECT	9.539 70.164 9.571 70.228 ;
			RECT	9.707 70.164 9.739 70.228 ;
			RECT	9.875 70.164 9.907 70.228 ;
			RECT	10.043 70.164 10.075 70.228 ;
			RECT	10.211 70.164 10.243 70.228 ;
			RECT	10.379 70.164 10.411 70.228 ;
			RECT	10.547 70.164 10.579 70.228 ;
			RECT	10.715 70.164 10.747 70.228 ;
			RECT	10.883 70.164 10.915 70.228 ;
			RECT	11.051 70.164 11.083 70.228 ;
			RECT	11.219 70.164 11.251 70.228 ;
			RECT	11.387 70.164 11.419 70.228 ;
			RECT	11.555 70.164 11.587 70.228 ;
			RECT	11.723 70.164 11.755 70.228 ;
			RECT	11.891 70.164 11.923 70.228 ;
			RECT	12.059 70.164 12.091 70.228 ;
			RECT	12.227 70.164 12.259 70.228 ;
			RECT	12.395 70.164 12.427 70.228 ;
			RECT	12.563 70.164 12.595 70.228 ;
			RECT	12.731 70.164 12.763 70.228 ;
			RECT	12.899 70.164 12.931 70.228 ;
			RECT	13.067 70.164 13.099 70.228 ;
			RECT	13.235 70.164 13.267 70.228 ;
			RECT	13.403 70.164 13.435 70.228 ;
			RECT	13.571 70.164 13.603 70.228 ;
			RECT	13.739 70.164 13.771 70.228 ;
			RECT	13.907 70.164 13.939 70.228 ;
			RECT	14.075 70.164 14.107 70.228 ;
			RECT	14.243 70.164 14.275 70.228 ;
			RECT	14.411 70.164 14.443 70.228 ;
			RECT	14.579 70.164 14.611 70.228 ;
			RECT	14.747 70.164 14.779 70.228 ;
			RECT	14.915 70.164 14.947 70.228 ;
			RECT	15.083 70.164 15.115 70.228 ;
			RECT	15.251 70.164 15.283 70.228 ;
			RECT	15.419 70.164 15.451 70.228 ;
			RECT	15.587 70.164 15.619 70.228 ;
			RECT	15.755 70.164 15.787 70.228 ;
			RECT	15.923 70.164 15.955 70.228 ;
			RECT	16.091 70.164 16.123 70.228 ;
			RECT	16.259 70.164 16.291 70.228 ;
			RECT	16.427 70.164 16.459 70.228 ;
			RECT	16.595 70.164 16.627 70.228 ;
			RECT	16.763 70.164 16.795 70.228 ;
			RECT	16.931 70.164 16.963 70.228 ;
			RECT	17.099 70.164 17.131 70.228 ;
			RECT	17.267 70.164 17.299 70.228 ;
			RECT	17.435 70.164 17.467 70.228 ;
			RECT	17.603 70.164 17.635 70.228 ;
			RECT	17.771 70.164 17.803 70.228 ;
			RECT	17.939 70.164 17.971 70.228 ;
			RECT	18.107 70.164 18.139 70.228 ;
			RECT	18.275 70.164 18.307 70.228 ;
			RECT	18.443 70.164 18.475 70.228 ;
			RECT	18.611 70.164 18.643 70.228 ;
			RECT	18.779 70.164 18.811 70.228 ;
			RECT	18.947 70.164 18.979 70.228 ;
			RECT	19.115 70.164 19.147 70.228 ;
			RECT	19.283 70.164 19.315 70.228 ;
			RECT	19.451 70.164 19.483 70.228 ;
			RECT	19.619 70.164 19.651 70.228 ;
			RECT	19.787 70.164 19.819 70.228 ;
			RECT	19.955 70.164 19.987 70.228 ;
			RECT	20.123 70.164 20.155 70.228 ;
			RECT	20.291 70.164 20.323 70.228 ;
			RECT	20.459 70.164 20.491 70.228 ;
			RECT	20.627 70.164 20.659 70.228 ;
			RECT	20.795 70.164 20.827 70.228 ;
			RECT	20.963 70.164 20.995 70.228 ;
			RECT	21.131 70.164 21.163 70.228 ;
			RECT	21.299 70.164 21.331 70.228 ;
			RECT	21.467 70.164 21.499 70.228 ;
			RECT	21.635 70.164 21.667 70.228 ;
			RECT	21.803 70.164 21.835 70.228 ;
			RECT	21.971 70.164 22.003 70.228 ;
			RECT	22.139 70.164 22.171 70.228 ;
			RECT	22.307 70.164 22.339 70.228 ;
			RECT	22.475 70.164 22.507 70.228 ;
			RECT	22.643 70.164 22.675 70.228 ;
			RECT	22.811 70.164 22.843 70.228 ;
			RECT	22.979 70.164 23.011 70.228 ;
			RECT	23.147 70.164 23.179 70.228 ;
			RECT	23.315 70.164 23.347 70.228 ;
			RECT	23.483 70.164 23.515 70.228 ;
			RECT	23.651 70.164 23.683 70.228 ;
			RECT	23.819 70.164 23.851 70.228 ;
			RECT	23.987 70.164 24.019 70.228 ;
			RECT	24.155 70.164 24.187 70.228 ;
			RECT	24.323 70.164 24.355 70.228 ;
			RECT	24.491 70.164 24.523 70.228 ;
			RECT	24.659 70.164 24.691 70.228 ;
			RECT	24.827 70.164 24.859 70.228 ;
			RECT	24.995 70.164 25.027 70.228 ;
			RECT	25.163 70.164 25.195 70.228 ;
			RECT	25.331 70.164 25.363 70.228 ;
			RECT	25.499 70.164 25.531 70.228 ;
			RECT	25.667 70.164 25.699 70.228 ;
			RECT	25.835 70.164 25.867 70.228 ;
			RECT	26.003 70.164 26.035 70.228 ;
			RECT	26.171 70.164 26.203 70.228 ;
			RECT	26.339 70.164 26.371 70.228 ;
			RECT	26.507 70.164 26.539 70.228 ;
			RECT	26.675 70.164 26.707 70.228 ;
			RECT	26.843 70.164 26.875 70.228 ;
			RECT	27.011 70.164 27.043 70.228 ;
			RECT	27.179 70.164 27.211 70.228 ;
			RECT	27.347 70.164 27.379 70.228 ;
			RECT	27.515 70.164 27.547 70.228 ;
			RECT	27.683 70.164 27.715 70.228 ;
			RECT	27.851 70.164 27.883 70.228 ;
			RECT	28.019 70.164 28.051 70.228 ;
			RECT	28.187 70.164 28.219 70.228 ;
			RECT	28.355 70.164 28.387 70.228 ;
			RECT	28.523 70.164 28.555 70.228 ;
			RECT	28.691 70.164 28.723 70.228 ;
			RECT	28.859 70.164 28.891 70.228 ;
			RECT	29.027 70.164 29.059 70.228 ;
			RECT	29.195 70.164 29.227 70.228 ;
			RECT	29.363 70.164 29.395 70.228 ;
			RECT	29.531 70.164 29.563 70.228 ;
			RECT	29.699 70.164 29.731 70.228 ;
			RECT	29.867 70.164 29.899 70.228 ;
			RECT	30.035 70.164 30.067 70.228 ;
			RECT	30.203 70.164 30.235 70.228 ;
			RECT	30.371 70.164 30.403 70.228 ;
			RECT	30.539 70.164 30.571 70.228 ;
			RECT	30.707 70.164 30.739 70.228 ;
			RECT	30.875 70.164 30.907 70.228 ;
			RECT	31.043 70.164 31.075 70.228 ;
			RECT	31.211 70.164 31.243 70.228 ;
			RECT	31.379 70.164 31.411 70.228 ;
			RECT	31.547 70.164 31.579 70.228 ;
			RECT	31.715 70.164 31.747 70.228 ;
			RECT	31.883 70.164 31.915 70.228 ;
			RECT	32.051 70.164 32.083 70.228 ;
			RECT	32.219 70.164 32.251 70.228 ;
			RECT	32.387 70.164 32.419 70.228 ;
			RECT	32.555 70.164 32.587 70.228 ;
			RECT	32.723 70.164 32.755 70.228 ;
			RECT	32.891 70.164 32.923 70.228 ;
			RECT	33.059 70.164 33.091 70.228 ;
			RECT	33.227 70.164 33.259 70.228 ;
			RECT	33.395 70.164 33.427 70.228 ;
			RECT	33.563 70.164 33.595 70.228 ;
			RECT	33.731 70.164 33.763 70.228 ;
			RECT	33.899 70.164 33.931 70.228 ;
			RECT	34.067 70.164 34.099 70.228 ;
			RECT	34.235 70.164 34.267 70.228 ;
			RECT	34.403 70.164 34.435 70.228 ;
			RECT	34.571 70.164 34.603 70.228 ;
			RECT	34.739 70.164 34.771 70.228 ;
			RECT	34.907 70.164 34.939 70.228 ;
			RECT	35.075 70.164 35.107 70.228 ;
			RECT	35.243 70.164 35.275 70.228 ;
			RECT	35.411 70.164 35.443 70.228 ;
			RECT	35.579 70.164 35.611 70.228 ;
			RECT	35.747 70.164 35.779 70.228 ;
			RECT	35.915 70.164 35.947 70.228 ;
			RECT	36.083 70.164 36.115 70.228 ;
			RECT	36.251 70.164 36.283 70.228 ;
			RECT	36.419 70.164 36.451 70.228 ;
			RECT	36.587 70.164 36.619 70.228 ;
			RECT	36.755 70.164 36.787 70.228 ;
			RECT	36.923 70.164 36.955 70.228 ;
			RECT	37.091 70.164 37.123 70.228 ;
			RECT	37.259 70.164 37.291 70.228 ;
			RECT	37.427 70.164 37.459 70.228 ;
			RECT	37.595 70.164 37.627 70.228 ;
			RECT	37.763 70.164 37.795 70.228 ;
			RECT	37.931 70.164 37.963 70.228 ;
			RECT	38.099 70.164 38.131 70.228 ;
			RECT	38.267 70.164 38.299 70.228 ;
			RECT	38.435 70.164 38.467 70.228 ;
			RECT	38.603 70.164 38.635 70.228 ;
			RECT	38.771 70.164 38.803 70.228 ;
			RECT	38.939 70.164 38.971 70.228 ;
			RECT	39.107 70.164 39.139 70.228 ;
			RECT	39.275 70.164 39.307 70.228 ;
			RECT	39.443 70.164 39.475 70.228 ;
			RECT	39.611 70.164 39.643 70.228 ;
			RECT	39.779 70.164 39.811 70.228 ;
			RECT	39.947 70.164 39.979 70.228 ;
			RECT	40.115 70.164 40.147 70.228 ;
			RECT	40.283 70.164 40.315 70.228 ;
			RECT	40.451 70.164 40.483 70.228 ;
			RECT	40.619 70.164 40.651 70.228 ;
			RECT	40.787 70.164 40.819 70.228 ;
			RECT	40.955 70.164 40.987 70.228 ;
			RECT	41.123 70.164 41.155 70.228 ;
			RECT	41.291 70.164 41.323 70.228 ;
			RECT	41.459 70.164 41.491 70.228 ;
			RECT	41.627 70.164 41.659 70.228 ;
			RECT	41.795 70.164 41.827 70.228 ;
			RECT	41.963 70.164 41.995 70.228 ;
			RECT	42.131 70.164 42.163 70.228 ;
			RECT	42.299 70.164 42.331 70.228 ;
			RECT	42.467 70.164 42.499 70.228 ;
			RECT	42.635 70.164 42.667 70.228 ;
			RECT	42.803 70.164 42.835 70.228 ;
			RECT	42.971 70.164 43.003 70.228 ;
			RECT	43.139 70.164 43.171 70.228 ;
			RECT	43.307 70.164 43.339 70.228 ;
			RECT	43.475 70.164 43.507 70.228 ;
			RECT	43.643 70.164 43.675 70.228 ;
			RECT	43.811 70.164 43.843 70.228 ;
			RECT	43.979 70.164 44.011 70.228 ;
			RECT	44.147 70.164 44.179 70.228 ;
			RECT	44.315 70.164 44.347 70.228 ;
			RECT	44.483 70.164 44.515 70.228 ;
			RECT	44.651 70.164 44.683 70.228 ;
			RECT	44.819 70.164 44.851 70.228 ;
			RECT	44.987 70.164 45.019 70.228 ;
			RECT	45.155 70.164 45.187 70.228 ;
			RECT	45.323 70.164 45.355 70.228 ;
			RECT	45.491 70.164 45.523 70.228 ;
			RECT	45.659 70.164 45.691 70.228 ;
			RECT	45.827 70.164 45.859 70.228 ;
			RECT	45.995 70.164 46.027 70.228 ;
			RECT	46.163 70.164 46.195 70.228 ;
			RECT	46.331 70.164 46.363 70.228 ;
			RECT	46.499 70.164 46.531 70.228 ;
			RECT	46.667 70.164 46.699 70.228 ;
			RECT	46.835 70.164 46.867 70.228 ;
			RECT	47.003 70.164 47.035 70.228 ;
			RECT	47.171 70.164 47.203 70.228 ;
			RECT	47.339 70.164 47.371 70.228 ;
			RECT	47.507 70.164 47.539 70.228 ;
			RECT	47.675 70.164 47.707 70.228 ;
			RECT	47.843 70.164 47.875 70.228 ;
			RECT	48.011 70.164 48.043 70.228 ;
			RECT	48.179 70.164 48.211 70.228 ;
			RECT	48.347 70.164 48.379 70.228 ;
			RECT	48.515 70.164 48.547 70.228 ;
			RECT	48.683 70.164 48.715 70.228 ;
			RECT	48.851 70.164 48.883 70.228 ;
			RECT	49.019 70.164 49.051 70.228 ;
			RECT	49.187 70.164 49.219 70.228 ;
			RECT	49.318 70.18 49.35 70.212 ;
			RECT	49.439 70.18 49.471 70.212 ;
			RECT	49.569 70.164 49.601 70.228 ;
			RECT	51.881 70.164 51.913 70.228 ;
			RECT	53.132 70.164 53.196 70.228 ;
			RECT	53.812 70.164 53.844 70.228 ;
			RECT	54.251 70.164 54.283 70.228 ;
			RECT	55.562 70.164 55.626 70.228 ;
			RECT	58.603 70.164 58.635 70.228 ;
			RECT	58.733 70.18 58.765 70.212 ;
			RECT	58.854 70.18 58.886 70.212 ;
			RECT	58.985 70.164 59.017 70.228 ;
			RECT	59.153 70.164 59.185 70.228 ;
			RECT	59.321 70.164 59.353 70.228 ;
			RECT	59.489 70.164 59.521 70.228 ;
			RECT	59.657 70.164 59.689 70.228 ;
			RECT	59.825 70.164 59.857 70.228 ;
			RECT	59.993 70.164 60.025 70.228 ;
			RECT	60.161 70.164 60.193 70.228 ;
			RECT	60.329 70.164 60.361 70.228 ;
			RECT	60.497 70.164 60.529 70.228 ;
			RECT	60.665 70.164 60.697 70.228 ;
			RECT	60.833 70.164 60.865 70.228 ;
			RECT	61.001 70.164 61.033 70.228 ;
			RECT	61.169 70.164 61.201 70.228 ;
			RECT	61.337 70.164 61.369 70.228 ;
			RECT	61.505 70.164 61.537 70.228 ;
			RECT	61.673 70.164 61.705 70.228 ;
			RECT	61.841 70.164 61.873 70.228 ;
			RECT	62.009 70.164 62.041 70.228 ;
			RECT	62.177 70.164 62.209 70.228 ;
			RECT	62.345 70.164 62.377 70.228 ;
			RECT	62.513 70.164 62.545 70.228 ;
			RECT	62.681 70.164 62.713 70.228 ;
			RECT	62.849 70.164 62.881 70.228 ;
			RECT	63.017 70.164 63.049 70.228 ;
			RECT	63.185 70.164 63.217 70.228 ;
			RECT	63.353 70.164 63.385 70.228 ;
			RECT	63.521 70.164 63.553 70.228 ;
			RECT	63.689 70.164 63.721 70.228 ;
			RECT	63.857 70.164 63.889 70.228 ;
			RECT	64.025 70.164 64.057 70.228 ;
			RECT	64.193 70.164 64.225 70.228 ;
			RECT	64.361 70.164 64.393 70.228 ;
			RECT	64.529 70.164 64.561 70.228 ;
			RECT	64.697 70.164 64.729 70.228 ;
			RECT	64.865 70.164 64.897 70.228 ;
			RECT	65.033 70.164 65.065 70.228 ;
			RECT	65.201 70.164 65.233 70.228 ;
			RECT	65.369 70.164 65.401 70.228 ;
			RECT	65.537 70.164 65.569 70.228 ;
			RECT	65.705 70.164 65.737 70.228 ;
			RECT	65.873 70.164 65.905 70.228 ;
			RECT	66.041 70.164 66.073 70.228 ;
			RECT	66.209 70.164 66.241 70.228 ;
			RECT	66.377 70.164 66.409 70.228 ;
			RECT	66.545 70.164 66.577 70.228 ;
			RECT	66.713 70.164 66.745 70.228 ;
			RECT	66.881 70.164 66.913 70.228 ;
			RECT	67.049 70.164 67.081 70.228 ;
			RECT	67.217 70.164 67.249 70.228 ;
			RECT	67.385 70.164 67.417 70.228 ;
			RECT	67.553 70.164 67.585 70.228 ;
			RECT	67.721 70.164 67.753 70.228 ;
			RECT	67.889 70.164 67.921 70.228 ;
			RECT	68.057 70.164 68.089 70.228 ;
			RECT	68.225 70.164 68.257 70.228 ;
			RECT	68.393 70.164 68.425 70.228 ;
			RECT	68.561 70.164 68.593 70.228 ;
			RECT	68.729 70.164 68.761 70.228 ;
			RECT	68.897 70.164 68.929 70.228 ;
			RECT	69.065 70.164 69.097 70.228 ;
			RECT	69.233 70.164 69.265 70.228 ;
			RECT	69.401 70.164 69.433 70.228 ;
			RECT	69.569 70.164 69.601 70.228 ;
			RECT	69.737 70.164 69.769 70.228 ;
			RECT	69.905 70.164 69.937 70.228 ;
			RECT	70.073 70.164 70.105 70.228 ;
			RECT	70.241 70.164 70.273 70.228 ;
			RECT	70.409 70.164 70.441 70.228 ;
			RECT	70.577 70.164 70.609 70.228 ;
			RECT	70.745 70.164 70.777 70.228 ;
			RECT	70.913 70.164 70.945 70.228 ;
			RECT	71.081 70.164 71.113 70.228 ;
			RECT	71.249 70.164 71.281 70.228 ;
			RECT	71.417 70.164 71.449 70.228 ;
			RECT	71.585 70.164 71.617 70.228 ;
			RECT	71.753 70.164 71.785 70.228 ;
			RECT	71.921 70.164 71.953 70.228 ;
			RECT	72.089 70.164 72.121 70.228 ;
			RECT	72.257 70.164 72.289 70.228 ;
			RECT	72.425 70.164 72.457 70.228 ;
			RECT	72.593 70.164 72.625 70.228 ;
			RECT	72.761 70.164 72.793 70.228 ;
			RECT	72.929 70.164 72.961 70.228 ;
			RECT	73.097 70.164 73.129 70.228 ;
			RECT	73.265 70.164 73.297 70.228 ;
			RECT	73.433 70.164 73.465 70.228 ;
			RECT	73.601 70.164 73.633 70.228 ;
			RECT	73.769 70.164 73.801 70.228 ;
			RECT	73.937 70.164 73.969 70.228 ;
			RECT	74.105 70.164 74.137 70.228 ;
			RECT	74.273 70.164 74.305 70.228 ;
			RECT	74.441 70.164 74.473 70.228 ;
			RECT	74.609 70.164 74.641 70.228 ;
			RECT	74.777 70.164 74.809 70.228 ;
			RECT	74.945 70.164 74.977 70.228 ;
			RECT	75.113 70.164 75.145 70.228 ;
			RECT	75.281 70.164 75.313 70.228 ;
			RECT	75.449 70.164 75.481 70.228 ;
			RECT	75.617 70.164 75.649 70.228 ;
			RECT	75.785 70.164 75.817 70.228 ;
			RECT	75.953 70.164 75.985 70.228 ;
			RECT	76.121 70.164 76.153 70.228 ;
			RECT	76.289 70.164 76.321 70.228 ;
			RECT	76.457 70.164 76.489 70.228 ;
			RECT	76.625 70.164 76.657 70.228 ;
			RECT	76.793 70.164 76.825 70.228 ;
			RECT	76.961 70.164 76.993 70.228 ;
			RECT	77.129 70.164 77.161 70.228 ;
			RECT	77.297 70.164 77.329 70.228 ;
			RECT	77.465 70.164 77.497 70.228 ;
			RECT	77.633 70.164 77.665 70.228 ;
			RECT	77.801 70.164 77.833 70.228 ;
			RECT	77.969 70.164 78.001 70.228 ;
			RECT	78.137 70.164 78.169 70.228 ;
			RECT	78.305 70.164 78.337 70.228 ;
			RECT	78.473 70.164 78.505 70.228 ;
			RECT	78.641 70.164 78.673 70.228 ;
			RECT	78.809 70.164 78.841 70.228 ;
			RECT	78.977 70.164 79.009 70.228 ;
			RECT	79.145 70.164 79.177 70.228 ;
			RECT	79.313 70.164 79.345 70.228 ;
			RECT	79.481 70.164 79.513 70.228 ;
			RECT	79.649 70.164 79.681 70.228 ;
			RECT	79.817 70.164 79.849 70.228 ;
			RECT	79.985 70.164 80.017 70.228 ;
			RECT	80.153 70.164 80.185 70.228 ;
			RECT	80.321 70.164 80.353 70.228 ;
			RECT	80.489 70.164 80.521 70.228 ;
			RECT	80.657 70.164 80.689 70.228 ;
			RECT	80.825 70.164 80.857 70.228 ;
			RECT	80.993 70.164 81.025 70.228 ;
			RECT	81.161 70.164 81.193 70.228 ;
			RECT	81.329 70.164 81.361 70.228 ;
			RECT	81.497 70.164 81.529 70.228 ;
			RECT	81.665 70.164 81.697 70.228 ;
			RECT	81.833 70.164 81.865 70.228 ;
			RECT	82.001 70.164 82.033 70.228 ;
			RECT	82.169 70.164 82.201 70.228 ;
			RECT	82.337 70.164 82.369 70.228 ;
			RECT	82.505 70.164 82.537 70.228 ;
			RECT	82.673 70.164 82.705 70.228 ;
			RECT	82.841 70.164 82.873 70.228 ;
			RECT	83.009 70.164 83.041 70.228 ;
			RECT	83.177 70.164 83.209 70.228 ;
			RECT	83.345 70.164 83.377 70.228 ;
			RECT	83.513 70.164 83.545 70.228 ;
			RECT	83.681 70.164 83.713 70.228 ;
			RECT	83.849 70.164 83.881 70.228 ;
			RECT	84.017 70.164 84.049 70.228 ;
			RECT	84.185 70.164 84.217 70.228 ;
			RECT	84.353 70.164 84.385 70.228 ;
			RECT	84.521 70.164 84.553 70.228 ;
			RECT	84.689 70.164 84.721 70.228 ;
			RECT	84.857 70.164 84.889 70.228 ;
			RECT	85.025 70.164 85.057 70.228 ;
			RECT	85.193 70.164 85.225 70.228 ;
			RECT	85.361 70.164 85.393 70.228 ;
			RECT	85.529 70.164 85.561 70.228 ;
			RECT	85.697 70.164 85.729 70.228 ;
			RECT	85.865 70.164 85.897 70.228 ;
			RECT	86.033 70.164 86.065 70.228 ;
			RECT	86.201 70.164 86.233 70.228 ;
			RECT	86.369 70.164 86.401 70.228 ;
			RECT	86.537 70.164 86.569 70.228 ;
			RECT	86.705 70.164 86.737 70.228 ;
			RECT	86.873 70.164 86.905 70.228 ;
			RECT	87.041 70.164 87.073 70.228 ;
			RECT	87.209 70.164 87.241 70.228 ;
			RECT	87.377 70.164 87.409 70.228 ;
			RECT	87.545 70.164 87.577 70.228 ;
			RECT	87.713 70.164 87.745 70.228 ;
			RECT	87.881 70.164 87.913 70.228 ;
			RECT	88.049 70.164 88.081 70.228 ;
			RECT	88.217 70.164 88.249 70.228 ;
			RECT	88.385 70.164 88.417 70.228 ;
			RECT	88.553 70.164 88.585 70.228 ;
			RECT	88.721 70.164 88.753 70.228 ;
			RECT	88.889 70.164 88.921 70.228 ;
			RECT	89.057 70.164 89.089 70.228 ;
			RECT	89.225 70.164 89.257 70.228 ;
			RECT	89.393 70.164 89.425 70.228 ;
			RECT	89.561 70.164 89.593 70.228 ;
			RECT	89.729 70.164 89.761 70.228 ;
			RECT	89.897 70.164 89.929 70.228 ;
			RECT	90.065 70.164 90.097 70.228 ;
			RECT	90.233 70.164 90.265 70.228 ;
			RECT	90.401 70.164 90.433 70.228 ;
			RECT	90.569 70.164 90.601 70.228 ;
			RECT	90.737 70.164 90.769 70.228 ;
			RECT	90.905 70.164 90.937 70.228 ;
			RECT	91.073 70.164 91.105 70.228 ;
			RECT	91.241 70.164 91.273 70.228 ;
			RECT	91.409 70.164 91.441 70.228 ;
			RECT	91.577 70.164 91.609 70.228 ;
			RECT	91.745 70.164 91.777 70.228 ;
			RECT	91.913 70.164 91.945 70.228 ;
			RECT	92.081 70.164 92.113 70.228 ;
			RECT	92.249 70.164 92.281 70.228 ;
			RECT	92.417 70.164 92.449 70.228 ;
			RECT	92.585 70.164 92.617 70.228 ;
			RECT	92.753 70.164 92.785 70.228 ;
			RECT	92.921 70.164 92.953 70.228 ;
			RECT	93.089 70.164 93.121 70.228 ;
			RECT	93.257 70.164 93.289 70.228 ;
			RECT	93.425 70.164 93.457 70.228 ;
			RECT	93.593 70.164 93.625 70.228 ;
			RECT	93.761 70.164 93.793 70.228 ;
			RECT	93.929 70.164 93.961 70.228 ;
			RECT	94.097 70.164 94.129 70.228 ;
			RECT	94.265 70.164 94.297 70.228 ;
			RECT	94.433 70.164 94.465 70.228 ;
			RECT	94.601 70.164 94.633 70.228 ;
			RECT	94.769 70.164 94.801 70.228 ;
			RECT	94.937 70.164 94.969 70.228 ;
			RECT	95.105 70.164 95.137 70.228 ;
			RECT	95.273 70.164 95.305 70.228 ;
			RECT	95.441 70.164 95.473 70.228 ;
			RECT	95.609 70.164 95.641 70.228 ;
			RECT	95.777 70.164 95.809 70.228 ;
			RECT	95.945 70.164 95.977 70.228 ;
			RECT	96.113 70.164 96.145 70.228 ;
			RECT	96.281 70.164 96.313 70.228 ;
			RECT	96.449 70.164 96.481 70.228 ;
			RECT	96.617 70.164 96.649 70.228 ;
			RECT	96.785 70.164 96.817 70.228 ;
			RECT	96.953 70.164 96.985 70.228 ;
			RECT	97.121 70.164 97.153 70.228 ;
			RECT	97.289 70.164 97.321 70.228 ;
			RECT	97.457 70.164 97.489 70.228 ;
			RECT	97.625 70.164 97.657 70.228 ;
			RECT	97.793 70.164 97.825 70.228 ;
			RECT	97.961 70.164 97.993 70.228 ;
			RECT	98.129 70.164 98.161 70.228 ;
			RECT	98.297 70.164 98.329 70.228 ;
			RECT	98.465 70.164 98.497 70.228 ;
			RECT	98.633 70.164 98.665 70.228 ;
			RECT	98.801 70.164 98.833 70.228 ;
			RECT	98.969 70.164 99.001 70.228 ;
			RECT	99.137 70.164 99.169 70.228 ;
			RECT	99.305 70.164 99.337 70.228 ;
			RECT	99.473 70.164 99.505 70.228 ;
			RECT	99.641 70.164 99.673 70.228 ;
			RECT	99.809 70.164 99.841 70.228 ;
			RECT	99.977 70.164 100.009 70.228 ;
			RECT	100.145 70.164 100.177 70.228 ;
			RECT	100.313 70.164 100.345 70.228 ;
			RECT	100.481 70.164 100.513 70.228 ;
			RECT	100.649 70.164 100.681 70.228 ;
			RECT	100.817 70.164 100.849 70.228 ;
			RECT	100.985 70.164 101.017 70.228 ;
			RECT	101.153 70.164 101.185 70.228 ;
			RECT	101.321 70.164 101.353 70.228 ;
			RECT	101.489 70.164 101.521 70.228 ;
			RECT	101.657 70.164 101.689 70.228 ;
			RECT	101.825 70.164 101.857 70.228 ;
			RECT	101.993 70.164 102.025 70.228 ;
			RECT	102.123 70.18 102.155 70.212 ;
			RECT	102.245 70.175 102.277 70.207 ;
			RECT	102.375 70.164 102.407 70.228 ;
			RECT	103.795 70.164 103.827 70.228 ;
			RECT	103.925 70.175 103.957 70.207 ;
			RECT	104.047 70.18 104.079 70.212 ;
			RECT	104.177 70.164 104.209 70.228 ;
			RECT	104.345 70.164 104.377 70.228 ;
			RECT	104.513 70.164 104.545 70.228 ;
			RECT	104.681 70.164 104.713 70.228 ;
			RECT	104.849 70.164 104.881 70.228 ;
			RECT	105.017 70.164 105.049 70.228 ;
			RECT	105.185 70.164 105.217 70.228 ;
			RECT	105.353 70.164 105.385 70.228 ;
			RECT	105.521 70.164 105.553 70.228 ;
			RECT	105.689 70.164 105.721 70.228 ;
			RECT	105.857 70.164 105.889 70.228 ;
			RECT	106.025 70.164 106.057 70.228 ;
			RECT	106.193 70.164 106.225 70.228 ;
			RECT	106.361 70.164 106.393 70.228 ;
			RECT	106.529 70.164 106.561 70.228 ;
			RECT	106.697 70.164 106.729 70.228 ;
			RECT	106.865 70.164 106.897 70.228 ;
			RECT	107.033 70.164 107.065 70.228 ;
			RECT	107.201 70.164 107.233 70.228 ;
			RECT	107.369 70.164 107.401 70.228 ;
			RECT	107.537 70.164 107.569 70.228 ;
			RECT	107.705 70.164 107.737 70.228 ;
			RECT	107.873 70.164 107.905 70.228 ;
			RECT	108.041 70.164 108.073 70.228 ;
			RECT	108.209 70.164 108.241 70.228 ;
			RECT	108.377 70.164 108.409 70.228 ;
			RECT	108.545 70.164 108.577 70.228 ;
			RECT	108.713 70.164 108.745 70.228 ;
			RECT	108.881 70.164 108.913 70.228 ;
			RECT	109.049 70.164 109.081 70.228 ;
			RECT	109.217 70.164 109.249 70.228 ;
			RECT	109.385 70.164 109.417 70.228 ;
			RECT	109.553 70.164 109.585 70.228 ;
			RECT	109.721 70.164 109.753 70.228 ;
			RECT	109.889 70.164 109.921 70.228 ;
			RECT	110.057 70.164 110.089 70.228 ;
			RECT	110.225 70.164 110.257 70.228 ;
			RECT	110.393 70.164 110.425 70.228 ;
			RECT	110.561 70.164 110.593 70.228 ;
			RECT	110.729 70.164 110.761 70.228 ;
			RECT	110.897 70.164 110.929 70.228 ;
			RECT	111.065 70.164 111.097 70.228 ;
			RECT	111.233 70.164 111.265 70.228 ;
			RECT	111.401 70.164 111.433 70.228 ;
			RECT	111.569 70.164 111.601 70.228 ;
			RECT	111.737 70.164 111.769 70.228 ;
			RECT	111.905 70.164 111.937 70.228 ;
			RECT	112.073 70.164 112.105 70.228 ;
			RECT	112.241 70.164 112.273 70.228 ;
			RECT	112.409 70.164 112.441 70.228 ;
			RECT	112.577 70.164 112.609 70.228 ;
			RECT	112.745 70.164 112.777 70.228 ;
			RECT	112.913 70.164 112.945 70.228 ;
			RECT	113.081 70.164 113.113 70.228 ;
			RECT	113.249 70.164 113.281 70.228 ;
			RECT	113.417 70.164 113.449 70.228 ;
			RECT	113.585 70.164 113.617 70.228 ;
			RECT	113.753 70.164 113.785 70.228 ;
			RECT	113.921 70.164 113.953 70.228 ;
			RECT	114.089 70.164 114.121 70.228 ;
			RECT	114.257 70.164 114.289 70.228 ;
			RECT	114.425 70.164 114.457 70.228 ;
			RECT	114.593 70.164 114.625 70.228 ;
			RECT	114.761 70.164 114.793 70.228 ;
			RECT	114.929 70.164 114.961 70.228 ;
			RECT	115.097 70.164 115.129 70.228 ;
			RECT	115.265 70.164 115.297 70.228 ;
			RECT	115.433 70.164 115.465 70.228 ;
			RECT	115.601 70.164 115.633 70.228 ;
			RECT	115.769 70.164 115.801 70.228 ;
			RECT	115.937 70.164 115.969 70.228 ;
			RECT	116.105 70.164 116.137 70.228 ;
			RECT	116.273 70.164 116.305 70.228 ;
			RECT	116.441 70.164 116.473 70.228 ;
			RECT	116.609 70.164 116.641 70.228 ;
			RECT	116.777 70.164 116.809 70.228 ;
			RECT	116.945 70.164 116.977 70.228 ;
			RECT	117.113 70.164 117.145 70.228 ;
			RECT	117.281 70.164 117.313 70.228 ;
			RECT	117.449 70.164 117.481 70.228 ;
			RECT	117.617 70.164 117.649 70.228 ;
			RECT	117.785 70.164 117.817 70.228 ;
			RECT	117.953 70.164 117.985 70.228 ;
			RECT	118.121 70.164 118.153 70.228 ;
			RECT	118.289 70.164 118.321 70.228 ;
			RECT	118.457 70.164 118.489 70.228 ;
			RECT	118.625 70.164 118.657 70.228 ;
			RECT	118.793 70.164 118.825 70.228 ;
			RECT	118.961 70.164 118.993 70.228 ;
			RECT	119.129 70.164 119.161 70.228 ;
			RECT	119.297 70.164 119.329 70.228 ;
			RECT	119.465 70.164 119.497 70.228 ;
			RECT	119.633 70.164 119.665 70.228 ;
			RECT	119.801 70.164 119.833 70.228 ;
			RECT	119.969 70.164 120.001 70.228 ;
			RECT	120.137 70.164 120.169 70.228 ;
			RECT	120.305 70.164 120.337 70.228 ;
			RECT	120.473 70.164 120.505 70.228 ;
			RECT	120.641 70.164 120.673 70.228 ;
			RECT	120.809 70.164 120.841 70.228 ;
			RECT	120.977 70.164 121.009 70.228 ;
			RECT	121.145 70.164 121.177 70.228 ;
			RECT	121.313 70.164 121.345 70.228 ;
			RECT	121.481 70.164 121.513 70.228 ;
			RECT	121.649 70.164 121.681 70.228 ;
			RECT	121.817 70.164 121.849 70.228 ;
			RECT	121.985 70.164 122.017 70.228 ;
			RECT	122.153 70.164 122.185 70.228 ;
			RECT	122.321 70.164 122.353 70.228 ;
			RECT	122.489 70.164 122.521 70.228 ;
			RECT	122.657 70.164 122.689 70.228 ;
			RECT	122.825 70.164 122.857 70.228 ;
			RECT	122.993 70.164 123.025 70.228 ;
			RECT	123.161 70.164 123.193 70.228 ;
			RECT	123.329 70.164 123.361 70.228 ;
			RECT	123.497 70.164 123.529 70.228 ;
			RECT	123.665 70.164 123.697 70.228 ;
			RECT	123.833 70.164 123.865 70.228 ;
			RECT	124.001 70.164 124.033 70.228 ;
			RECT	124.169 70.164 124.201 70.228 ;
			RECT	124.337 70.164 124.369 70.228 ;
			RECT	124.505 70.164 124.537 70.228 ;
			RECT	124.673 70.164 124.705 70.228 ;
			RECT	124.841 70.164 124.873 70.228 ;
			RECT	125.009 70.164 125.041 70.228 ;
			RECT	125.177 70.164 125.209 70.228 ;
			RECT	125.345 70.164 125.377 70.228 ;
			RECT	125.513 70.164 125.545 70.228 ;
			RECT	125.681 70.164 125.713 70.228 ;
			RECT	125.849 70.164 125.881 70.228 ;
			RECT	126.017 70.164 126.049 70.228 ;
			RECT	126.185 70.164 126.217 70.228 ;
			RECT	126.353 70.164 126.385 70.228 ;
			RECT	126.521 70.164 126.553 70.228 ;
			RECT	126.689 70.164 126.721 70.228 ;
			RECT	126.857 70.164 126.889 70.228 ;
			RECT	127.025 70.164 127.057 70.228 ;
			RECT	127.193 70.164 127.225 70.228 ;
			RECT	127.361 70.164 127.393 70.228 ;
			RECT	127.529 70.164 127.561 70.228 ;
			RECT	127.697 70.164 127.729 70.228 ;
			RECT	127.865 70.164 127.897 70.228 ;
			RECT	128.033 70.164 128.065 70.228 ;
			RECT	128.201 70.164 128.233 70.228 ;
			RECT	128.369 70.164 128.401 70.228 ;
			RECT	128.537 70.164 128.569 70.228 ;
			RECT	128.705 70.164 128.737 70.228 ;
			RECT	128.873 70.164 128.905 70.228 ;
			RECT	129.041 70.164 129.073 70.228 ;
			RECT	129.209 70.164 129.241 70.228 ;
			RECT	129.377 70.164 129.409 70.228 ;
			RECT	129.545 70.164 129.577 70.228 ;
			RECT	129.713 70.164 129.745 70.228 ;
			RECT	129.881 70.164 129.913 70.228 ;
			RECT	130.049 70.164 130.081 70.228 ;
			RECT	130.217 70.164 130.249 70.228 ;
			RECT	130.385 70.164 130.417 70.228 ;
			RECT	130.553 70.164 130.585 70.228 ;
			RECT	130.721 70.164 130.753 70.228 ;
			RECT	130.889 70.164 130.921 70.228 ;
			RECT	131.057 70.164 131.089 70.228 ;
			RECT	131.225 70.164 131.257 70.228 ;
			RECT	131.393 70.164 131.425 70.228 ;
			RECT	131.561 70.164 131.593 70.228 ;
			RECT	131.729 70.164 131.761 70.228 ;
			RECT	131.897 70.164 131.929 70.228 ;
			RECT	132.065 70.164 132.097 70.228 ;
			RECT	132.233 70.164 132.265 70.228 ;
			RECT	132.401 70.164 132.433 70.228 ;
			RECT	132.569 70.164 132.601 70.228 ;
			RECT	132.737 70.164 132.769 70.228 ;
			RECT	132.905 70.164 132.937 70.228 ;
			RECT	133.073 70.164 133.105 70.228 ;
			RECT	133.241 70.164 133.273 70.228 ;
			RECT	133.409 70.164 133.441 70.228 ;
			RECT	133.577 70.164 133.609 70.228 ;
			RECT	133.745 70.164 133.777 70.228 ;
			RECT	133.913 70.164 133.945 70.228 ;
			RECT	134.081 70.164 134.113 70.228 ;
			RECT	134.249 70.164 134.281 70.228 ;
			RECT	134.417 70.164 134.449 70.228 ;
			RECT	134.585 70.164 134.617 70.228 ;
			RECT	134.753 70.164 134.785 70.228 ;
			RECT	134.921 70.164 134.953 70.228 ;
			RECT	135.089 70.164 135.121 70.228 ;
			RECT	135.257 70.164 135.289 70.228 ;
			RECT	135.425 70.164 135.457 70.228 ;
			RECT	135.593 70.164 135.625 70.228 ;
			RECT	135.761 70.164 135.793 70.228 ;
			RECT	135.929 70.164 135.961 70.228 ;
			RECT	136.097 70.164 136.129 70.228 ;
			RECT	136.265 70.164 136.297 70.228 ;
			RECT	136.433 70.164 136.465 70.228 ;
			RECT	136.601 70.164 136.633 70.228 ;
			RECT	136.769 70.164 136.801 70.228 ;
			RECT	136.937 70.164 136.969 70.228 ;
			RECT	137.105 70.164 137.137 70.228 ;
			RECT	137.273 70.164 137.305 70.228 ;
			RECT	137.441 70.164 137.473 70.228 ;
			RECT	137.609 70.164 137.641 70.228 ;
			RECT	137.777 70.164 137.809 70.228 ;
			RECT	137.945 70.164 137.977 70.228 ;
			RECT	138.113 70.164 138.145 70.228 ;
			RECT	138.281 70.164 138.313 70.228 ;
			RECT	138.449 70.164 138.481 70.228 ;
			RECT	138.617 70.164 138.649 70.228 ;
			RECT	138.785 70.164 138.817 70.228 ;
			RECT	138.953 70.164 138.985 70.228 ;
			RECT	139.121 70.164 139.153 70.228 ;
			RECT	139.289 70.164 139.321 70.228 ;
			RECT	139.457 70.164 139.489 70.228 ;
			RECT	139.625 70.164 139.657 70.228 ;
			RECT	139.793 70.164 139.825 70.228 ;
			RECT	139.961 70.164 139.993 70.228 ;
			RECT	140.129 70.164 140.161 70.228 ;
			RECT	140.297 70.164 140.329 70.228 ;
			RECT	140.465 70.164 140.497 70.228 ;
			RECT	140.633 70.164 140.665 70.228 ;
			RECT	140.801 70.164 140.833 70.228 ;
			RECT	140.969 70.164 141.001 70.228 ;
			RECT	141.137 70.164 141.169 70.228 ;
			RECT	141.305 70.164 141.337 70.228 ;
			RECT	141.473 70.164 141.505 70.228 ;
			RECT	141.641 70.164 141.673 70.228 ;
			RECT	141.809 70.164 141.841 70.228 ;
			RECT	141.977 70.164 142.009 70.228 ;
			RECT	142.145 70.164 142.177 70.228 ;
			RECT	142.313 70.164 142.345 70.228 ;
			RECT	142.481 70.164 142.513 70.228 ;
			RECT	142.649 70.164 142.681 70.228 ;
			RECT	142.817 70.164 142.849 70.228 ;
			RECT	142.985 70.164 143.017 70.228 ;
			RECT	143.153 70.164 143.185 70.228 ;
			RECT	143.321 70.164 143.353 70.228 ;
			RECT	143.489 70.164 143.521 70.228 ;
			RECT	143.657 70.164 143.689 70.228 ;
			RECT	143.825 70.164 143.857 70.228 ;
			RECT	143.993 70.164 144.025 70.228 ;
			RECT	144.161 70.164 144.193 70.228 ;
			RECT	144.329 70.164 144.361 70.228 ;
			RECT	144.497 70.164 144.529 70.228 ;
			RECT	144.665 70.164 144.697 70.228 ;
			RECT	144.833 70.164 144.865 70.228 ;
			RECT	145.001 70.164 145.033 70.228 ;
			RECT	145.169 70.164 145.201 70.228 ;
			RECT	145.337 70.164 145.369 70.228 ;
			RECT	145.505 70.164 145.537 70.228 ;
			RECT	145.673 70.164 145.705 70.228 ;
			RECT	145.841 70.164 145.873 70.228 ;
			RECT	146.009 70.164 146.041 70.228 ;
			RECT	146.177 70.164 146.209 70.228 ;
			RECT	146.345 70.164 146.377 70.228 ;
			RECT	146.513 70.164 146.545 70.228 ;
			RECT	146.681 70.164 146.713 70.228 ;
			RECT	146.849 70.164 146.881 70.228 ;
			RECT	147.017 70.164 147.049 70.228 ;
			RECT	147.185 70.164 147.217 70.228 ;
			RECT	147.316 70.18 147.348 70.212 ;
			RECT	147.437 70.18 147.469 70.212 ;
			RECT	147.567 70.164 147.599 70.228 ;
			RECT	149.879 70.164 149.911 70.228 ;
			RECT	151.13 70.164 151.194 70.228 ;
			RECT	151.81 70.164 151.842 70.228 ;
			RECT	152.249 70.164 152.281 70.228 ;
			RECT	153.56 70.164 153.624 70.228 ;
			RECT	156.601 70.164 156.633 70.228 ;
			RECT	156.731 70.18 156.763 70.212 ;
			RECT	156.852 70.18 156.884 70.212 ;
			RECT	156.983 70.164 157.015 70.228 ;
			RECT	157.151 70.164 157.183 70.228 ;
			RECT	157.319 70.164 157.351 70.228 ;
			RECT	157.487 70.164 157.519 70.228 ;
			RECT	157.655 70.164 157.687 70.228 ;
			RECT	157.823 70.164 157.855 70.228 ;
			RECT	157.991 70.164 158.023 70.228 ;
			RECT	158.159 70.164 158.191 70.228 ;
			RECT	158.327 70.164 158.359 70.228 ;
			RECT	158.495 70.164 158.527 70.228 ;
			RECT	158.663 70.164 158.695 70.228 ;
			RECT	158.831 70.164 158.863 70.228 ;
			RECT	158.999 70.164 159.031 70.228 ;
			RECT	159.167 70.164 159.199 70.228 ;
			RECT	159.335 70.164 159.367 70.228 ;
			RECT	159.503 70.164 159.535 70.228 ;
			RECT	159.671 70.164 159.703 70.228 ;
			RECT	159.839 70.164 159.871 70.228 ;
			RECT	160.007 70.164 160.039 70.228 ;
			RECT	160.175 70.164 160.207 70.228 ;
			RECT	160.343 70.164 160.375 70.228 ;
			RECT	160.511 70.164 160.543 70.228 ;
			RECT	160.679 70.164 160.711 70.228 ;
			RECT	160.847 70.164 160.879 70.228 ;
			RECT	161.015 70.164 161.047 70.228 ;
			RECT	161.183 70.164 161.215 70.228 ;
			RECT	161.351 70.164 161.383 70.228 ;
			RECT	161.519 70.164 161.551 70.228 ;
			RECT	161.687 70.164 161.719 70.228 ;
			RECT	161.855 70.164 161.887 70.228 ;
			RECT	162.023 70.164 162.055 70.228 ;
			RECT	162.191 70.164 162.223 70.228 ;
			RECT	162.359 70.164 162.391 70.228 ;
			RECT	162.527 70.164 162.559 70.228 ;
			RECT	162.695 70.164 162.727 70.228 ;
			RECT	162.863 70.164 162.895 70.228 ;
			RECT	163.031 70.164 163.063 70.228 ;
			RECT	163.199 70.164 163.231 70.228 ;
			RECT	163.367 70.164 163.399 70.228 ;
			RECT	163.535 70.164 163.567 70.228 ;
			RECT	163.703 70.164 163.735 70.228 ;
			RECT	163.871 70.164 163.903 70.228 ;
			RECT	164.039 70.164 164.071 70.228 ;
			RECT	164.207 70.164 164.239 70.228 ;
			RECT	164.375 70.164 164.407 70.228 ;
			RECT	164.543 70.164 164.575 70.228 ;
			RECT	164.711 70.164 164.743 70.228 ;
			RECT	164.879 70.164 164.911 70.228 ;
			RECT	165.047 70.164 165.079 70.228 ;
			RECT	165.215 70.164 165.247 70.228 ;
			RECT	165.383 70.164 165.415 70.228 ;
			RECT	165.551 70.164 165.583 70.228 ;
			RECT	165.719 70.164 165.751 70.228 ;
			RECT	165.887 70.164 165.919 70.228 ;
			RECT	166.055 70.164 166.087 70.228 ;
			RECT	166.223 70.164 166.255 70.228 ;
			RECT	166.391 70.164 166.423 70.228 ;
			RECT	166.559 70.164 166.591 70.228 ;
			RECT	166.727 70.164 166.759 70.228 ;
			RECT	166.895 70.164 166.927 70.228 ;
			RECT	167.063 70.164 167.095 70.228 ;
			RECT	167.231 70.164 167.263 70.228 ;
			RECT	167.399 70.164 167.431 70.228 ;
			RECT	167.567 70.164 167.599 70.228 ;
			RECT	167.735 70.164 167.767 70.228 ;
			RECT	167.903 70.164 167.935 70.228 ;
			RECT	168.071 70.164 168.103 70.228 ;
			RECT	168.239 70.164 168.271 70.228 ;
			RECT	168.407 70.164 168.439 70.228 ;
			RECT	168.575 70.164 168.607 70.228 ;
			RECT	168.743 70.164 168.775 70.228 ;
			RECT	168.911 70.164 168.943 70.228 ;
			RECT	169.079 70.164 169.111 70.228 ;
			RECT	169.247 70.164 169.279 70.228 ;
			RECT	169.415 70.164 169.447 70.228 ;
			RECT	169.583 70.164 169.615 70.228 ;
			RECT	169.751 70.164 169.783 70.228 ;
			RECT	169.919 70.164 169.951 70.228 ;
			RECT	170.087 70.164 170.119 70.228 ;
			RECT	170.255 70.164 170.287 70.228 ;
			RECT	170.423 70.164 170.455 70.228 ;
			RECT	170.591 70.164 170.623 70.228 ;
			RECT	170.759 70.164 170.791 70.228 ;
			RECT	170.927 70.164 170.959 70.228 ;
			RECT	171.095 70.164 171.127 70.228 ;
			RECT	171.263 70.164 171.295 70.228 ;
			RECT	171.431 70.164 171.463 70.228 ;
			RECT	171.599 70.164 171.631 70.228 ;
			RECT	171.767 70.164 171.799 70.228 ;
			RECT	171.935 70.164 171.967 70.228 ;
			RECT	172.103 70.164 172.135 70.228 ;
			RECT	172.271 70.164 172.303 70.228 ;
			RECT	172.439 70.164 172.471 70.228 ;
			RECT	172.607 70.164 172.639 70.228 ;
			RECT	172.775 70.164 172.807 70.228 ;
			RECT	172.943 70.164 172.975 70.228 ;
			RECT	173.111 70.164 173.143 70.228 ;
			RECT	173.279 70.164 173.311 70.228 ;
			RECT	173.447 70.164 173.479 70.228 ;
			RECT	173.615 70.164 173.647 70.228 ;
			RECT	173.783 70.164 173.815 70.228 ;
			RECT	173.951 70.164 173.983 70.228 ;
			RECT	174.119 70.164 174.151 70.228 ;
			RECT	174.287 70.164 174.319 70.228 ;
			RECT	174.455 70.164 174.487 70.228 ;
			RECT	174.623 70.164 174.655 70.228 ;
			RECT	174.791 70.164 174.823 70.228 ;
			RECT	174.959 70.164 174.991 70.228 ;
			RECT	175.127 70.164 175.159 70.228 ;
			RECT	175.295 70.164 175.327 70.228 ;
			RECT	175.463 70.164 175.495 70.228 ;
			RECT	175.631 70.164 175.663 70.228 ;
			RECT	175.799 70.164 175.831 70.228 ;
			RECT	175.967 70.164 175.999 70.228 ;
			RECT	176.135 70.164 176.167 70.228 ;
			RECT	176.303 70.164 176.335 70.228 ;
			RECT	176.471 70.164 176.503 70.228 ;
			RECT	176.639 70.164 176.671 70.228 ;
			RECT	176.807 70.164 176.839 70.228 ;
			RECT	176.975 70.164 177.007 70.228 ;
			RECT	177.143 70.164 177.175 70.228 ;
			RECT	177.311 70.164 177.343 70.228 ;
			RECT	177.479 70.164 177.511 70.228 ;
			RECT	177.647 70.164 177.679 70.228 ;
			RECT	177.815 70.164 177.847 70.228 ;
			RECT	177.983 70.164 178.015 70.228 ;
			RECT	178.151 70.164 178.183 70.228 ;
			RECT	178.319 70.164 178.351 70.228 ;
			RECT	178.487 70.164 178.519 70.228 ;
			RECT	178.655 70.164 178.687 70.228 ;
			RECT	178.823 70.164 178.855 70.228 ;
			RECT	178.991 70.164 179.023 70.228 ;
			RECT	179.159 70.164 179.191 70.228 ;
			RECT	179.327 70.164 179.359 70.228 ;
			RECT	179.495 70.164 179.527 70.228 ;
			RECT	179.663 70.164 179.695 70.228 ;
			RECT	179.831 70.164 179.863 70.228 ;
			RECT	179.999 70.164 180.031 70.228 ;
			RECT	180.167 70.164 180.199 70.228 ;
			RECT	180.335 70.164 180.367 70.228 ;
			RECT	180.503 70.164 180.535 70.228 ;
			RECT	180.671 70.164 180.703 70.228 ;
			RECT	180.839 70.164 180.871 70.228 ;
			RECT	181.007 70.164 181.039 70.228 ;
			RECT	181.175 70.164 181.207 70.228 ;
			RECT	181.343 70.164 181.375 70.228 ;
			RECT	181.511 70.164 181.543 70.228 ;
			RECT	181.679 70.164 181.711 70.228 ;
			RECT	181.847 70.164 181.879 70.228 ;
			RECT	182.015 70.164 182.047 70.228 ;
			RECT	182.183 70.164 182.215 70.228 ;
			RECT	182.351 70.164 182.383 70.228 ;
			RECT	182.519 70.164 182.551 70.228 ;
			RECT	182.687 70.164 182.719 70.228 ;
			RECT	182.855 70.164 182.887 70.228 ;
			RECT	183.023 70.164 183.055 70.228 ;
			RECT	183.191 70.164 183.223 70.228 ;
			RECT	183.359 70.164 183.391 70.228 ;
			RECT	183.527 70.164 183.559 70.228 ;
			RECT	183.695 70.164 183.727 70.228 ;
			RECT	183.863 70.164 183.895 70.228 ;
			RECT	184.031 70.164 184.063 70.228 ;
			RECT	184.199 70.164 184.231 70.228 ;
			RECT	184.367 70.164 184.399 70.228 ;
			RECT	184.535 70.164 184.567 70.228 ;
			RECT	184.703 70.164 184.735 70.228 ;
			RECT	184.871 70.164 184.903 70.228 ;
			RECT	185.039 70.164 185.071 70.228 ;
			RECT	185.207 70.164 185.239 70.228 ;
			RECT	185.375 70.164 185.407 70.228 ;
			RECT	185.543 70.164 185.575 70.228 ;
			RECT	185.711 70.164 185.743 70.228 ;
			RECT	185.879 70.164 185.911 70.228 ;
			RECT	186.047 70.164 186.079 70.228 ;
			RECT	186.215 70.164 186.247 70.228 ;
			RECT	186.383 70.164 186.415 70.228 ;
			RECT	186.551 70.164 186.583 70.228 ;
			RECT	186.719 70.164 186.751 70.228 ;
			RECT	186.887 70.164 186.919 70.228 ;
			RECT	187.055 70.164 187.087 70.228 ;
			RECT	187.223 70.164 187.255 70.228 ;
			RECT	187.391 70.164 187.423 70.228 ;
			RECT	187.559 70.164 187.591 70.228 ;
			RECT	187.727 70.164 187.759 70.228 ;
			RECT	187.895 70.164 187.927 70.228 ;
			RECT	188.063 70.164 188.095 70.228 ;
			RECT	188.231 70.164 188.263 70.228 ;
			RECT	188.399 70.164 188.431 70.228 ;
			RECT	188.567 70.164 188.599 70.228 ;
			RECT	188.735 70.164 188.767 70.228 ;
			RECT	188.903 70.164 188.935 70.228 ;
			RECT	189.071 70.164 189.103 70.228 ;
			RECT	189.239 70.164 189.271 70.228 ;
			RECT	189.407 70.164 189.439 70.228 ;
			RECT	189.575 70.164 189.607 70.228 ;
			RECT	189.743 70.164 189.775 70.228 ;
			RECT	189.911 70.164 189.943 70.228 ;
			RECT	190.079 70.164 190.111 70.228 ;
			RECT	190.247 70.164 190.279 70.228 ;
			RECT	190.415 70.164 190.447 70.228 ;
			RECT	190.583 70.164 190.615 70.228 ;
			RECT	190.751 70.164 190.783 70.228 ;
			RECT	190.919 70.164 190.951 70.228 ;
			RECT	191.087 70.164 191.119 70.228 ;
			RECT	191.255 70.164 191.287 70.228 ;
			RECT	191.423 70.164 191.455 70.228 ;
			RECT	191.591 70.164 191.623 70.228 ;
			RECT	191.759 70.164 191.791 70.228 ;
			RECT	191.927 70.164 191.959 70.228 ;
			RECT	192.095 70.164 192.127 70.228 ;
			RECT	192.263 70.164 192.295 70.228 ;
			RECT	192.431 70.164 192.463 70.228 ;
			RECT	192.599 70.164 192.631 70.228 ;
			RECT	192.767 70.164 192.799 70.228 ;
			RECT	192.935 70.164 192.967 70.228 ;
			RECT	193.103 70.164 193.135 70.228 ;
			RECT	193.271 70.164 193.303 70.228 ;
			RECT	193.439 70.164 193.471 70.228 ;
			RECT	193.607 70.164 193.639 70.228 ;
			RECT	193.775 70.164 193.807 70.228 ;
			RECT	193.943 70.164 193.975 70.228 ;
			RECT	194.111 70.164 194.143 70.228 ;
			RECT	194.279 70.164 194.311 70.228 ;
			RECT	194.447 70.164 194.479 70.228 ;
			RECT	194.615 70.164 194.647 70.228 ;
			RECT	194.783 70.164 194.815 70.228 ;
			RECT	194.951 70.164 194.983 70.228 ;
			RECT	195.119 70.164 195.151 70.228 ;
			RECT	195.287 70.164 195.319 70.228 ;
			RECT	195.455 70.164 195.487 70.228 ;
			RECT	195.623 70.164 195.655 70.228 ;
			RECT	195.791 70.164 195.823 70.228 ;
			RECT	195.959 70.164 195.991 70.228 ;
			RECT	196.127 70.164 196.159 70.228 ;
			RECT	196.295 70.164 196.327 70.228 ;
			RECT	196.463 70.164 196.495 70.228 ;
			RECT	196.631 70.164 196.663 70.228 ;
			RECT	196.799 70.164 196.831 70.228 ;
			RECT	196.967 70.164 196.999 70.228 ;
			RECT	197.135 70.164 197.167 70.228 ;
			RECT	197.303 70.164 197.335 70.228 ;
			RECT	197.471 70.164 197.503 70.228 ;
			RECT	197.639 70.164 197.671 70.228 ;
			RECT	197.807 70.164 197.839 70.228 ;
			RECT	197.975 70.164 198.007 70.228 ;
			RECT	198.143 70.164 198.175 70.228 ;
			RECT	198.311 70.164 198.343 70.228 ;
			RECT	198.479 70.164 198.511 70.228 ;
			RECT	198.647 70.164 198.679 70.228 ;
			RECT	198.815 70.164 198.847 70.228 ;
			RECT	198.983 70.164 199.015 70.228 ;
			RECT	199.151 70.164 199.183 70.228 ;
			RECT	199.319 70.164 199.351 70.228 ;
			RECT	199.487 70.164 199.519 70.228 ;
			RECT	199.655 70.164 199.687 70.228 ;
			RECT	199.823 70.164 199.855 70.228 ;
			RECT	199.991 70.164 200.023 70.228 ;
			RECT	200.121 70.18 200.153 70.212 ;
			RECT	200.243 70.175 200.275 70.207 ;
			RECT	200.373 70.164 200.405 70.228 ;
			RECT	200.9 70.164 200.932 70.228 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 68.216 201.665 68.336 ;
			LAYER	J3 ;
			RECT	0.755 68.244 0.787 68.308 ;
			RECT	1.645 68.244 1.709 68.308 ;
			RECT	2.323 68.244 2.387 68.308 ;
			RECT	3.438 68.244 3.47 68.308 ;
			RECT	3.585 68.244 3.617 68.308 ;
			RECT	4.195 68.244 4.227 68.308 ;
			RECT	4.72 68.244 4.752 68.308 ;
			RECT	4.944 68.244 5.008 68.308 ;
			RECT	5.267 68.244 5.299 68.308 ;
			RECT	5.797 68.244 5.829 68.308 ;
			RECT	5.927 68.255 5.959 68.287 ;
			RECT	6.049 68.26 6.081 68.292 ;
			RECT	6.179 68.244 6.211 68.308 ;
			RECT	6.347 68.244 6.379 68.308 ;
			RECT	6.515 68.244 6.547 68.308 ;
			RECT	6.683 68.244 6.715 68.308 ;
			RECT	6.851 68.244 6.883 68.308 ;
			RECT	7.019 68.244 7.051 68.308 ;
			RECT	7.187 68.244 7.219 68.308 ;
			RECT	7.355 68.244 7.387 68.308 ;
			RECT	7.523 68.244 7.555 68.308 ;
			RECT	7.691 68.244 7.723 68.308 ;
			RECT	7.859 68.244 7.891 68.308 ;
			RECT	8.027 68.244 8.059 68.308 ;
			RECT	8.195 68.244 8.227 68.308 ;
			RECT	8.363 68.244 8.395 68.308 ;
			RECT	8.531 68.244 8.563 68.308 ;
			RECT	8.699 68.244 8.731 68.308 ;
			RECT	8.867 68.244 8.899 68.308 ;
			RECT	9.035 68.244 9.067 68.308 ;
			RECT	9.203 68.244 9.235 68.308 ;
			RECT	9.371 68.244 9.403 68.308 ;
			RECT	9.539 68.244 9.571 68.308 ;
			RECT	9.707 68.244 9.739 68.308 ;
			RECT	9.875 68.244 9.907 68.308 ;
			RECT	10.043 68.244 10.075 68.308 ;
			RECT	10.211 68.244 10.243 68.308 ;
			RECT	10.379 68.244 10.411 68.308 ;
			RECT	10.547 68.244 10.579 68.308 ;
			RECT	10.715 68.244 10.747 68.308 ;
			RECT	10.883 68.244 10.915 68.308 ;
			RECT	11.051 68.244 11.083 68.308 ;
			RECT	11.219 68.244 11.251 68.308 ;
			RECT	11.387 68.244 11.419 68.308 ;
			RECT	11.555 68.244 11.587 68.308 ;
			RECT	11.723 68.244 11.755 68.308 ;
			RECT	11.891 68.244 11.923 68.308 ;
			RECT	12.059 68.244 12.091 68.308 ;
			RECT	12.227 68.244 12.259 68.308 ;
			RECT	12.395 68.244 12.427 68.308 ;
			RECT	12.563 68.244 12.595 68.308 ;
			RECT	12.731 68.244 12.763 68.308 ;
			RECT	12.899 68.244 12.931 68.308 ;
			RECT	13.067 68.244 13.099 68.308 ;
			RECT	13.235 68.244 13.267 68.308 ;
			RECT	13.403 68.244 13.435 68.308 ;
			RECT	13.571 68.244 13.603 68.308 ;
			RECT	13.739 68.244 13.771 68.308 ;
			RECT	13.907 68.244 13.939 68.308 ;
			RECT	14.075 68.244 14.107 68.308 ;
			RECT	14.243 68.244 14.275 68.308 ;
			RECT	14.411 68.244 14.443 68.308 ;
			RECT	14.579 68.244 14.611 68.308 ;
			RECT	14.747 68.244 14.779 68.308 ;
			RECT	14.915 68.244 14.947 68.308 ;
			RECT	15.083 68.244 15.115 68.308 ;
			RECT	15.251 68.244 15.283 68.308 ;
			RECT	15.419 68.244 15.451 68.308 ;
			RECT	15.587 68.244 15.619 68.308 ;
			RECT	15.755 68.244 15.787 68.308 ;
			RECT	15.923 68.244 15.955 68.308 ;
			RECT	16.091 68.244 16.123 68.308 ;
			RECT	16.259 68.244 16.291 68.308 ;
			RECT	16.427 68.244 16.459 68.308 ;
			RECT	16.595 68.244 16.627 68.308 ;
			RECT	16.763 68.244 16.795 68.308 ;
			RECT	16.931 68.244 16.963 68.308 ;
			RECT	17.099 68.244 17.131 68.308 ;
			RECT	17.267 68.244 17.299 68.308 ;
			RECT	17.435 68.244 17.467 68.308 ;
			RECT	17.603 68.244 17.635 68.308 ;
			RECT	17.771 68.244 17.803 68.308 ;
			RECT	17.939 68.244 17.971 68.308 ;
			RECT	18.107 68.244 18.139 68.308 ;
			RECT	18.275 68.244 18.307 68.308 ;
			RECT	18.443 68.244 18.475 68.308 ;
			RECT	18.611 68.244 18.643 68.308 ;
			RECT	18.779 68.244 18.811 68.308 ;
			RECT	18.947 68.244 18.979 68.308 ;
			RECT	19.115 68.244 19.147 68.308 ;
			RECT	19.283 68.244 19.315 68.308 ;
			RECT	19.451 68.244 19.483 68.308 ;
			RECT	19.619 68.244 19.651 68.308 ;
			RECT	19.787 68.244 19.819 68.308 ;
			RECT	19.955 68.244 19.987 68.308 ;
			RECT	20.123 68.244 20.155 68.308 ;
			RECT	20.291 68.244 20.323 68.308 ;
			RECT	20.459 68.244 20.491 68.308 ;
			RECT	20.627 68.244 20.659 68.308 ;
			RECT	20.795 68.244 20.827 68.308 ;
			RECT	20.963 68.244 20.995 68.308 ;
			RECT	21.131 68.244 21.163 68.308 ;
			RECT	21.299 68.244 21.331 68.308 ;
			RECT	21.467 68.244 21.499 68.308 ;
			RECT	21.635 68.244 21.667 68.308 ;
			RECT	21.803 68.244 21.835 68.308 ;
			RECT	21.971 68.244 22.003 68.308 ;
			RECT	22.139 68.244 22.171 68.308 ;
			RECT	22.307 68.244 22.339 68.308 ;
			RECT	22.475 68.244 22.507 68.308 ;
			RECT	22.643 68.244 22.675 68.308 ;
			RECT	22.811 68.244 22.843 68.308 ;
			RECT	22.979 68.244 23.011 68.308 ;
			RECT	23.147 68.244 23.179 68.308 ;
			RECT	23.315 68.244 23.347 68.308 ;
			RECT	23.483 68.244 23.515 68.308 ;
			RECT	23.651 68.244 23.683 68.308 ;
			RECT	23.819 68.244 23.851 68.308 ;
			RECT	23.987 68.244 24.019 68.308 ;
			RECT	24.155 68.244 24.187 68.308 ;
			RECT	24.323 68.244 24.355 68.308 ;
			RECT	24.491 68.244 24.523 68.308 ;
			RECT	24.659 68.244 24.691 68.308 ;
			RECT	24.827 68.244 24.859 68.308 ;
			RECT	24.995 68.244 25.027 68.308 ;
			RECT	25.163 68.244 25.195 68.308 ;
			RECT	25.331 68.244 25.363 68.308 ;
			RECT	25.499 68.244 25.531 68.308 ;
			RECT	25.667 68.244 25.699 68.308 ;
			RECT	25.835 68.244 25.867 68.308 ;
			RECT	26.003 68.244 26.035 68.308 ;
			RECT	26.171 68.244 26.203 68.308 ;
			RECT	26.339 68.244 26.371 68.308 ;
			RECT	26.507 68.244 26.539 68.308 ;
			RECT	26.675 68.244 26.707 68.308 ;
			RECT	26.843 68.244 26.875 68.308 ;
			RECT	27.011 68.244 27.043 68.308 ;
			RECT	27.179 68.244 27.211 68.308 ;
			RECT	27.347 68.244 27.379 68.308 ;
			RECT	27.515 68.244 27.547 68.308 ;
			RECT	27.683 68.244 27.715 68.308 ;
			RECT	27.851 68.244 27.883 68.308 ;
			RECT	28.019 68.244 28.051 68.308 ;
			RECT	28.187 68.244 28.219 68.308 ;
			RECT	28.355 68.244 28.387 68.308 ;
			RECT	28.523 68.244 28.555 68.308 ;
			RECT	28.691 68.244 28.723 68.308 ;
			RECT	28.859 68.244 28.891 68.308 ;
			RECT	29.027 68.244 29.059 68.308 ;
			RECT	29.195 68.244 29.227 68.308 ;
			RECT	29.363 68.244 29.395 68.308 ;
			RECT	29.531 68.244 29.563 68.308 ;
			RECT	29.699 68.244 29.731 68.308 ;
			RECT	29.867 68.244 29.899 68.308 ;
			RECT	30.035 68.244 30.067 68.308 ;
			RECT	30.203 68.244 30.235 68.308 ;
			RECT	30.371 68.244 30.403 68.308 ;
			RECT	30.539 68.244 30.571 68.308 ;
			RECT	30.707 68.244 30.739 68.308 ;
			RECT	30.875 68.244 30.907 68.308 ;
			RECT	31.043 68.244 31.075 68.308 ;
			RECT	31.211 68.244 31.243 68.308 ;
			RECT	31.379 68.244 31.411 68.308 ;
			RECT	31.547 68.244 31.579 68.308 ;
			RECT	31.715 68.244 31.747 68.308 ;
			RECT	31.883 68.244 31.915 68.308 ;
			RECT	32.051 68.244 32.083 68.308 ;
			RECT	32.219 68.244 32.251 68.308 ;
			RECT	32.387 68.244 32.419 68.308 ;
			RECT	32.555 68.244 32.587 68.308 ;
			RECT	32.723 68.244 32.755 68.308 ;
			RECT	32.891 68.244 32.923 68.308 ;
			RECT	33.059 68.244 33.091 68.308 ;
			RECT	33.227 68.244 33.259 68.308 ;
			RECT	33.395 68.244 33.427 68.308 ;
			RECT	33.563 68.244 33.595 68.308 ;
			RECT	33.731 68.244 33.763 68.308 ;
			RECT	33.899 68.244 33.931 68.308 ;
			RECT	34.067 68.244 34.099 68.308 ;
			RECT	34.235 68.244 34.267 68.308 ;
			RECT	34.403 68.244 34.435 68.308 ;
			RECT	34.571 68.244 34.603 68.308 ;
			RECT	34.739 68.244 34.771 68.308 ;
			RECT	34.907 68.244 34.939 68.308 ;
			RECT	35.075 68.244 35.107 68.308 ;
			RECT	35.243 68.244 35.275 68.308 ;
			RECT	35.411 68.244 35.443 68.308 ;
			RECT	35.579 68.244 35.611 68.308 ;
			RECT	35.747 68.244 35.779 68.308 ;
			RECT	35.915 68.244 35.947 68.308 ;
			RECT	36.083 68.244 36.115 68.308 ;
			RECT	36.251 68.244 36.283 68.308 ;
			RECT	36.419 68.244 36.451 68.308 ;
			RECT	36.587 68.244 36.619 68.308 ;
			RECT	36.755 68.244 36.787 68.308 ;
			RECT	36.923 68.244 36.955 68.308 ;
			RECT	37.091 68.244 37.123 68.308 ;
			RECT	37.259 68.244 37.291 68.308 ;
			RECT	37.427 68.244 37.459 68.308 ;
			RECT	37.595 68.244 37.627 68.308 ;
			RECT	37.763 68.244 37.795 68.308 ;
			RECT	37.931 68.244 37.963 68.308 ;
			RECT	38.099 68.244 38.131 68.308 ;
			RECT	38.267 68.244 38.299 68.308 ;
			RECT	38.435 68.244 38.467 68.308 ;
			RECT	38.603 68.244 38.635 68.308 ;
			RECT	38.771 68.244 38.803 68.308 ;
			RECT	38.939 68.244 38.971 68.308 ;
			RECT	39.107 68.244 39.139 68.308 ;
			RECT	39.275 68.244 39.307 68.308 ;
			RECT	39.443 68.244 39.475 68.308 ;
			RECT	39.611 68.244 39.643 68.308 ;
			RECT	39.779 68.244 39.811 68.308 ;
			RECT	39.947 68.244 39.979 68.308 ;
			RECT	40.115 68.244 40.147 68.308 ;
			RECT	40.283 68.244 40.315 68.308 ;
			RECT	40.451 68.244 40.483 68.308 ;
			RECT	40.619 68.244 40.651 68.308 ;
			RECT	40.787 68.244 40.819 68.308 ;
			RECT	40.955 68.244 40.987 68.308 ;
			RECT	41.123 68.244 41.155 68.308 ;
			RECT	41.291 68.244 41.323 68.308 ;
			RECT	41.459 68.244 41.491 68.308 ;
			RECT	41.627 68.244 41.659 68.308 ;
			RECT	41.795 68.244 41.827 68.308 ;
			RECT	41.963 68.244 41.995 68.308 ;
			RECT	42.131 68.244 42.163 68.308 ;
			RECT	42.299 68.244 42.331 68.308 ;
			RECT	42.467 68.244 42.499 68.308 ;
			RECT	42.635 68.244 42.667 68.308 ;
			RECT	42.803 68.244 42.835 68.308 ;
			RECT	42.971 68.244 43.003 68.308 ;
			RECT	43.139 68.244 43.171 68.308 ;
			RECT	43.307 68.244 43.339 68.308 ;
			RECT	43.475 68.244 43.507 68.308 ;
			RECT	43.643 68.244 43.675 68.308 ;
			RECT	43.811 68.244 43.843 68.308 ;
			RECT	43.979 68.244 44.011 68.308 ;
			RECT	44.147 68.244 44.179 68.308 ;
			RECT	44.315 68.244 44.347 68.308 ;
			RECT	44.483 68.244 44.515 68.308 ;
			RECT	44.651 68.244 44.683 68.308 ;
			RECT	44.819 68.244 44.851 68.308 ;
			RECT	44.987 68.244 45.019 68.308 ;
			RECT	45.155 68.244 45.187 68.308 ;
			RECT	45.323 68.244 45.355 68.308 ;
			RECT	45.491 68.244 45.523 68.308 ;
			RECT	45.659 68.244 45.691 68.308 ;
			RECT	45.827 68.244 45.859 68.308 ;
			RECT	45.995 68.244 46.027 68.308 ;
			RECT	46.163 68.244 46.195 68.308 ;
			RECT	46.331 68.244 46.363 68.308 ;
			RECT	46.499 68.244 46.531 68.308 ;
			RECT	46.667 68.244 46.699 68.308 ;
			RECT	46.835 68.244 46.867 68.308 ;
			RECT	47.003 68.244 47.035 68.308 ;
			RECT	47.171 68.244 47.203 68.308 ;
			RECT	47.339 68.244 47.371 68.308 ;
			RECT	47.507 68.244 47.539 68.308 ;
			RECT	47.675 68.244 47.707 68.308 ;
			RECT	47.843 68.244 47.875 68.308 ;
			RECT	48.011 68.244 48.043 68.308 ;
			RECT	48.179 68.244 48.211 68.308 ;
			RECT	48.347 68.244 48.379 68.308 ;
			RECT	48.515 68.244 48.547 68.308 ;
			RECT	48.683 68.244 48.715 68.308 ;
			RECT	48.851 68.244 48.883 68.308 ;
			RECT	49.019 68.244 49.051 68.308 ;
			RECT	49.187 68.244 49.219 68.308 ;
			RECT	49.318 68.26 49.35 68.292 ;
			RECT	49.439 68.26 49.471 68.292 ;
			RECT	49.569 68.244 49.601 68.308 ;
			RECT	51.881 68.244 51.913 68.308 ;
			RECT	53.132 68.244 53.196 68.308 ;
			RECT	53.812 68.244 53.844 68.308 ;
			RECT	54.251 68.244 54.283 68.308 ;
			RECT	55.562 68.244 55.626 68.308 ;
			RECT	58.603 68.244 58.635 68.308 ;
			RECT	58.733 68.26 58.765 68.292 ;
			RECT	58.854 68.26 58.886 68.292 ;
			RECT	58.985 68.244 59.017 68.308 ;
			RECT	59.153 68.244 59.185 68.308 ;
			RECT	59.321 68.244 59.353 68.308 ;
			RECT	59.489 68.244 59.521 68.308 ;
			RECT	59.657 68.244 59.689 68.308 ;
			RECT	59.825 68.244 59.857 68.308 ;
			RECT	59.993 68.244 60.025 68.308 ;
			RECT	60.161 68.244 60.193 68.308 ;
			RECT	60.329 68.244 60.361 68.308 ;
			RECT	60.497 68.244 60.529 68.308 ;
			RECT	60.665 68.244 60.697 68.308 ;
			RECT	60.833 68.244 60.865 68.308 ;
			RECT	61.001 68.244 61.033 68.308 ;
			RECT	61.169 68.244 61.201 68.308 ;
			RECT	61.337 68.244 61.369 68.308 ;
			RECT	61.505 68.244 61.537 68.308 ;
			RECT	61.673 68.244 61.705 68.308 ;
			RECT	61.841 68.244 61.873 68.308 ;
			RECT	62.009 68.244 62.041 68.308 ;
			RECT	62.177 68.244 62.209 68.308 ;
			RECT	62.345 68.244 62.377 68.308 ;
			RECT	62.513 68.244 62.545 68.308 ;
			RECT	62.681 68.244 62.713 68.308 ;
			RECT	62.849 68.244 62.881 68.308 ;
			RECT	63.017 68.244 63.049 68.308 ;
			RECT	63.185 68.244 63.217 68.308 ;
			RECT	63.353 68.244 63.385 68.308 ;
			RECT	63.521 68.244 63.553 68.308 ;
			RECT	63.689 68.244 63.721 68.308 ;
			RECT	63.857 68.244 63.889 68.308 ;
			RECT	64.025 68.244 64.057 68.308 ;
			RECT	64.193 68.244 64.225 68.308 ;
			RECT	64.361 68.244 64.393 68.308 ;
			RECT	64.529 68.244 64.561 68.308 ;
			RECT	64.697 68.244 64.729 68.308 ;
			RECT	64.865 68.244 64.897 68.308 ;
			RECT	65.033 68.244 65.065 68.308 ;
			RECT	65.201 68.244 65.233 68.308 ;
			RECT	65.369 68.244 65.401 68.308 ;
			RECT	65.537 68.244 65.569 68.308 ;
			RECT	65.705 68.244 65.737 68.308 ;
			RECT	65.873 68.244 65.905 68.308 ;
			RECT	66.041 68.244 66.073 68.308 ;
			RECT	66.209 68.244 66.241 68.308 ;
			RECT	66.377 68.244 66.409 68.308 ;
			RECT	66.545 68.244 66.577 68.308 ;
			RECT	66.713 68.244 66.745 68.308 ;
			RECT	66.881 68.244 66.913 68.308 ;
			RECT	67.049 68.244 67.081 68.308 ;
			RECT	67.217 68.244 67.249 68.308 ;
			RECT	67.385 68.244 67.417 68.308 ;
			RECT	67.553 68.244 67.585 68.308 ;
			RECT	67.721 68.244 67.753 68.308 ;
			RECT	67.889 68.244 67.921 68.308 ;
			RECT	68.057 68.244 68.089 68.308 ;
			RECT	68.225 68.244 68.257 68.308 ;
			RECT	68.393 68.244 68.425 68.308 ;
			RECT	68.561 68.244 68.593 68.308 ;
			RECT	68.729 68.244 68.761 68.308 ;
			RECT	68.897 68.244 68.929 68.308 ;
			RECT	69.065 68.244 69.097 68.308 ;
			RECT	69.233 68.244 69.265 68.308 ;
			RECT	69.401 68.244 69.433 68.308 ;
			RECT	69.569 68.244 69.601 68.308 ;
			RECT	69.737 68.244 69.769 68.308 ;
			RECT	69.905 68.244 69.937 68.308 ;
			RECT	70.073 68.244 70.105 68.308 ;
			RECT	70.241 68.244 70.273 68.308 ;
			RECT	70.409 68.244 70.441 68.308 ;
			RECT	70.577 68.244 70.609 68.308 ;
			RECT	70.745 68.244 70.777 68.308 ;
			RECT	70.913 68.244 70.945 68.308 ;
			RECT	71.081 68.244 71.113 68.308 ;
			RECT	71.249 68.244 71.281 68.308 ;
			RECT	71.417 68.244 71.449 68.308 ;
			RECT	71.585 68.244 71.617 68.308 ;
			RECT	71.753 68.244 71.785 68.308 ;
			RECT	71.921 68.244 71.953 68.308 ;
			RECT	72.089 68.244 72.121 68.308 ;
			RECT	72.257 68.244 72.289 68.308 ;
			RECT	72.425 68.244 72.457 68.308 ;
			RECT	72.593 68.244 72.625 68.308 ;
			RECT	72.761 68.244 72.793 68.308 ;
			RECT	72.929 68.244 72.961 68.308 ;
			RECT	73.097 68.244 73.129 68.308 ;
			RECT	73.265 68.244 73.297 68.308 ;
			RECT	73.433 68.244 73.465 68.308 ;
			RECT	73.601 68.244 73.633 68.308 ;
			RECT	73.769 68.244 73.801 68.308 ;
			RECT	73.937 68.244 73.969 68.308 ;
			RECT	74.105 68.244 74.137 68.308 ;
			RECT	74.273 68.244 74.305 68.308 ;
			RECT	74.441 68.244 74.473 68.308 ;
			RECT	74.609 68.244 74.641 68.308 ;
			RECT	74.777 68.244 74.809 68.308 ;
			RECT	74.945 68.244 74.977 68.308 ;
			RECT	75.113 68.244 75.145 68.308 ;
			RECT	75.281 68.244 75.313 68.308 ;
			RECT	75.449 68.244 75.481 68.308 ;
			RECT	75.617 68.244 75.649 68.308 ;
			RECT	75.785 68.244 75.817 68.308 ;
			RECT	75.953 68.244 75.985 68.308 ;
			RECT	76.121 68.244 76.153 68.308 ;
			RECT	76.289 68.244 76.321 68.308 ;
			RECT	76.457 68.244 76.489 68.308 ;
			RECT	76.625 68.244 76.657 68.308 ;
			RECT	76.793 68.244 76.825 68.308 ;
			RECT	76.961 68.244 76.993 68.308 ;
			RECT	77.129 68.244 77.161 68.308 ;
			RECT	77.297 68.244 77.329 68.308 ;
			RECT	77.465 68.244 77.497 68.308 ;
			RECT	77.633 68.244 77.665 68.308 ;
			RECT	77.801 68.244 77.833 68.308 ;
			RECT	77.969 68.244 78.001 68.308 ;
			RECT	78.137 68.244 78.169 68.308 ;
			RECT	78.305 68.244 78.337 68.308 ;
			RECT	78.473 68.244 78.505 68.308 ;
			RECT	78.641 68.244 78.673 68.308 ;
			RECT	78.809 68.244 78.841 68.308 ;
			RECT	78.977 68.244 79.009 68.308 ;
			RECT	79.145 68.244 79.177 68.308 ;
			RECT	79.313 68.244 79.345 68.308 ;
			RECT	79.481 68.244 79.513 68.308 ;
			RECT	79.649 68.244 79.681 68.308 ;
			RECT	79.817 68.244 79.849 68.308 ;
			RECT	79.985 68.244 80.017 68.308 ;
			RECT	80.153 68.244 80.185 68.308 ;
			RECT	80.321 68.244 80.353 68.308 ;
			RECT	80.489 68.244 80.521 68.308 ;
			RECT	80.657 68.244 80.689 68.308 ;
			RECT	80.825 68.244 80.857 68.308 ;
			RECT	80.993 68.244 81.025 68.308 ;
			RECT	81.161 68.244 81.193 68.308 ;
			RECT	81.329 68.244 81.361 68.308 ;
			RECT	81.497 68.244 81.529 68.308 ;
			RECT	81.665 68.244 81.697 68.308 ;
			RECT	81.833 68.244 81.865 68.308 ;
			RECT	82.001 68.244 82.033 68.308 ;
			RECT	82.169 68.244 82.201 68.308 ;
			RECT	82.337 68.244 82.369 68.308 ;
			RECT	82.505 68.244 82.537 68.308 ;
			RECT	82.673 68.244 82.705 68.308 ;
			RECT	82.841 68.244 82.873 68.308 ;
			RECT	83.009 68.244 83.041 68.308 ;
			RECT	83.177 68.244 83.209 68.308 ;
			RECT	83.345 68.244 83.377 68.308 ;
			RECT	83.513 68.244 83.545 68.308 ;
			RECT	83.681 68.244 83.713 68.308 ;
			RECT	83.849 68.244 83.881 68.308 ;
			RECT	84.017 68.244 84.049 68.308 ;
			RECT	84.185 68.244 84.217 68.308 ;
			RECT	84.353 68.244 84.385 68.308 ;
			RECT	84.521 68.244 84.553 68.308 ;
			RECT	84.689 68.244 84.721 68.308 ;
			RECT	84.857 68.244 84.889 68.308 ;
			RECT	85.025 68.244 85.057 68.308 ;
			RECT	85.193 68.244 85.225 68.308 ;
			RECT	85.361 68.244 85.393 68.308 ;
			RECT	85.529 68.244 85.561 68.308 ;
			RECT	85.697 68.244 85.729 68.308 ;
			RECT	85.865 68.244 85.897 68.308 ;
			RECT	86.033 68.244 86.065 68.308 ;
			RECT	86.201 68.244 86.233 68.308 ;
			RECT	86.369 68.244 86.401 68.308 ;
			RECT	86.537 68.244 86.569 68.308 ;
			RECT	86.705 68.244 86.737 68.308 ;
			RECT	86.873 68.244 86.905 68.308 ;
			RECT	87.041 68.244 87.073 68.308 ;
			RECT	87.209 68.244 87.241 68.308 ;
			RECT	87.377 68.244 87.409 68.308 ;
			RECT	87.545 68.244 87.577 68.308 ;
			RECT	87.713 68.244 87.745 68.308 ;
			RECT	87.881 68.244 87.913 68.308 ;
			RECT	88.049 68.244 88.081 68.308 ;
			RECT	88.217 68.244 88.249 68.308 ;
			RECT	88.385 68.244 88.417 68.308 ;
			RECT	88.553 68.244 88.585 68.308 ;
			RECT	88.721 68.244 88.753 68.308 ;
			RECT	88.889 68.244 88.921 68.308 ;
			RECT	89.057 68.244 89.089 68.308 ;
			RECT	89.225 68.244 89.257 68.308 ;
			RECT	89.393 68.244 89.425 68.308 ;
			RECT	89.561 68.244 89.593 68.308 ;
			RECT	89.729 68.244 89.761 68.308 ;
			RECT	89.897 68.244 89.929 68.308 ;
			RECT	90.065 68.244 90.097 68.308 ;
			RECT	90.233 68.244 90.265 68.308 ;
			RECT	90.401 68.244 90.433 68.308 ;
			RECT	90.569 68.244 90.601 68.308 ;
			RECT	90.737 68.244 90.769 68.308 ;
			RECT	90.905 68.244 90.937 68.308 ;
			RECT	91.073 68.244 91.105 68.308 ;
			RECT	91.241 68.244 91.273 68.308 ;
			RECT	91.409 68.244 91.441 68.308 ;
			RECT	91.577 68.244 91.609 68.308 ;
			RECT	91.745 68.244 91.777 68.308 ;
			RECT	91.913 68.244 91.945 68.308 ;
			RECT	92.081 68.244 92.113 68.308 ;
			RECT	92.249 68.244 92.281 68.308 ;
			RECT	92.417 68.244 92.449 68.308 ;
			RECT	92.585 68.244 92.617 68.308 ;
			RECT	92.753 68.244 92.785 68.308 ;
			RECT	92.921 68.244 92.953 68.308 ;
			RECT	93.089 68.244 93.121 68.308 ;
			RECT	93.257 68.244 93.289 68.308 ;
			RECT	93.425 68.244 93.457 68.308 ;
			RECT	93.593 68.244 93.625 68.308 ;
			RECT	93.761 68.244 93.793 68.308 ;
			RECT	93.929 68.244 93.961 68.308 ;
			RECT	94.097 68.244 94.129 68.308 ;
			RECT	94.265 68.244 94.297 68.308 ;
			RECT	94.433 68.244 94.465 68.308 ;
			RECT	94.601 68.244 94.633 68.308 ;
			RECT	94.769 68.244 94.801 68.308 ;
			RECT	94.937 68.244 94.969 68.308 ;
			RECT	95.105 68.244 95.137 68.308 ;
			RECT	95.273 68.244 95.305 68.308 ;
			RECT	95.441 68.244 95.473 68.308 ;
			RECT	95.609 68.244 95.641 68.308 ;
			RECT	95.777 68.244 95.809 68.308 ;
			RECT	95.945 68.244 95.977 68.308 ;
			RECT	96.113 68.244 96.145 68.308 ;
			RECT	96.281 68.244 96.313 68.308 ;
			RECT	96.449 68.244 96.481 68.308 ;
			RECT	96.617 68.244 96.649 68.308 ;
			RECT	96.785 68.244 96.817 68.308 ;
			RECT	96.953 68.244 96.985 68.308 ;
			RECT	97.121 68.244 97.153 68.308 ;
			RECT	97.289 68.244 97.321 68.308 ;
			RECT	97.457 68.244 97.489 68.308 ;
			RECT	97.625 68.244 97.657 68.308 ;
			RECT	97.793 68.244 97.825 68.308 ;
			RECT	97.961 68.244 97.993 68.308 ;
			RECT	98.129 68.244 98.161 68.308 ;
			RECT	98.297 68.244 98.329 68.308 ;
			RECT	98.465 68.244 98.497 68.308 ;
			RECT	98.633 68.244 98.665 68.308 ;
			RECT	98.801 68.244 98.833 68.308 ;
			RECT	98.969 68.244 99.001 68.308 ;
			RECT	99.137 68.244 99.169 68.308 ;
			RECT	99.305 68.244 99.337 68.308 ;
			RECT	99.473 68.244 99.505 68.308 ;
			RECT	99.641 68.244 99.673 68.308 ;
			RECT	99.809 68.244 99.841 68.308 ;
			RECT	99.977 68.244 100.009 68.308 ;
			RECT	100.145 68.244 100.177 68.308 ;
			RECT	100.313 68.244 100.345 68.308 ;
			RECT	100.481 68.244 100.513 68.308 ;
			RECT	100.649 68.244 100.681 68.308 ;
			RECT	100.817 68.244 100.849 68.308 ;
			RECT	100.985 68.244 101.017 68.308 ;
			RECT	101.153 68.244 101.185 68.308 ;
			RECT	101.321 68.244 101.353 68.308 ;
			RECT	101.489 68.244 101.521 68.308 ;
			RECT	101.657 68.244 101.689 68.308 ;
			RECT	101.825 68.244 101.857 68.308 ;
			RECT	101.993 68.244 102.025 68.308 ;
			RECT	102.123 68.26 102.155 68.292 ;
			RECT	102.245 68.255 102.277 68.287 ;
			RECT	102.375 68.244 102.407 68.308 ;
			RECT	103.795 68.244 103.827 68.308 ;
			RECT	103.925 68.255 103.957 68.287 ;
			RECT	104.047 68.26 104.079 68.292 ;
			RECT	104.177 68.244 104.209 68.308 ;
			RECT	104.345 68.244 104.377 68.308 ;
			RECT	104.513 68.244 104.545 68.308 ;
			RECT	104.681 68.244 104.713 68.308 ;
			RECT	104.849 68.244 104.881 68.308 ;
			RECT	105.017 68.244 105.049 68.308 ;
			RECT	105.185 68.244 105.217 68.308 ;
			RECT	105.353 68.244 105.385 68.308 ;
			RECT	105.521 68.244 105.553 68.308 ;
			RECT	105.689 68.244 105.721 68.308 ;
			RECT	105.857 68.244 105.889 68.308 ;
			RECT	106.025 68.244 106.057 68.308 ;
			RECT	106.193 68.244 106.225 68.308 ;
			RECT	106.361 68.244 106.393 68.308 ;
			RECT	106.529 68.244 106.561 68.308 ;
			RECT	106.697 68.244 106.729 68.308 ;
			RECT	106.865 68.244 106.897 68.308 ;
			RECT	107.033 68.244 107.065 68.308 ;
			RECT	107.201 68.244 107.233 68.308 ;
			RECT	107.369 68.244 107.401 68.308 ;
			RECT	107.537 68.244 107.569 68.308 ;
			RECT	107.705 68.244 107.737 68.308 ;
			RECT	107.873 68.244 107.905 68.308 ;
			RECT	108.041 68.244 108.073 68.308 ;
			RECT	108.209 68.244 108.241 68.308 ;
			RECT	108.377 68.244 108.409 68.308 ;
			RECT	108.545 68.244 108.577 68.308 ;
			RECT	108.713 68.244 108.745 68.308 ;
			RECT	108.881 68.244 108.913 68.308 ;
			RECT	109.049 68.244 109.081 68.308 ;
			RECT	109.217 68.244 109.249 68.308 ;
			RECT	109.385 68.244 109.417 68.308 ;
			RECT	109.553 68.244 109.585 68.308 ;
			RECT	109.721 68.244 109.753 68.308 ;
			RECT	109.889 68.244 109.921 68.308 ;
			RECT	110.057 68.244 110.089 68.308 ;
			RECT	110.225 68.244 110.257 68.308 ;
			RECT	110.393 68.244 110.425 68.308 ;
			RECT	110.561 68.244 110.593 68.308 ;
			RECT	110.729 68.244 110.761 68.308 ;
			RECT	110.897 68.244 110.929 68.308 ;
			RECT	111.065 68.244 111.097 68.308 ;
			RECT	111.233 68.244 111.265 68.308 ;
			RECT	111.401 68.244 111.433 68.308 ;
			RECT	111.569 68.244 111.601 68.308 ;
			RECT	111.737 68.244 111.769 68.308 ;
			RECT	111.905 68.244 111.937 68.308 ;
			RECT	112.073 68.244 112.105 68.308 ;
			RECT	112.241 68.244 112.273 68.308 ;
			RECT	112.409 68.244 112.441 68.308 ;
			RECT	112.577 68.244 112.609 68.308 ;
			RECT	112.745 68.244 112.777 68.308 ;
			RECT	112.913 68.244 112.945 68.308 ;
			RECT	113.081 68.244 113.113 68.308 ;
			RECT	113.249 68.244 113.281 68.308 ;
			RECT	113.417 68.244 113.449 68.308 ;
			RECT	113.585 68.244 113.617 68.308 ;
			RECT	113.753 68.244 113.785 68.308 ;
			RECT	113.921 68.244 113.953 68.308 ;
			RECT	114.089 68.244 114.121 68.308 ;
			RECT	114.257 68.244 114.289 68.308 ;
			RECT	114.425 68.244 114.457 68.308 ;
			RECT	114.593 68.244 114.625 68.308 ;
			RECT	114.761 68.244 114.793 68.308 ;
			RECT	114.929 68.244 114.961 68.308 ;
			RECT	115.097 68.244 115.129 68.308 ;
			RECT	115.265 68.244 115.297 68.308 ;
			RECT	115.433 68.244 115.465 68.308 ;
			RECT	115.601 68.244 115.633 68.308 ;
			RECT	115.769 68.244 115.801 68.308 ;
			RECT	115.937 68.244 115.969 68.308 ;
			RECT	116.105 68.244 116.137 68.308 ;
			RECT	116.273 68.244 116.305 68.308 ;
			RECT	116.441 68.244 116.473 68.308 ;
			RECT	116.609 68.244 116.641 68.308 ;
			RECT	116.777 68.244 116.809 68.308 ;
			RECT	116.945 68.244 116.977 68.308 ;
			RECT	117.113 68.244 117.145 68.308 ;
			RECT	117.281 68.244 117.313 68.308 ;
			RECT	117.449 68.244 117.481 68.308 ;
			RECT	117.617 68.244 117.649 68.308 ;
			RECT	117.785 68.244 117.817 68.308 ;
			RECT	117.953 68.244 117.985 68.308 ;
			RECT	118.121 68.244 118.153 68.308 ;
			RECT	118.289 68.244 118.321 68.308 ;
			RECT	118.457 68.244 118.489 68.308 ;
			RECT	118.625 68.244 118.657 68.308 ;
			RECT	118.793 68.244 118.825 68.308 ;
			RECT	118.961 68.244 118.993 68.308 ;
			RECT	119.129 68.244 119.161 68.308 ;
			RECT	119.297 68.244 119.329 68.308 ;
			RECT	119.465 68.244 119.497 68.308 ;
			RECT	119.633 68.244 119.665 68.308 ;
			RECT	119.801 68.244 119.833 68.308 ;
			RECT	119.969 68.244 120.001 68.308 ;
			RECT	120.137 68.244 120.169 68.308 ;
			RECT	120.305 68.244 120.337 68.308 ;
			RECT	120.473 68.244 120.505 68.308 ;
			RECT	120.641 68.244 120.673 68.308 ;
			RECT	120.809 68.244 120.841 68.308 ;
			RECT	120.977 68.244 121.009 68.308 ;
			RECT	121.145 68.244 121.177 68.308 ;
			RECT	121.313 68.244 121.345 68.308 ;
			RECT	121.481 68.244 121.513 68.308 ;
			RECT	121.649 68.244 121.681 68.308 ;
			RECT	121.817 68.244 121.849 68.308 ;
			RECT	121.985 68.244 122.017 68.308 ;
			RECT	122.153 68.244 122.185 68.308 ;
			RECT	122.321 68.244 122.353 68.308 ;
			RECT	122.489 68.244 122.521 68.308 ;
			RECT	122.657 68.244 122.689 68.308 ;
			RECT	122.825 68.244 122.857 68.308 ;
			RECT	122.993 68.244 123.025 68.308 ;
			RECT	123.161 68.244 123.193 68.308 ;
			RECT	123.329 68.244 123.361 68.308 ;
			RECT	123.497 68.244 123.529 68.308 ;
			RECT	123.665 68.244 123.697 68.308 ;
			RECT	123.833 68.244 123.865 68.308 ;
			RECT	124.001 68.244 124.033 68.308 ;
			RECT	124.169 68.244 124.201 68.308 ;
			RECT	124.337 68.244 124.369 68.308 ;
			RECT	124.505 68.244 124.537 68.308 ;
			RECT	124.673 68.244 124.705 68.308 ;
			RECT	124.841 68.244 124.873 68.308 ;
			RECT	125.009 68.244 125.041 68.308 ;
			RECT	125.177 68.244 125.209 68.308 ;
			RECT	125.345 68.244 125.377 68.308 ;
			RECT	125.513 68.244 125.545 68.308 ;
			RECT	125.681 68.244 125.713 68.308 ;
			RECT	125.849 68.244 125.881 68.308 ;
			RECT	126.017 68.244 126.049 68.308 ;
			RECT	126.185 68.244 126.217 68.308 ;
			RECT	126.353 68.244 126.385 68.308 ;
			RECT	126.521 68.244 126.553 68.308 ;
			RECT	126.689 68.244 126.721 68.308 ;
			RECT	126.857 68.244 126.889 68.308 ;
			RECT	127.025 68.244 127.057 68.308 ;
			RECT	127.193 68.244 127.225 68.308 ;
			RECT	127.361 68.244 127.393 68.308 ;
			RECT	127.529 68.244 127.561 68.308 ;
			RECT	127.697 68.244 127.729 68.308 ;
			RECT	127.865 68.244 127.897 68.308 ;
			RECT	128.033 68.244 128.065 68.308 ;
			RECT	128.201 68.244 128.233 68.308 ;
			RECT	128.369 68.244 128.401 68.308 ;
			RECT	128.537 68.244 128.569 68.308 ;
			RECT	128.705 68.244 128.737 68.308 ;
			RECT	128.873 68.244 128.905 68.308 ;
			RECT	129.041 68.244 129.073 68.308 ;
			RECT	129.209 68.244 129.241 68.308 ;
			RECT	129.377 68.244 129.409 68.308 ;
			RECT	129.545 68.244 129.577 68.308 ;
			RECT	129.713 68.244 129.745 68.308 ;
			RECT	129.881 68.244 129.913 68.308 ;
			RECT	130.049 68.244 130.081 68.308 ;
			RECT	130.217 68.244 130.249 68.308 ;
			RECT	130.385 68.244 130.417 68.308 ;
			RECT	130.553 68.244 130.585 68.308 ;
			RECT	130.721 68.244 130.753 68.308 ;
			RECT	130.889 68.244 130.921 68.308 ;
			RECT	131.057 68.244 131.089 68.308 ;
			RECT	131.225 68.244 131.257 68.308 ;
			RECT	131.393 68.244 131.425 68.308 ;
			RECT	131.561 68.244 131.593 68.308 ;
			RECT	131.729 68.244 131.761 68.308 ;
			RECT	131.897 68.244 131.929 68.308 ;
			RECT	132.065 68.244 132.097 68.308 ;
			RECT	132.233 68.244 132.265 68.308 ;
			RECT	132.401 68.244 132.433 68.308 ;
			RECT	132.569 68.244 132.601 68.308 ;
			RECT	132.737 68.244 132.769 68.308 ;
			RECT	132.905 68.244 132.937 68.308 ;
			RECT	133.073 68.244 133.105 68.308 ;
			RECT	133.241 68.244 133.273 68.308 ;
			RECT	133.409 68.244 133.441 68.308 ;
			RECT	133.577 68.244 133.609 68.308 ;
			RECT	133.745 68.244 133.777 68.308 ;
			RECT	133.913 68.244 133.945 68.308 ;
			RECT	134.081 68.244 134.113 68.308 ;
			RECT	134.249 68.244 134.281 68.308 ;
			RECT	134.417 68.244 134.449 68.308 ;
			RECT	134.585 68.244 134.617 68.308 ;
			RECT	134.753 68.244 134.785 68.308 ;
			RECT	134.921 68.244 134.953 68.308 ;
			RECT	135.089 68.244 135.121 68.308 ;
			RECT	135.257 68.244 135.289 68.308 ;
			RECT	135.425 68.244 135.457 68.308 ;
			RECT	135.593 68.244 135.625 68.308 ;
			RECT	135.761 68.244 135.793 68.308 ;
			RECT	135.929 68.244 135.961 68.308 ;
			RECT	136.097 68.244 136.129 68.308 ;
			RECT	136.265 68.244 136.297 68.308 ;
			RECT	136.433 68.244 136.465 68.308 ;
			RECT	136.601 68.244 136.633 68.308 ;
			RECT	136.769 68.244 136.801 68.308 ;
			RECT	136.937 68.244 136.969 68.308 ;
			RECT	137.105 68.244 137.137 68.308 ;
			RECT	137.273 68.244 137.305 68.308 ;
			RECT	137.441 68.244 137.473 68.308 ;
			RECT	137.609 68.244 137.641 68.308 ;
			RECT	137.777 68.244 137.809 68.308 ;
			RECT	137.945 68.244 137.977 68.308 ;
			RECT	138.113 68.244 138.145 68.308 ;
			RECT	138.281 68.244 138.313 68.308 ;
			RECT	138.449 68.244 138.481 68.308 ;
			RECT	138.617 68.244 138.649 68.308 ;
			RECT	138.785 68.244 138.817 68.308 ;
			RECT	138.953 68.244 138.985 68.308 ;
			RECT	139.121 68.244 139.153 68.308 ;
			RECT	139.289 68.244 139.321 68.308 ;
			RECT	139.457 68.244 139.489 68.308 ;
			RECT	139.625 68.244 139.657 68.308 ;
			RECT	139.793 68.244 139.825 68.308 ;
			RECT	139.961 68.244 139.993 68.308 ;
			RECT	140.129 68.244 140.161 68.308 ;
			RECT	140.297 68.244 140.329 68.308 ;
			RECT	140.465 68.244 140.497 68.308 ;
			RECT	140.633 68.244 140.665 68.308 ;
			RECT	140.801 68.244 140.833 68.308 ;
			RECT	140.969 68.244 141.001 68.308 ;
			RECT	141.137 68.244 141.169 68.308 ;
			RECT	141.305 68.244 141.337 68.308 ;
			RECT	141.473 68.244 141.505 68.308 ;
			RECT	141.641 68.244 141.673 68.308 ;
			RECT	141.809 68.244 141.841 68.308 ;
			RECT	141.977 68.244 142.009 68.308 ;
			RECT	142.145 68.244 142.177 68.308 ;
			RECT	142.313 68.244 142.345 68.308 ;
			RECT	142.481 68.244 142.513 68.308 ;
			RECT	142.649 68.244 142.681 68.308 ;
			RECT	142.817 68.244 142.849 68.308 ;
			RECT	142.985 68.244 143.017 68.308 ;
			RECT	143.153 68.244 143.185 68.308 ;
			RECT	143.321 68.244 143.353 68.308 ;
			RECT	143.489 68.244 143.521 68.308 ;
			RECT	143.657 68.244 143.689 68.308 ;
			RECT	143.825 68.244 143.857 68.308 ;
			RECT	143.993 68.244 144.025 68.308 ;
			RECT	144.161 68.244 144.193 68.308 ;
			RECT	144.329 68.244 144.361 68.308 ;
			RECT	144.497 68.244 144.529 68.308 ;
			RECT	144.665 68.244 144.697 68.308 ;
			RECT	144.833 68.244 144.865 68.308 ;
			RECT	145.001 68.244 145.033 68.308 ;
			RECT	145.169 68.244 145.201 68.308 ;
			RECT	145.337 68.244 145.369 68.308 ;
			RECT	145.505 68.244 145.537 68.308 ;
			RECT	145.673 68.244 145.705 68.308 ;
			RECT	145.841 68.244 145.873 68.308 ;
			RECT	146.009 68.244 146.041 68.308 ;
			RECT	146.177 68.244 146.209 68.308 ;
			RECT	146.345 68.244 146.377 68.308 ;
			RECT	146.513 68.244 146.545 68.308 ;
			RECT	146.681 68.244 146.713 68.308 ;
			RECT	146.849 68.244 146.881 68.308 ;
			RECT	147.017 68.244 147.049 68.308 ;
			RECT	147.185 68.244 147.217 68.308 ;
			RECT	147.316 68.26 147.348 68.292 ;
			RECT	147.437 68.26 147.469 68.292 ;
			RECT	147.567 68.244 147.599 68.308 ;
			RECT	149.879 68.244 149.911 68.308 ;
			RECT	151.13 68.244 151.194 68.308 ;
			RECT	151.81 68.244 151.842 68.308 ;
			RECT	152.249 68.244 152.281 68.308 ;
			RECT	153.56 68.244 153.624 68.308 ;
			RECT	156.601 68.244 156.633 68.308 ;
			RECT	156.731 68.26 156.763 68.292 ;
			RECT	156.852 68.26 156.884 68.292 ;
			RECT	156.983 68.244 157.015 68.308 ;
			RECT	157.151 68.244 157.183 68.308 ;
			RECT	157.319 68.244 157.351 68.308 ;
			RECT	157.487 68.244 157.519 68.308 ;
			RECT	157.655 68.244 157.687 68.308 ;
			RECT	157.823 68.244 157.855 68.308 ;
			RECT	157.991 68.244 158.023 68.308 ;
			RECT	158.159 68.244 158.191 68.308 ;
			RECT	158.327 68.244 158.359 68.308 ;
			RECT	158.495 68.244 158.527 68.308 ;
			RECT	158.663 68.244 158.695 68.308 ;
			RECT	158.831 68.244 158.863 68.308 ;
			RECT	158.999 68.244 159.031 68.308 ;
			RECT	159.167 68.244 159.199 68.308 ;
			RECT	159.335 68.244 159.367 68.308 ;
			RECT	159.503 68.244 159.535 68.308 ;
			RECT	159.671 68.244 159.703 68.308 ;
			RECT	159.839 68.244 159.871 68.308 ;
			RECT	160.007 68.244 160.039 68.308 ;
			RECT	160.175 68.244 160.207 68.308 ;
			RECT	160.343 68.244 160.375 68.308 ;
			RECT	160.511 68.244 160.543 68.308 ;
			RECT	160.679 68.244 160.711 68.308 ;
			RECT	160.847 68.244 160.879 68.308 ;
			RECT	161.015 68.244 161.047 68.308 ;
			RECT	161.183 68.244 161.215 68.308 ;
			RECT	161.351 68.244 161.383 68.308 ;
			RECT	161.519 68.244 161.551 68.308 ;
			RECT	161.687 68.244 161.719 68.308 ;
			RECT	161.855 68.244 161.887 68.308 ;
			RECT	162.023 68.244 162.055 68.308 ;
			RECT	162.191 68.244 162.223 68.308 ;
			RECT	162.359 68.244 162.391 68.308 ;
			RECT	162.527 68.244 162.559 68.308 ;
			RECT	162.695 68.244 162.727 68.308 ;
			RECT	162.863 68.244 162.895 68.308 ;
			RECT	163.031 68.244 163.063 68.308 ;
			RECT	163.199 68.244 163.231 68.308 ;
			RECT	163.367 68.244 163.399 68.308 ;
			RECT	163.535 68.244 163.567 68.308 ;
			RECT	163.703 68.244 163.735 68.308 ;
			RECT	163.871 68.244 163.903 68.308 ;
			RECT	164.039 68.244 164.071 68.308 ;
			RECT	164.207 68.244 164.239 68.308 ;
			RECT	164.375 68.244 164.407 68.308 ;
			RECT	164.543 68.244 164.575 68.308 ;
			RECT	164.711 68.244 164.743 68.308 ;
			RECT	164.879 68.244 164.911 68.308 ;
			RECT	165.047 68.244 165.079 68.308 ;
			RECT	165.215 68.244 165.247 68.308 ;
			RECT	165.383 68.244 165.415 68.308 ;
			RECT	165.551 68.244 165.583 68.308 ;
			RECT	165.719 68.244 165.751 68.308 ;
			RECT	165.887 68.244 165.919 68.308 ;
			RECT	166.055 68.244 166.087 68.308 ;
			RECT	166.223 68.244 166.255 68.308 ;
			RECT	166.391 68.244 166.423 68.308 ;
			RECT	166.559 68.244 166.591 68.308 ;
			RECT	166.727 68.244 166.759 68.308 ;
			RECT	166.895 68.244 166.927 68.308 ;
			RECT	167.063 68.244 167.095 68.308 ;
			RECT	167.231 68.244 167.263 68.308 ;
			RECT	167.399 68.244 167.431 68.308 ;
			RECT	167.567 68.244 167.599 68.308 ;
			RECT	167.735 68.244 167.767 68.308 ;
			RECT	167.903 68.244 167.935 68.308 ;
			RECT	168.071 68.244 168.103 68.308 ;
			RECT	168.239 68.244 168.271 68.308 ;
			RECT	168.407 68.244 168.439 68.308 ;
			RECT	168.575 68.244 168.607 68.308 ;
			RECT	168.743 68.244 168.775 68.308 ;
			RECT	168.911 68.244 168.943 68.308 ;
			RECT	169.079 68.244 169.111 68.308 ;
			RECT	169.247 68.244 169.279 68.308 ;
			RECT	169.415 68.244 169.447 68.308 ;
			RECT	169.583 68.244 169.615 68.308 ;
			RECT	169.751 68.244 169.783 68.308 ;
			RECT	169.919 68.244 169.951 68.308 ;
			RECT	170.087 68.244 170.119 68.308 ;
			RECT	170.255 68.244 170.287 68.308 ;
			RECT	170.423 68.244 170.455 68.308 ;
			RECT	170.591 68.244 170.623 68.308 ;
			RECT	170.759 68.244 170.791 68.308 ;
			RECT	170.927 68.244 170.959 68.308 ;
			RECT	171.095 68.244 171.127 68.308 ;
			RECT	171.263 68.244 171.295 68.308 ;
			RECT	171.431 68.244 171.463 68.308 ;
			RECT	171.599 68.244 171.631 68.308 ;
			RECT	171.767 68.244 171.799 68.308 ;
			RECT	171.935 68.244 171.967 68.308 ;
			RECT	172.103 68.244 172.135 68.308 ;
			RECT	172.271 68.244 172.303 68.308 ;
			RECT	172.439 68.244 172.471 68.308 ;
			RECT	172.607 68.244 172.639 68.308 ;
			RECT	172.775 68.244 172.807 68.308 ;
			RECT	172.943 68.244 172.975 68.308 ;
			RECT	173.111 68.244 173.143 68.308 ;
			RECT	173.279 68.244 173.311 68.308 ;
			RECT	173.447 68.244 173.479 68.308 ;
			RECT	173.615 68.244 173.647 68.308 ;
			RECT	173.783 68.244 173.815 68.308 ;
			RECT	173.951 68.244 173.983 68.308 ;
			RECT	174.119 68.244 174.151 68.308 ;
			RECT	174.287 68.244 174.319 68.308 ;
			RECT	174.455 68.244 174.487 68.308 ;
			RECT	174.623 68.244 174.655 68.308 ;
			RECT	174.791 68.244 174.823 68.308 ;
			RECT	174.959 68.244 174.991 68.308 ;
			RECT	175.127 68.244 175.159 68.308 ;
			RECT	175.295 68.244 175.327 68.308 ;
			RECT	175.463 68.244 175.495 68.308 ;
			RECT	175.631 68.244 175.663 68.308 ;
			RECT	175.799 68.244 175.831 68.308 ;
			RECT	175.967 68.244 175.999 68.308 ;
			RECT	176.135 68.244 176.167 68.308 ;
			RECT	176.303 68.244 176.335 68.308 ;
			RECT	176.471 68.244 176.503 68.308 ;
			RECT	176.639 68.244 176.671 68.308 ;
			RECT	176.807 68.244 176.839 68.308 ;
			RECT	176.975 68.244 177.007 68.308 ;
			RECT	177.143 68.244 177.175 68.308 ;
			RECT	177.311 68.244 177.343 68.308 ;
			RECT	177.479 68.244 177.511 68.308 ;
			RECT	177.647 68.244 177.679 68.308 ;
			RECT	177.815 68.244 177.847 68.308 ;
			RECT	177.983 68.244 178.015 68.308 ;
			RECT	178.151 68.244 178.183 68.308 ;
			RECT	178.319 68.244 178.351 68.308 ;
			RECT	178.487 68.244 178.519 68.308 ;
			RECT	178.655 68.244 178.687 68.308 ;
			RECT	178.823 68.244 178.855 68.308 ;
			RECT	178.991 68.244 179.023 68.308 ;
			RECT	179.159 68.244 179.191 68.308 ;
			RECT	179.327 68.244 179.359 68.308 ;
			RECT	179.495 68.244 179.527 68.308 ;
			RECT	179.663 68.244 179.695 68.308 ;
			RECT	179.831 68.244 179.863 68.308 ;
			RECT	179.999 68.244 180.031 68.308 ;
			RECT	180.167 68.244 180.199 68.308 ;
			RECT	180.335 68.244 180.367 68.308 ;
			RECT	180.503 68.244 180.535 68.308 ;
			RECT	180.671 68.244 180.703 68.308 ;
			RECT	180.839 68.244 180.871 68.308 ;
			RECT	181.007 68.244 181.039 68.308 ;
			RECT	181.175 68.244 181.207 68.308 ;
			RECT	181.343 68.244 181.375 68.308 ;
			RECT	181.511 68.244 181.543 68.308 ;
			RECT	181.679 68.244 181.711 68.308 ;
			RECT	181.847 68.244 181.879 68.308 ;
			RECT	182.015 68.244 182.047 68.308 ;
			RECT	182.183 68.244 182.215 68.308 ;
			RECT	182.351 68.244 182.383 68.308 ;
			RECT	182.519 68.244 182.551 68.308 ;
			RECT	182.687 68.244 182.719 68.308 ;
			RECT	182.855 68.244 182.887 68.308 ;
			RECT	183.023 68.244 183.055 68.308 ;
			RECT	183.191 68.244 183.223 68.308 ;
			RECT	183.359 68.244 183.391 68.308 ;
			RECT	183.527 68.244 183.559 68.308 ;
			RECT	183.695 68.244 183.727 68.308 ;
			RECT	183.863 68.244 183.895 68.308 ;
			RECT	184.031 68.244 184.063 68.308 ;
			RECT	184.199 68.244 184.231 68.308 ;
			RECT	184.367 68.244 184.399 68.308 ;
			RECT	184.535 68.244 184.567 68.308 ;
			RECT	184.703 68.244 184.735 68.308 ;
			RECT	184.871 68.244 184.903 68.308 ;
			RECT	185.039 68.244 185.071 68.308 ;
			RECT	185.207 68.244 185.239 68.308 ;
			RECT	185.375 68.244 185.407 68.308 ;
			RECT	185.543 68.244 185.575 68.308 ;
			RECT	185.711 68.244 185.743 68.308 ;
			RECT	185.879 68.244 185.911 68.308 ;
			RECT	186.047 68.244 186.079 68.308 ;
			RECT	186.215 68.244 186.247 68.308 ;
			RECT	186.383 68.244 186.415 68.308 ;
			RECT	186.551 68.244 186.583 68.308 ;
			RECT	186.719 68.244 186.751 68.308 ;
			RECT	186.887 68.244 186.919 68.308 ;
			RECT	187.055 68.244 187.087 68.308 ;
			RECT	187.223 68.244 187.255 68.308 ;
			RECT	187.391 68.244 187.423 68.308 ;
			RECT	187.559 68.244 187.591 68.308 ;
			RECT	187.727 68.244 187.759 68.308 ;
			RECT	187.895 68.244 187.927 68.308 ;
			RECT	188.063 68.244 188.095 68.308 ;
			RECT	188.231 68.244 188.263 68.308 ;
			RECT	188.399 68.244 188.431 68.308 ;
			RECT	188.567 68.244 188.599 68.308 ;
			RECT	188.735 68.244 188.767 68.308 ;
			RECT	188.903 68.244 188.935 68.308 ;
			RECT	189.071 68.244 189.103 68.308 ;
			RECT	189.239 68.244 189.271 68.308 ;
			RECT	189.407 68.244 189.439 68.308 ;
			RECT	189.575 68.244 189.607 68.308 ;
			RECT	189.743 68.244 189.775 68.308 ;
			RECT	189.911 68.244 189.943 68.308 ;
			RECT	190.079 68.244 190.111 68.308 ;
			RECT	190.247 68.244 190.279 68.308 ;
			RECT	190.415 68.244 190.447 68.308 ;
			RECT	190.583 68.244 190.615 68.308 ;
			RECT	190.751 68.244 190.783 68.308 ;
			RECT	190.919 68.244 190.951 68.308 ;
			RECT	191.087 68.244 191.119 68.308 ;
			RECT	191.255 68.244 191.287 68.308 ;
			RECT	191.423 68.244 191.455 68.308 ;
			RECT	191.591 68.244 191.623 68.308 ;
			RECT	191.759 68.244 191.791 68.308 ;
			RECT	191.927 68.244 191.959 68.308 ;
			RECT	192.095 68.244 192.127 68.308 ;
			RECT	192.263 68.244 192.295 68.308 ;
			RECT	192.431 68.244 192.463 68.308 ;
			RECT	192.599 68.244 192.631 68.308 ;
			RECT	192.767 68.244 192.799 68.308 ;
			RECT	192.935 68.244 192.967 68.308 ;
			RECT	193.103 68.244 193.135 68.308 ;
			RECT	193.271 68.244 193.303 68.308 ;
			RECT	193.439 68.244 193.471 68.308 ;
			RECT	193.607 68.244 193.639 68.308 ;
			RECT	193.775 68.244 193.807 68.308 ;
			RECT	193.943 68.244 193.975 68.308 ;
			RECT	194.111 68.244 194.143 68.308 ;
			RECT	194.279 68.244 194.311 68.308 ;
			RECT	194.447 68.244 194.479 68.308 ;
			RECT	194.615 68.244 194.647 68.308 ;
			RECT	194.783 68.244 194.815 68.308 ;
			RECT	194.951 68.244 194.983 68.308 ;
			RECT	195.119 68.244 195.151 68.308 ;
			RECT	195.287 68.244 195.319 68.308 ;
			RECT	195.455 68.244 195.487 68.308 ;
			RECT	195.623 68.244 195.655 68.308 ;
			RECT	195.791 68.244 195.823 68.308 ;
			RECT	195.959 68.244 195.991 68.308 ;
			RECT	196.127 68.244 196.159 68.308 ;
			RECT	196.295 68.244 196.327 68.308 ;
			RECT	196.463 68.244 196.495 68.308 ;
			RECT	196.631 68.244 196.663 68.308 ;
			RECT	196.799 68.244 196.831 68.308 ;
			RECT	196.967 68.244 196.999 68.308 ;
			RECT	197.135 68.244 197.167 68.308 ;
			RECT	197.303 68.244 197.335 68.308 ;
			RECT	197.471 68.244 197.503 68.308 ;
			RECT	197.639 68.244 197.671 68.308 ;
			RECT	197.807 68.244 197.839 68.308 ;
			RECT	197.975 68.244 198.007 68.308 ;
			RECT	198.143 68.244 198.175 68.308 ;
			RECT	198.311 68.244 198.343 68.308 ;
			RECT	198.479 68.244 198.511 68.308 ;
			RECT	198.647 68.244 198.679 68.308 ;
			RECT	198.815 68.244 198.847 68.308 ;
			RECT	198.983 68.244 199.015 68.308 ;
			RECT	199.151 68.244 199.183 68.308 ;
			RECT	199.319 68.244 199.351 68.308 ;
			RECT	199.487 68.244 199.519 68.308 ;
			RECT	199.655 68.244 199.687 68.308 ;
			RECT	199.823 68.244 199.855 68.308 ;
			RECT	199.991 68.244 200.023 68.308 ;
			RECT	200.121 68.26 200.153 68.292 ;
			RECT	200.243 68.255 200.275 68.287 ;
			RECT	200.373 68.244 200.405 68.308 ;
			RECT	200.9 68.244 200.932 68.308 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 66.296 201.665 66.416 ;
			LAYER	J3 ;
			RECT	0.755 66.324 0.787 66.388 ;
			RECT	1.645 66.324 1.709 66.388 ;
			RECT	2.323 66.324 2.387 66.388 ;
			RECT	3.438 66.324 3.47 66.388 ;
			RECT	3.585 66.324 3.617 66.388 ;
			RECT	4.195 66.324 4.227 66.388 ;
			RECT	4.72 66.324 4.752 66.388 ;
			RECT	4.944 66.324 5.008 66.388 ;
			RECT	5.267 66.324 5.299 66.388 ;
			RECT	5.797 66.324 5.829 66.388 ;
			RECT	5.927 66.335 5.959 66.367 ;
			RECT	6.049 66.34 6.081 66.372 ;
			RECT	6.179 66.324 6.211 66.388 ;
			RECT	6.347 66.324 6.379 66.388 ;
			RECT	6.515 66.324 6.547 66.388 ;
			RECT	6.683 66.324 6.715 66.388 ;
			RECT	6.851 66.324 6.883 66.388 ;
			RECT	7.019 66.324 7.051 66.388 ;
			RECT	7.187 66.324 7.219 66.388 ;
			RECT	7.355 66.324 7.387 66.388 ;
			RECT	7.523 66.324 7.555 66.388 ;
			RECT	7.691 66.324 7.723 66.388 ;
			RECT	7.859 66.324 7.891 66.388 ;
			RECT	8.027 66.324 8.059 66.388 ;
			RECT	8.195 66.324 8.227 66.388 ;
			RECT	8.363 66.324 8.395 66.388 ;
			RECT	8.531 66.324 8.563 66.388 ;
			RECT	8.699 66.324 8.731 66.388 ;
			RECT	8.867 66.324 8.899 66.388 ;
			RECT	9.035 66.324 9.067 66.388 ;
			RECT	9.203 66.324 9.235 66.388 ;
			RECT	9.371 66.324 9.403 66.388 ;
			RECT	9.539 66.324 9.571 66.388 ;
			RECT	9.707 66.324 9.739 66.388 ;
			RECT	9.875 66.324 9.907 66.388 ;
			RECT	10.043 66.324 10.075 66.388 ;
			RECT	10.211 66.324 10.243 66.388 ;
			RECT	10.379 66.324 10.411 66.388 ;
			RECT	10.547 66.324 10.579 66.388 ;
			RECT	10.715 66.324 10.747 66.388 ;
			RECT	10.883 66.324 10.915 66.388 ;
			RECT	11.051 66.324 11.083 66.388 ;
			RECT	11.219 66.324 11.251 66.388 ;
			RECT	11.387 66.324 11.419 66.388 ;
			RECT	11.555 66.324 11.587 66.388 ;
			RECT	11.723 66.324 11.755 66.388 ;
			RECT	11.891 66.324 11.923 66.388 ;
			RECT	12.059 66.324 12.091 66.388 ;
			RECT	12.227 66.324 12.259 66.388 ;
			RECT	12.395 66.324 12.427 66.388 ;
			RECT	12.563 66.324 12.595 66.388 ;
			RECT	12.731 66.324 12.763 66.388 ;
			RECT	12.899 66.324 12.931 66.388 ;
			RECT	13.067 66.324 13.099 66.388 ;
			RECT	13.235 66.324 13.267 66.388 ;
			RECT	13.403 66.324 13.435 66.388 ;
			RECT	13.571 66.324 13.603 66.388 ;
			RECT	13.739 66.324 13.771 66.388 ;
			RECT	13.907 66.324 13.939 66.388 ;
			RECT	14.075 66.324 14.107 66.388 ;
			RECT	14.243 66.324 14.275 66.388 ;
			RECT	14.411 66.324 14.443 66.388 ;
			RECT	14.579 66.324 14.611 66.388 ;
			RECT	14.747 66.324 14.779 66.388 ;
			RECT	14.915 66.324 14.947 66.388 ;
			RECT	15.083 66.324 15.115 66.388 ;
			RECT	15.251 66.324 15.283 66.388 ;
			RECT	15.419 66.324 15.451 66.388 ;
			RECT	15.587 66.324 15.619 66.388 ;
			RECT	15.755 66.324 15.787 66.388 ;
			RECT	15.923 66.324 15.955 66.388 ;
			RECT	16.091 66.324 16.123 66.388 ;
			RECT	16.259 66.324 16.291 66.388 ;
			RECT	16.427 66.324 16.459 66.388 ;
			RECT	16.595 66.324 16.627 66.388 ;
			RECT	16.763 66.324 16.795 66.388 ;
			RECT	16.931 66.324 16.963 66.388 ;
			RECT	17.099 66.324 17.131 66.388 ;
			RECT	17.267 66.324 17.299 66.388 ;
			RECT	17.435 66.324 17.467 66.388 ;
			RECT	17.603 66.324 17.635 66.388 ;
			RECT	17.771 66.324 17.803 66.388 ;
			RECT	17.939 66.324 17.971 66.388 ;
			RECT	18.107 66.324 18.139 66.388 ;
			RECT	18.275 66.324 18.307 66.388 ;
			RECT	18.443 66.324 18.475 66.388 ;
			RECT	18.611 66.324 18.643 66.388 ;
			RECT	18.779 66.324 18.811 66.388 ;
			RECT	18.947 66.324 18.979 66.388 ;
			RECT	19.115 66.324 19.147 66.388 ;
			RECT	19.283 66.324 19.315 66.388 ;
			RECT	19.451 66.324 19.483 66.388 ;
			RECT	19.619 66.324 19.651 66.388 ;
			RECT	19.787 66.324 19.819 66.388 ;
			RECT	19.955 66.324 19.987 66.388 ;
			RECT	20.123 66.324 20.155 66.388 ;
			RECT	20.291 66.324 20.323 66.388 ;
			RECT	20.459 66.324 20.491 66.388 ;
			RECT	20.627 66.324 20.659 66.388 ;
			RECT	20.795 66.324 20.827 66.388 ;
			RECT	20.963 66.324 20.995 66.388 ;
			RECT	21.131 66.324 21.163 66.388 ;
			RECT	21.299 66.324 21.331 66.388 ;
			RECT	21.467 66.324 21.499 66.388 ;
			RECT	21.635 66.324 21.667 66.388 ;
			RECT	21.803 66.324 21.835 66.388 ;
			RECT	21.971 66.324 22.003 66.388 ;
			RECT	22.139 66.324 22.171 66.388 ;
			RECT	22.307 66.324 22.339 66.388 ;
			RECT	22.475 66.324 22.507 66.388 ;
			RECT	22.643 66.324 22.675 66.388 ;
			RECT	22.811 66.324 22.843 66.388 ;
			RECT	22.979 66.324 23.011 66.388 ;
			RECT	23.147 66.324 23.179 66.388 ;
			RECT	23.315 66.324 23.347 66.388 ;
			RECT	23.483 66.324 23.515 66.388 ;
			RECT	23.651 66.324 23.683 66.388 ;
			RECT	23.819 66.324 23.851 66.388 ;
			RECT	23.987 66.324 24.019 66.388 ;
			RECT	24.155 66.324 24.187 66.388 ;
			RECT	24.323 66.324 24.355 66.388 ;
			RECT	24.491 66.324 24.523 66.388 ;
			RECT	24.659 66.324 24.691 66.388 ;
			RECT	24.827 66.324 24.859 66.388 ;
			RECT	24.995 66.324 25.027 66.388 ;
			RECT	25.163 66.324 25.195 66.388 ;
			RECT	25.331 66.324 25.363 66.388 ;
			RECT	25.499 66.324 25.531 66.388 ;
			RECT	25.667 66.324 25.699 66.388 ;
			RECT	25.835 66.324 25.867 66.388 ;
			RECT	26.003 66.324 26.035 66.388 ;
			RECT	26.171 66.324 26.203 66.388 ;
			RECT	26.339 66.324 26.371 66.388 ;
			RECT	26.507 66.324 26.539 66.388 ;
			RECT	26.675 66.324 26.707 66.388 ;
			RECT	26.843 66.324 26.875 66.388 ;
			RECT	27.011 66.324 27.043 66.388 ;
			RECT	27.179 66.324 27.211 66.388 ;
			RECT	27.347 66.324 27.379 66.388 ;
			RECT	27.515 66.324 27.547 66.388 ;
			RECT	27.683 66.324 27.715 66.388 ;
			RECT	27.851 66.324 27.883 66.388 ;
			RECT	28.019 66.324 28.051 66.388 ;
			RECT	28.187 66.324 28.219 66.388 ;
			RECT	28.355 66.324 28.387 66.388 ;
			RECT	28.523 66.324 28.555 66.388 ;
			RECT	28.691 66.324 28.723 66.388 ;
			RECT	28.859 66.324 28.891 66.388 ;
			RECT	29.027 66.324 29.059 66.388 ;
			RECT	29.195 66.324 29.227 66.388 ;
			RECT	29.363 66.324 29.395 66.388 ;
			RECT	29.531 66.324 29.563 66.388 ;
			RECT	29.699 66.324 29.731 66.388 ;
			RECT	29.867 66.324 29.899 66.388 ;
			RECT	30.035 66.324 30.067 66.388 ;
			RECT	30.203 66.324 30.235 66.388 ;
			RECT	30.371 66.324 30.403 66.388 ;
			RECT	30.539 66.324 30.571 66.388 ;
			RECT	30.707 66.324 30.739 66.388 ;
			RECT	30.875 66.324 30.907 66.388 ;
			RECT	31.043 66.324 31.075 66.388 ;
			RECT	31.211 66.324 31.243 66.388 ;
			RECT	31.379 66.324 31.411 66.388 ;
			RECT	31.547 66.324 31.579 66.388 ;
			RECT	31.715 66.324 31.747 66.388 ;
			RECT	31.883 66.324 31.915 66.388 ;
			RECT	32.051 66.324 32.083 66.388 ;
			RECT	32.219 66.324 32.251 66.388 ;
			RECT	32.387 66.324 32.419 66.388 ;
			RECT	32.555 66.324 32.587 66.388 ;
			RECT	32.723 66.324 32.755 66.388 ;
			RECT	32.891 66.324 32.923 66.388 ;
			RECT	33.059 66.324 33.091 66.388 ;
			RECT	33.227 66.324 33.259 66.388 ;
			RECT	33.395 66.324 33.427 66.388 ;
			RECT	33.563 66.324 33.595 66.388 ;
			RECT	33.731 66.324 33.763 66.388 ;
			RECT	33.899 66.324 33.931 66.388 ;
			RECT	34.067 66.324 34.099 66.388 ;
			RECT	34.235 66.324 34.267 66.388 ;
			RECT	34.403 66.324 34.435 66.388 ;
			RECT	34.571 66.324 34.603 66.388 ;
			RECT	34.739 66.324 34.771 66.388 ;
			RECT	34.907 66.324 34.939 66.388 ;
			RECT	35.075 66.324 35.107 66.388 ;
			RECT	35.243 66.324 35.275 66.388 ;
			RECT	35.411 66.324 35.443 66.388 ;
			RECT	35.579 66.324 35.611 66.388 ;
			RECT	35.747 66.324 35.779 66.388 ;
			RECT	35.915 66.324 35.947 66.388 ;
			RECT	36.083 66.324 36.115 66.388 ;
			RECT	36.251 66.324 36.283 66.388 ;
			RECT	36.419 66.324 36.451 66.388 ;
			RECT	36.587 66.324 36.619 66.388 ;
			RECT	36.755 66.324 36.787 66.388 ;
			RECT	36.923 66.324 36.955 66.388 ;
			RECT	37.091 66.324 37.123 66.388 ;
			RECT	37.259 66.324 37.291 66.388 ;
			RECT	37.427 66.324 37.459 66.388 ;
			RECT	37.595 66.324 37.627 66.388 ;
			RECT	37.763 66.324 37.795 66.388 ;
			RECT	37.931 66.324 37.963 66.388 ;
			RECT	38.099 66.324 38.131 66.388 ;
			RECT	38.267 66.324 38.299 66.388 ;
			RECT	38.435 66.324 38.467 66.388 ;
			RECT	38.603 66.324 38.635 66.388 ;
			RECT	38.771 66.324 38.803 66.388 ;
			RECT	38.939 66.324 38.971 66.388 ;
			RECT	39.107 66.324 39.139 66.388 ;
			RECT	39.275 66.324 39.307 66.388 ;
			RECT	39.443 66.324 39.475 66.388 ;
			RECT	39.611 66.324 39.643 66.388 ;
			RECT	39.779 66.324 39.811 66.388 ;
			RECT	39.947 66.324 39.979 66.388 ;
			RECT	40.115 66.324 40.147 66.388 ;
			RECT	40.283 66.324 40.315 66.388 ;
			RECT	40.451 66.324 40.483 66.388 ;
			RECT	40.619 66.324 40.651 66.388 ;
			RECT	40.787 66.324 40.819 66.388 ;
			RECT	40.955 66.324 40.987 66.388 ;
			RECT	41.123 66.324 41.155 66.388 ;
			RECT	41.291 66.324 41.323 66.388 ;
			RECT	41.459 66.324 41.491 66.388 ;
			RECT	41.627 66.324 41.659 66.388 ;
			RECT	41.795 66.324 41.827 66.388 ;
			RECT	41.963 66.324 41.995 66.388 ;
			RECT	42.131 66.324 42.163 66.388 ;
			RECT	42.299 66.324 42.331 66.388 ;
			RECT	42.467 66.324 42.499 66.388 ;
			RECT	42.635 66.324 42.667 66.388 ;
			RECT	42.803 66.324 42.835 66.388 ;
			RECT	42.971 66.324 43.003 66.388 ;
			RECT	43.139 66.324 43.171 66.388 ;
			RECT	43.307 66.324 43.339 66.388 ;
			RECT	43.475 66.324 43.507 66.388 ;
			RECT	43.643 66.324 43.675 66.388 ;
			RECT	43.811 66.324 43.843 66.388 ;
			RECT	43.979 66.324 44.011 66.388 ;
			RECT	44.147 66.324 44.179 66.388 ;
			RECT	44.315 66.324 44.347 66.388 ;
			RECT	44.483 66.324 44.515 66.388 ;
			RECT	44.651 66.324 44.683 66.388 ;
			RECT	44.819 66.324 44.851 66.388 ;
			RECT	44.987 66.324 45.019 66.388 ;
			RECT	45.155 66.324 45.187 66.388 ;
			RECT	45.323 66.324 45.355 66.388 ;
			RECT	45.491 66.324 45.523 66.388 ;
			RECT	45.659 66.324 45.691 66.388 ;
			RECT	45.827 66.324 45.859 66.388 ;
			RECT	45.995 66.324 46.027 66.388 ;
			RECT	46.163 66.324 46.195 66.388 ;
			RECT	46.331 66.324 46.363 66.388 ;
			RECT	46.499 66.324 46.531 66.388 ;
			RECT	46.667 66.324 46.699 66.388 ;
			RECT	46.835 66.324 46.867 66.388 ;
			RECT	47.003 66.324 47.035 66.388 ;
			RECT	47.171 66.324 47.203 66.388 ;
			RECT	47.339 66.324 47.371 66.388 ;
			RECT	47.507 66.324 47.539 66.388 ;
			RECT	47.675 66.324 47.707 66.388 ;
			RECT	47.843 66.324 47.875 66.388 ;
			RECT	48.011 66.324 48.043 66.388 ;
			RECT	48.179 66.324 48.211 66.388 ;
			RECT	48.347 66.324 48.379 66.388 ;
			RECT	48.515 66.324 48.547 66.388 ;
			RECT	48.683 66.324 48.715 66.388 ;
			RECT	48.851 66.324 48.883 66.388 ;
			RECT	49.019 66.324 49.051 66.388 ;
			RECT	49.187 66.324 49.219 66.388 ;
			RECT	49.318 66.34 49.35 66.372 ;
			RECT	49.439 66.34 49.471 66.372 ;
			RECT	49.569 66.324 49.601 66.388 ;
			RECT	51.881 66.324 51.913 66.388 ;
			RECT	53.132 66.324 53.196 66.388 ;
			RECT	53.812 66.324 53.844 66.388 ;
			RECT	54.251 66.324 54.283 66.388 ;
			RECT	55.562 66.324 55.626 66.388 ;
			RECT	58.603 66.324 58.635 66.388 ;
			RECT	58.733 66.34 58.765 66.372 ;
			RECT	58.854 66.34 58.886 66.372 ;
			RECT	58.985 66.324 59.017 66.388 ;
			RECT	59.153 66.324 59.185 66.388 ;
			RECT	59.321 66.324 59.353 66.388 ;
			RECT	59.489 66.324 59.521 66.388 ;
			RECT	59.657 66.324 59.689 66.388 ;
			RECT	59.825 66.324 59.857 66.388 ;
			RECT	59.993 66.324 60.025 66.388 ;
			RECT	60.161 66.324 60.193 66.388 ;
			RECT	60.329 66.324 60.361 66.388 ;
			RECT	60.497 66.324 60.529 66.388 ;
			RECT	60.665 66.324 60.697 66.388 ;
			RECT	60.833 66.324 60.865 66.388 ;
			RECT	61.001 66.324 61.033 66.388 ;
			RECT	61.169 66.324 61.201 66.388 ;
			RECT	61.337 66.324 61.369 66.388 ;
			RECT	61.505 66.324 61.537 66.388 ;
			RECT	61.673 66.324 61.705 66.388 ;
			RECT	61.841 66.324 61.873 66.388 ;
			RECT	62.009 66.324 62.041 66.388 ;
			RECT	62.177 66.324 62.209 66.388 ;
			RECT	62.345 66.324 62.377 66.388 ;
			RECT	62.513 66.324 62.545 66.388 ;
			RECT	62.681 66.324 62.713 66.388 ;
			RECT	62.849 66.324 62.881 66.388 ;
			RECT	63.017 66.324 63.049 66.388 ;
			RECT	63.185 66.324 63.217 66.388 ;
			RECT	63.353 66.324 63.385 66.388 ;
			RECT	63.521 66.324 63.553 66.388 ;
			RECT	63.689 66.324 63.721 66.388 ;
			RECT	63.857 66.324 63.889 66.388 ;
			RECT	64.025 66.324 64.057 66.388 ;
			RECT	64.193 66.324 64.225 66.388 ;
			RECT	64.361 66.324 64.393 66.388 ;
			RECT	64.529 66.324 64.561 66.388 ;
			RECT	64.697 66.324 64.729 66.388 ;
			RECT	64.865 66.324 64.897 66.388 ;
			RECT	65.033 66.324 65.065 66.388 ;
			RECT	65.201 66.324 65.233 66.388 ;
			RECT	65.369 66.324 65.401 66.388 ;
			RECT	65.537 66.324 65.569 66.388 ;
			RECT	65.705 66.324 65.737 66.388 ;
			RECT	65.873 66.324 65.905 66.388 ;
			RECT	66.041 66.324 66.073 66.388 ;
			RECT	66.209 66.324 66.241 66.388 ;
			RECT	66.377 66.324 66.409 66.388 ;
			RECT	66.545 66.324 66.577 66.388 ;
			RECT	66.713 66.324 66.745 66.388 ;
			RECT	66.881 66.324 66.913 66.388 ;
			RECT	67.049 66.324 67.081 66.388 ;
			RECT	67.217 66.324 67.249 66.388 ;
			RECT	67.385 66.324 67.417 66.388 ;
			RECT	67.553 66.324 67.585 66.388 ;
			RECT	67.721 66.324 67.753 66.388 ;
			RECT	67.889 66.324 67.921 66.388 ;
			RECT	68.057 66.324 68.089 66.388 ;
			RECT	68.225 66.324 68.257 66.388 ;
			RECT	68.393 66.324 68.425 66.388 ;
			RECT	68.561 66.324 68.593 66.388 ;
			RECT	68.729 66.324 68.761 66.388 ;
			RECT	68.897 66.324 68.929 66.388 ;
			RECT	69.065 66.324 69.097 66.388 ;
			RECT	69.233 66.324 69.265 66.388 ;
			RECT	69.401 66.324 69.433 66.388 ;
			RECT	69.569 66.324 69.601 66.388 ;
			RECT	69.737 66.324 69.769 66.388 ;
			RECT	69.905 66.324 69.937 66.388 ;
			RECT	70.073 66.324 70.105 66.388 ;
			RECT	70.241 66.324 70.273 66.388 ;
			RECT	70.409 66.324 70.441 66.388 ;
			RECT	70.577 66.324 70.609 66.388 ;
			RECT	70.745 66.324 70.777 66.388 ;
			RECT	70.913 66.324 70.945 66.388 ;
			RECT	71.081 66.324 71.113 66.388 ;
			RECT	71.249 66.324 71.281 66.388 ;
			RECT	71.417 66.324 71.449 66.388 ;
			RECT	71.585 66.324 71.617 66.388 ;
			RECT	71.753 66.324 71.785 66.388 ;
			RECT	71.921 66.324 71.953 66.388 ;
			RECT	72.089 66.324 72.121 66.388 ;
			RECT	72.257 66.324 72.289 66.388 ;
			RECT	72.425 66.324 72.457 66.388 ;
			RECT	72.593 66.324 72.625 66.388 ;
			RECT	72.761 66.324 72.793 66.388 ;
			RECT	72.929 66.324 72.961 66.388 ;
			RECT	73.097 66.324 73.129 66.388 ;
			RECT	73.265 66.324 73.297 66.388 ;
			RECT	73.433 66.324 73.465 66.388 ;
			RECT	73.601 66.324 73.633 66.388 ;
			RECT	73.769 66.324 73.801 66.388 ;
			RECT	73.937 66.324 73.969 66.388 ;
			RECT	74.105 66.324 74.137 66.388 ;
			RECT	74.273 66.324 74.305 66.388 ;
			RECT	74.441 66.324 74.473 66.388 ;
			RECT	74.609 66.324 74.641 66.388 ;
			RECT	74.777 66.324 74.809 66.388 ;
			RECT	74.945 66.324 74.977 66.388 ;
			RECT	75.113 66.324 75.145 66.388 ;
			RECT	75.281 66.324 75.313 66.388 ;
			RECT	75.449 66.324 75.481 66.388 ;
			RECT	75.617 66.324 75.649 66.388 ;
			RECT	75.785 66.324 75.817 66.388 ;
			RECT	75.953 66.324 75.985 66.388 ;
			RECT	76.121 66.324 76.153 66.388 ;
			RECT	76.289 66.324 76.321 66.388 ;
			RECT	76.457 66.324 76.489 66.388 ;
			RECT	76.625 66.324 76.657 66.388 ;
			RECT	76.793 66.324 76.825 66.388 ;
			RECT	76.961 66.324 76.993 66.388 ;
			RECT	77.129 66.324 77.161 66.388 ;
			RECT	77.297 66.324 77.329 66.388 ;
			RECT	77.465 66.324 77.497 66.388 ;
			RECT	77.633 66.324 77.665 66.388 ;
			RECT	77.801 66.324 77.833 66.388 ;
			RECT	77.969 66.324 78.001 66.388 ;
			RECT	78.137 66.324 78.169 66.388 ;
			RECT	78.305 66.324 78.337 66.388 ;
			RECT	78.473 66.324 78.505 66.388 ;
			RECT	78.641 66.324 78.673 66.388 ;
			RECT	78.809 66.324 78.841 66.388 ;
			RECT	78.977 66.324 79.009 66.388 ;
			RECT	79.145 66.324 79.177 66.388 ;
			RECT	79.313 66.324 79.345 66.388 ;
			RECT	79.481 66.324 79.513 66.388 ;
			RECT	79.649 66.324 79.681 66.388 ;
			RECT	79.817 66.324 79.849 66.388 ;
			RECT	79.985 66.324 80.017 66.388 ;
			RECT	80.153 66.324 80.185 66.388 ;
			RECT	80.321 66.324 80.353 66.388 ;
			RECT	80.489 66.324 80.521 66.388 ;
			RECT	80.657 66.324 80.689 66.388 ;
			RECT	80.825 66.324 80.857 66.388 ;
			RECT	80.993 66.324 81.025 66.388 ;
			RECT	81.161 66.324 81.193 66.388 ;
			RECT	81.329 66.324 81.361 66.388 ;
			RECT	81.497 66.324 81.529 66.388 ;
			RECT	81.665 66.324 81.697 66.388 ;
			RECT	81.833 66.324 81.865 66.388 ;
			RECT	82.001 66.324 82.033 66.388 ;
			RECT	82.169 66.324 82.201 66.388 ;
			RECT	82.337 66.324 82.369 66.388 ;
			RECT	82.505 66.324 82.537 66.388 ;
			RECT	82.673 66.324 82.705 66.388 ;
			RECT	82.841 66.324 82.873 66.388 ;
			RECT	83.009 66.324 83.041 66.388 ;
			RECT	83.177 66.324 83.209 66.388 ;
			RECT	83.345 66.324 83.377 66.388 ;
			RECT	83.513 66.324 83.545 66.388 ;
			RECT	83.681 66.324 83.713 66.388 ;
			RECT	83.849 66.324 83.881 66.388 ;
			RECT	84.017 66.324 84.049 66.388 ;
			RECT	84.185 66.324 84.217 66.388 ;
			RECT	84.353 66.324 84.385 66.388 ;
			RECT	84.521 66.324 84.553 66.388 ;
			RECT	84.689 66.324 84.721 66.388 ;
			RECT	84.857 66.324 84.889 66.388 ;
			RECT	85.025 66.324 85.057 66.388 ;
			RECT	85.193 66.324 85.225 66.388 ;
			RECT	85.361 66.324 85.393 66.388 ;
			RECT	85.529 66.324 85.561 66.388 ;
			RECT	85.697 66.324 85.729 66.388 ;
			RECT	85.865 66.324 85.897 66.388 ;
			RECT	86.033 66.324 86.065 66.388 ;
			RECT	86.201 66.324 86.233 66.388 ;
			RECT	86.369 66.324 86.401 66.388 ;
			RECT	86.537 66.324 86.569 66.388 ;
			RECT	86.705 66.324 86.737 66.388 ;
			RECT	86.873 66.324 86.905 66.388 ;
			RECT	87.041 66.324 87.073 66.388 ;
			RECT	87.209 66.324 87.241 66.388 ;
			RECT	87.377 66.324 87.409 66.388 ;
			RECT	87.545 66.324 87.577 66.388 ;
			RECT	87.713 66.324 87.745 66.388 ;
			RECT	87.881 66.324 87.913 66.388 ;
			RECT	88.049 66.324 88.081 66.388 ;
			RECT	88.217 66.324 88.249 66.388 ;
			RECT	88.385 66.324 88.417 66.388 ;
			RECT	88.553 66.324 88.585 66.388 ;
			RECT	88.721 66.324 88.753 66.388 ;
			RECT	88.889 66.324 88.921 66.388 ;
			RECT	89.057 66.324 89.089 66.388 ;
			RECT	89.225 66.324 89.257 66.388 ;
			RECT	89.393 66.324 89.425 66.388 ;
			RECT	89.561 66.324 89.593 66.388 ;
			RECT	89.729 66.324 89.761 66.388 ;
			RECT	89.897 66.324 89.929 66.388 ;
			RECT	90.065 66.324 90.097 66.388 ;
			RECT	90.233 66.324 90.265 66.388 ;
			RECT	90.401 66.324 90.433 66.388 ;
			RECT	90.569 66.324 90.601 66.388 ;
			RECT	90.737 66.324 90.769 66.388 ;
			RECT	90.905 66.324 90.937 66.388 ;
			RECT	91.073 66.324 91.105 66.388 ;
			RECT	91.241 66.324 91.273 66.388 ;
			RECT	91.409 66.324 91.441 66.388 ;
			RECT	91.577 66.324 91.609 66.388 ;
			RECT	91.745 66.324 91.777 66.388 ;
			RECT	91.913 66.324 91.945 66.388 ;
			RECT	92.081 66.324 92.113 66.388 ;
			RECT	92.249 66.324 92.281 66.388 ;
			RECT	92.417 66.324 92.449 66.388 ;
			RECT	92.585 66.324 92.617 66.388 ;
			RECT	92.753 66.324 92.785 66.388 ;
			RECT	92.921 66.324 92.953 66.388 ;
			RECT	93.089 66.324 93.121 66.388 ;
			RECT	93.257 66.324 93.289 66.388 ;
			RECT	93.425 66.324 93.457 66.388 ;
			RECT	93.593 66.324 93.625 66.388 ;
			RECT	93.761 66.324 93.793 66.388 ;
			RECT	93.929 66.324 93.961 66.388 ;
			RECT	94.097 66.324 94.129 66.388 ;
			RECT	94.265 66.324 94.297 66.388 ;
			RECT	94.433 66.324 94.465 66.388 ;
			RECT	94.601 66.324 94.633 66.388 ;
			RECT	94.769 66.324 94.801 66.388 ;
			RECT	94.937 66.324 94.969 66.388 ;
			RECT	95.105 66.324 95.137 66.388 ;
			RECT	95.273 66.324 95.305 66.388 ;
			RECT	95.441 66.324 95.473 66.388 ;
			RECT	95.609 66.324 95.641 66.388 ;
			RECT	95.777 66.324 95.809 66.388 ;
			RECT	95.945 66.324 95.977 66.388 ;
			RECT	96.113 66.324 96.145 66.388 ;
			RECT	96.281 66.324 96.313 66.388 ;
			RECT	96.449 66.324 96.481 66.388 ;
			RECT	96.617 66.324 96.649 66.388 ;
			RECT	96.785 66.324 96.817 66.388 ;
			RECT	96.953 66.324 96.985 66.388 ;
			RECT	97.121 66.324 97.153 66.388 ;
			RECT	97.289 66.324 97.321 66.388 ;
			RECT	97.457 66.324 97.489 66.388 ;
			RECT	97.625 66.324 97.657 66.388 ;
			RECT	97.793 66.324 97.825 66.388 ;
			RECT	97.961 66.324 97.993 66.388 ;
			RECT	98.129 66.324 98.161 66.388 ;
			RECT	98.297 66.324 98.329 66.388 ;
			RECT	98.465 66.324 98.497 66.388 ;
			RECT	98.633 66.324 98.665 66.388 ;
			RECT	98.801 66.324 98.833 66.388 ;
			RECT	98.969 66.324 99.001 66.388 ;
			RECT	99.137 66.324 99.169 66.388 ;
			RECT	99.305 66.324 99.337 66.388 ;
			RECT	99.473 66.324 99.505 66.388 ;
			RECT	99.641 66.324 99.673 66.388 ;
			RECT	99.809 66.324 99.841 66.388 ;
			RECT	99.977 66.324 100.009 66.388 ;
			RECT	100.145 66.324 100.177 66.388 ;
			RECT	100.313 66.324 100.345 66.388 ;
			RECT	100.481 66.324 100.513 66.388 ;
			RECT	100.649 66.324 100.681 66.388 ;
			RECT	100.817 66.324 100.849 66.388 ;
			RECT	100.985 66.324 101.017 66.388 ;
			RECT	101.153 66.324 101.185 66.388 ;
			RECT	101.321 66.324 101.353 66.388 ;
			RECT	101.489 66.324 101.521 66.388 ;
			RECT	101.657 66.324 101.689 66.388 ;
			RECT	101.825 66.324 101.857 66.388 ;
			RECT	101.993 66.324 102.025 66.388 ;
			RECT	102.123 66.34 102.155 66.372 ;
			RECT	102.245 66.335 102.277 66.367 ;
			RECT	102.375 66.324 102.407 66.388 ;
			RECT	103.795 66.324 103.827 66.388 ;
			RECT	103.925 66.335 103.957 66.367 ;
			RECT	104.047 66.34 104.079 66.372 ;
			RECT	104.177 66.324 104.209 66.388 ;
			RECT	104.345 66.324 104.377 66.388 ;
			RECT	104.513 66.324 104.545 66.388 ;
			RECT	104.681 66.324 104.713 66.388 ;
			RECT	104.849 66.324 104.881 66.388 ;
			RECT	105.017 66.324 105.049 66.388 ;
			RECT	105.185 66.324 105.217 66.388 ;
			RECT	105.353 66.324 105.385 66.388 ;
			RECT	105.521 66.324 105.553 66.388 ;
			RECT	105.689 66.324 105.721 66.388 ;
			RECT	105.857 66.324 105.889 66.388 ;
			RECT	106.025 66.324 106.057 66.388 ;
			RECT	106.193 66.324 106.225 66.388 ;
			RECT	106.361 66.324 106.393 66.388 ;
			RECT	106.529 66.324 106.561 66.388 ;
			RECT	106.697 66.324 106.729 66.388 ;
			RECT	106.865 66.324 106.897 66.388 ;
			RECT	107.033 66.324 107.065 66.388 ;
			RECT	107.201 66.324 107.233 66.388 ;
			RECT	107.369 66.324 107.401 66.388 ;
			RECT	107.537 66.324 107.569 66.388 ;
			RECT	107.705 66.324 107.737 66.388 ;
			RECT	107.873 66.324 107.905 66.388 ;
			RECT	108.041 66.324 108.073 66.388 ;
			RECT	108.209 66.324 108.241 66.388 ;
			RECT	108.377 66.324 108.409 66.388 ;
			RECT	108.545 66.324 108.577 66.388 ;
			RECT	108.713 66.324 108.745 66.388 ;
			RECT	108.881 66.324 108.913 66.388 ;
			RECT	109.049 66.324 109.081 66.388 ;
			RECT	109.217 66.324 109.249 66.388 ;
			RECT	109.385 66.324 109.417 66.388 ;
			RECT	109.553 66.324 109.585 66.388 ;
			RECT	109.721 66.324 109.753 66.388 ;
			RECT	109.889 66.324 109.921 66.388 ;
			RECT	110.057 66.324 110.089 66.388 ;
			RECT	110.225 66.324 110.257 66.388 ;
			RECT	110.393 66.324 110.425 66.388 ;
			RECT	110.561 66.324 110.593 66.388 ;
			RECT	110.729 66.324 110.761 66.388 ;
			RECT	110.897 66.324 110.929 66.388 ;
			RECT	111.065 66.324 111.097 66.388 ;
			RECT	111.233 66.324 111.265 66.388 ;
			RECT	111.401 66.324 111.433 66.388 ;
			RECT	111.569 66.324 111.601 66.388 ;
			RECT	111.737 66.324 111.769 66.388 ;
			RECT	111.905 66.324 111.937 66.388 ;
			RECT	112.073 66.324 112.105 66.388 ;
			RECT	112.241 66.324 112.273 66.388 ;
			RECT	112.409 66.324 112.441 66.388 ;
			RECT	112.577 66.324 112.609 66.388 ;
			RECT	112.745 66.324 112.777 66.388 ;
			RECT	112.913 66.324 112.945 66.388 ;
			RECT	113.081 66.324 113.113 66.388 ;
			RECT	113.249 66.324 113.281 66.388 ;
			RECT	113.417 66.324 113.449 66.388 ;
			RECT	113.585 66.324 113.617 66.388 ;
			RECT	113.753 66.324 113.785 66.388 ;
			RECT	113.921 66.324 113.953 66.388 ;
			RECT	114.089 66.324 114.121 66.388 ;
			RECT	114.257 66.324 114.289 66.388 ;
			RECT	114.425 66.324 114.457 66.388 ;
			RECT	114.593 66.324 114.625 66.388 ;
			RECT	114.761 66.324 114.793 66.388 ;
			RECT	114.929 66.324 114.961 66.388 ;
			RECT	115.097 66.324 115.129 66.388 ;
			RECT	115.265 66.324 115.297 66.388 ;
			RECT	115.433 66.324 115.465 66.388 ;
			RECT	115.601 66.324 115.633 66.388 ;
			RECT	115.769 66.324 115.801 66.388 ;
			RECT	115.937 66.324 115.969 66.388 ;
			RECT	116.105 66.324 116.137 66.388 ;
			RECT	116.273 66.324 116.305 66.388 ;
			RECT	116.441 66.324 116.473 66.388 ;
			RECT	116.609 66.324 116.641 66.388 ;
			RECT	116.777 66.324 116.809 66.388 ;
			RECT	116.945 66.324 116.977 66.388 ;
			RECT	117.113 66.324 117.145 66.388 ;
			RECT	117.281 66.324 117.313 66.388 ;
			RECT	117.449 66.324 117.481 66.388 ;
			RECT	117.617 66.324 117.649 66.388 ;
			RECT	117.785 66.324 117.817 66.388 ;
			RECT	117.953 66.324 117.985 66.388 ;
			RECT	118.121 66.324 118.153 66.388 ;
			RECT	118.289 66.324 118.321 66.388 ;
			RECT	118.457 66.324 118.489 66.388 ;
			RECT	118.625 66.324 118.657 66.388 ;
			RECT	118.793 66.324 118.825 66.388 ;
			RECT	118.961 66.324 118.993 66.388 ;
			RECT	119.129 66.324 119.161 66.388 ;
			RECT	119.297 66.324 119.329 66.388 ;
			RECT	119.465 66.324 119.497 66.388 ;
			RECT	119.633 66.324 119.665 66.388 ;
			RECT	119.801 66.324 119.833 66.388 ;
			RECT	119.969 66.324 120.001 66.388 ;
			RECT	120.137 66.324 120.169 66.388 ;
			RECT	120.305 66.324 120.337 66.388 ;
			RECT	120.473 66.324 120.505 66.388 ;
			RECT	120.641 66.324 120.673 66.388 ;
			RECT	120.809 66.324 120.841 66.388 ;
			RECT	120.977 66.324 121.009 66.388 ;
			RECT	121.145 66.324 121.177 66.388 ;
			RECT	121.313 66.324 121.345 66.388 ;
			RECT	121.481 66.324 121.513 66.388 ;
			RECT	121.649 66.324 121.681 66.388 ;
			RECT	121.817 66.324 121.849 66.388 ;
			RECT	121.985 66.324 122.017 66.388 ;
			RECT	122.153 66.324 122.185 66.388 ;
			RECT	122.321 66.324 122.353 66.388 ;
			RECT	122.489 66.324 122.521 66.388 ;
			RECT	122.657 66.324 122.689 66.388 ;
			RECT	122.825 66.324 122.857 66.388 ;
			RECT	122.993 66.324 123.025 66.388 ;
			RECT	123.161 66.324 123.193 66.388 ;
			RECT	123.329 66.324 123.361 66.388 ;
			RECT	123.497 66.324 123.529 66.388 ;
			RECT	123.665 66.324 123.697 66.388 ;
			RECT	123.833 66.324 123.865 66.388 ;
			RECT	124.001 66.324 124.033 66.388 ;
			RECT	124.169 66.324 124.201 66.388 ;
			RECT	124.337 66.324 124.369 66.388 ;
			RECT	124.505 66.324 124.537 66.388 ;
			RECT	124.673 66.324 124.705 66.388 ;
			RECT	124.841 66.324 124.873 66.388 ;
			RECT	125.009 66.324 125.041 66.388 ;
			RECT	125.177 66.324 125.209 66.388 ;
			RECT	125.345 66.324 125.377 66.388 ;
			RECT	125.513 66.324 125.545 66.388 ;
			RECT	125.681 66.324 125.713 66.388 ;
			RECT	125.849 66.324 125.881 66.388 ;
			RECT	126.017 66.324 126.049 66.388 ;
			RECT	126.185 66.324 126.217 66.388 ;
			RECT	126.353 66.324 126.385 66.388 ;
			RECT	126.521 66.324 126.553 66.388 ;
			RECT	126.689 66.324 126.721 66.388 ;
			RECT	126.857 66.324 126.889 66.388 ;
			RECT	127.025 66.324 127.057 66.388 ;
			RECT	127.193 66.324 127.225 66.388 ;
			RECT	127.361 66.324 127.393 66.388 ;
			RECT	127.529 66.324 127.561 66.388 ;
			RECT	127.697 66.324 127.729 66.388 ;
			RECT	127.865 66.324 127.897 66.388 ;
			RECT	128.033 66.324 128.065 66.388 ;
			RECT	128.201 66.324 128.233 66.388 ;
			RECT	128.369 66.324 128.401 66.388 ;
			RECT	128.537 66.324 128.569 66.388 ;
			RECT	128.705 66.324 128.737 66.388 ;
			RECT	128.873 66.324 128.905 66.388 ;
			RECT	129.041 66.324 129.073 66.388 ;
			RECT	129.209 66.324 129.241 66.388 ;
			RECT	129.377 66.324 129.409 66.388 ;
			RECT	129.545 66.324 129.577 66.388 ;
			RECT	129.713 66.324 129.745 66.388 ;
			RECT	129.881 66.324 129.913 66.388 ;
			RECT	130.049 66.324 130.081 66.388 ;
			RECT	130.217 66.324 130.249 66.388 ;
			RECT	130.385 66.324 130.417 66.388 ;
			RECT	130.553 66.324 130.585 66.388 ;
			RECT	130.721 66.324 130.753 66.388 ;
			RECT	130.889 66.324 130.921 66.388 ;
			RECT	131.057 66.324 131.089 66.388 ;
			RECT	131.225 66.324 131.257 66.388 ;
			RECT	131.393 66.324 131.425 66.388 ;
			RECT	131.561 66.324 131.593 66.388 ;
			RECT	131.729 66.324 131.761 66.388 ;
			RECT	131.897 66.324 131.929 66.388 ;
			RECT	132.065 66.324 132.097 66.388 ;
			RECT	132.233 66.324 132.265 66.388 ;
			RECT	132.401 66.324 132.433 66.388 ;
			RECT	132.569 66.324 132.601 66.388 ;
			RECT	132.737 66.324 132.769 66.388 ;
			RECT	132.905 66.324 132.937 66.388 ;
			RECT	133.073 66.324 133.105 66.388 ;
			RECT	133.241 66.324 133.273 66.388 ;
			RECT	133.409 66.324 133.441 66.388 ;
			RECT	133.577 66.324 133.609 66.388 ;
			RECT	133.745 66.324 133.777 66.388 ;
			RECT	133.913 66.324 133.945 66.388 ;
			RECT	134.081 66.324 134.113 66.388 ;
			RECT	134.249 66.324 134.281 66.388 ;
			RECT	134.417 66.324 134.449 66.388 ;
			RECT	134.585 66.324 134.617 66.388 ;
			RECT	134.753 66.324 134.785 66.388 ;
			RECT	134.921 66.324 134.953 66.388 ;
			RECT	135.089 66.324 135.121 66.388 ;
			RECT	135.257 66.324 135.289 66.388 ;
			RECT	135.425 66.324 135.457 66.388 ;
			RECT	135.593 66.324 135.625 66.388 ;
			RECT	135.761 66.324 135.793 66.388 ;
			RECT	135.929 66.324 135.961 66.388 ;
			RECT	136.097 66.324 136.129 66.388 ;
			RECT	136.265 66.324 136.297 66.388 ;
			RECT	136.433 66.324 136.465 66.388 ;
			RECT	136.601 66.324 136.633 66.388 ;
			RECT	136.769 66.324 136.801 66.388 ;
			RECT	136.937 66.324 136.969 66.388 ;
			RECT	137.105 66.324 137.137 66.388 ;
			RECT	137.273 66.324 137.305 66.388 ;
			RECT	137.441 66.324 137.473 66.388 ;
			RECT	137.609 66.324 137.641 66.388 ;
			RECT	137.777 66.324 137.809 66.388 ;
			RECT	137.945 66.324 137.977 66.388 ;
			RECT	138.113 66.324 138.145 66.388 ;
			RECT	138.281 66.324 138.313 66.388 ;
			RECT	138.449 66.324 138.481 66.388 ;
			RECT	138.617 66.324 138.649 66.388 ;
			RECT	138.785 66.324 138.817 66.388 ;
			RECT	138.953 66.324 138.985 66.388 ;
			RECT	139.121 66.324 139.153 66.388 ;
			RECT	139.289 66.324 139.321 66.388 ;
			RECT	139.457 66.324 139.489 66.388 ;
			RECT	139.625 66.324 139.657 66.388 ;
			RECT	139.793 66.324 139.825 66.388 ;
			RECT	139.961 66.324 139.993 66.388 ;
			RECT	140.129 66.324 140.161 66.388 ;
			RECT	140.297 66.324 140.329 66.388 ;
			RECT	140.465 66.324 140.497 66.388 ;
			RECT	140.633 66.324 140.665 66.388 ;
			RECT	140.801 66.324 140.833 66.388 ;
			RECT	140.969 66.324 141.001 66.388 ;
			RECT	141.137 66.324 141.169 66.388 ;
			RECT	141.305 66.324 141.337 66.388 ;
			RECT	141.473 66.324 141.505 66.388 ;
			RECT	141.641 66.324 141.673 66.388 ;
			RECT	141.809 66.324 141.841 66.388 ;
			RECT	141.977 66.324 142.009 66.388 ;
			RECT	142.145 66.324 142.177 66.388 ;
			RECT	142.313 66.324 142.345 66.388 ;
			RECT	142.481 66.324 142.513 66.388 ;
			RECT	142.649 66.324 142.681 66.388 ;
			RECT	142.817 66.324 142.849 66.388 ;
			RECT	142.985 66.324 143.017 66.388 ;
			RECT	143.153 66.324 143.185 66.388 ;
			RECT	143.321 66.324 143.353 66.388 ;
			RECT	143.489 66.324 143.521 66.388 ;
			RECT	143.657 66.324 143.689 66.388 ;
			RECT	143.825 66.324 143.857 66.388 ;
			RECT	143.993 66.324 144.025 66.388 ;
			RECT	144.161 66.324 144.193 66.388 ;
			RECT	144.329 66.324 144.361 66.388 ;
			RECT	144.497 66.324 144.529 66.388 ;
			RECT	144.665 66.324 144.697 66.388 ;
			RECT	144.833 66.324 144.865 66.388 ;
			RECT	145.001 66.324 145.033 66.388 ;
			RECT	145.169 66.324 145.201 66.388 ;
			RECT	145.337 66.324 145.369 66.388 ;
			RECT	145.505 66.324 145.537 66.388 ;
			RECT	145.673 66.324 145.705 66.388 ;
			RECT	145.841 66.324 145.873 66.388 ;
			RECT	146.009 66.324 146.041 66.388 ;
			RECT	146.177 66.324 146.209 66.388 ;
			RECT	146.345 66.324 146.377 66.388 ;
			RECT	146.513 66.324 146.545 66.388 ;
			RECT	146.681 66.324 146.713 66.388 ;
			RECT	146.849 66.324 146.881 66.388 ;
			RECT	147.017 66.324 147.049 66.388 ;
			RECT	147.185 66.324 147.217 66.388 ;
			RECT	147.316 66.34 147.348 66.372 ;
			RECT	147.437 66.34 147.469 66.372 ;
			RECT	147.567 66.324 147.599 66.388 ;
			RECT	149.879 66.324 149.911 66.388 ;
			RECT	151.13 66.324 151.194 66.388 ;
			RECT	151.81 66.324 151.842 66.388 ;
			RECT	152.249 66.324 152.281 66.388 ;
			RECT	153.56 66.324 153.624 66.388 ;
			RECT	156.601 66.324 156.633 66.388 ;
			RECT	156.731 66.34 156.763 66.372 ;
			RECT	156.852 66.34 156.884 66.372 ;
			RECT	156.983 66.324 157.015 66.388 ;
			RECT	157.151 66.324 157.183 66.388 ;
			RECT	157.319 66.324 157.351 66.388 ;
			RECT	157.487 66.324 157.519 66.388 ;
			RECT	157.655 66.324 157.687 66.388 ;
			RECT	157.823 66.324 157.855 66.388 ;
			RECT	157.991 66.324 158.023 66.388 ;
			RECT	158.159 66.324 158.191 66.388 ;
			RECT	158.327 66.324 158.359 66.388 ;
			RECT	158.495 66.324 158.527 66.388 ;
			RECT	158.663 66.324 158.695 66.388 ;
			RECT	158.831 66.324 158.863 66.388 ;
			RECT	158.999 66.324 159.031 66.388 ;
			RECT	159.167 66.324 159.199 66.388 ;
			RECT	159.335 66.324 159.367 66.388 ;
			RECT	159.503 66.324 159.535 66.388 ;
			RECT	159.671 66.324 159.703 66.388 ;
			RECT	159.839 66.324 159.871 66.388 ;
			RECT	160.007 66.324 160.039 66.388 ;
			RECT	160.175 66.324 160.207 66.388 ;
			RECT	160.343 66.324 160.375 66.388 ;
			RECT	160.511 66.324 160.543 66.388 ;
			RECT	160.679 66.324 160.711 66.388 ;
			RECT	160.847 66.324 160.879 66.388 ;
			RECT	161.015 66.324 161.047 66.388 ;
			RECT	161.183 66.324 161.215 66.388 ;
			RECT	161.351 66.324 161.383 66.388 ;
			RECT	161.519 66.324 161.551 66.388 ;
			RECT	161.687 66.324 161.719 66.388 ;
			RECT	161.855 66.324 161.887 66.388 ;
			RECT	162.023 66.324 162.055 66.388 ;
			RECT	162.191 66.324 162.223 66.388 ;
			RECT	162.359 66.324 162.391 66.388 ;
			RECT	162.527 66.324 162.559 66.388 ;
			RECT	162.695 66.324 162.727 66.388 ;
			RECT	162.863 66.324 162.895 66.388 ;
			RECT	163.031 66.324 163.063 66.388 ;
			RECT	163.199 66.324 163.231 66.388 ;
			RECT	163.367 66.324 163.399 66.388 ;
			RECT	163.535 66.324 163.567 66.388 ;
			RECT	163.703 66.324 163.735 66.388 ;
			RECT	163.871 66.324 163.903 66.388 ;
			RECT	164.039 66.324 164.071 66.388 ;
			RECT	164.207 66.324 164.239 66.388 ;
			RECT	164.375 66.324 164.407 66.388 ;
			RECT	164.543 66.324 164.575 66.388 ;
			RECT	164.711 66.324 164.743 66.388 ;
			RECT	164.879 66.324 164.911 66.388 ;
			RECT	165.047 66.324 165.079 66.388 ;
			RECT	165.215 66.324 165.247 66.388 ;
			RECT	165.383 66.324 165.415 66.388 ;
			RECT	165.551 66.324 165.583 66.388 ;
			RECT	165.719 66.324 165.751 66.388 ;
			RECT	165.887 66.324 165.919 66.388 ;
			RECT	166.055 66.324 166.087 66.388 ;
			RECT	166.223 66.324 166.255 66.388 ;
			RECT	166.391 66.324 166.423 66.388 ;
			RECT	166.559 66.324 166.591 66.388 ;
			RECT	166.727 66.324 166.759 66.388 ;
			RECT	166.895 66.324 166.927 66.388 ;
			RECT	167.063 66.324 167.095 66.388 ;
			RECT	167.231 66.324 167.263 66.388 ;
			RECT	167.399 66.324 167.431 66.388 ;
			RECT	167.567 66.324 167.599 66.388 ;
			RECT	167.735 66.324 167.767 66.388 ;
			RECT	167.903 66.324 167.935 66.388 ;
			RECT	168.071 66.324 168.103 66.388 ;
			RECT	168.239 66.324 168.271 66.388 ;
			RECT	168.407 66.324 168.439 66.388 ;
			RECT	168.575 66.324 168.607 66.388 ;
			RECT	168.743 66.324 168.775 66.388 ;
			RECT	168.911 66.324 168.943 66.388 ;
			RECT	169.079 66.324 169.111 66.388 ;
			RECT	169.247 66.324 169.279 66.388 ;
			RECT	169.415 66.324 169.447 66.388 ;
			RECT	169.583 66.324 169.615 66.388 ;
			RECT	169.751 66.324 169.783 66.388 ;
			RECT	169.919 66.324 169.951 66.388 ;
			RECT	170.087 66.324 170.119 66.388 ;
			RECT	170.255 66.324 170.287 66.388 ;
			RECT	170.423 66.324 170.455 66.388 ;
			RECT	170.591 66.324 170.623 66.388 ;
			RECT	170.759 66.324 170.791 66.388 ;
			RECT	170.927 66.324 170.959 66.388 ;
			RECT	171.095 66.324 171.127 66.388 ;
			RECT	171.263 66.324 171.295 66.388 ;
			RECT	171.431 66.324 171.463 66.388 ;
			RECT	171.599 66.324 171.631 66.388 ;
			RECT	171.767 66.324 171.799 66.388 ;
			RECT	171.935 66.324 171.967 66.388 ;
			RECT	172.103 66.324 172.135 66.388 ;
			RECT	172.271 66.324 172.303 66.388 ;
			RECT	172.439 66.324 172.471 66.388 ;
			RECT	172.607 66.324 172.639 66.388 ;
			RECT	172.775 66.324 172.807 66.388 ;
			RECT	172.943 66.324 172.975 66.388 ;
			RECT	173.111 66.324 173.143 66.388 ;
			RECT	173.279 66.324 173.311 66.388 ;
			RECT	173.447 66.324 173.479 66.388 ;
			RECT	173.615 66.324 173.647 66.388 ;
			RECT	173.783 66.324 173.815 66.388 ;
			RECT	173.951 66.324 173.983 66.388 ;
			RECT	174.119 66.324 174.151 66.388 ;
			RECT	174.287 66.324 174.319 66.388 ;
			RECT	174.455 66.324 174.487 66.388 ;
			RECT	174.623 66.324 174.655 66.388 ;
			RECT	174.791 66.324 174.823 66.388 ;
			RECT	174.959 66.324 174.991 66.388 ;
			RECT	175.127 66.324 175.159 66.388 ;
			RECT	175.295 66.324 175.327 66.388 ;
			RECT	175.463 66.324 175.495 66.388 ;
			RECT	175.631 66.324 175.663 66.388 ;
			RECT	175.799 66.324 175.831 66.388 ;
			RECT	175.967 66.324 175.999 66.388 ;
			RECT	176.135 66.324 176.167 66.388 ;
			RECT	176.303 66.324 176.335 66.388 ;
			RECT	176.471 66.324 176.503 66.388 ;
			RECT	176.639 66.324 176.671 66.388 ;
			RECT	176.807 66.324 176.839 66.388 ;
			RECT	176.975 66.324 177.007 66.388 ;
			RECT	177.143 66.324 177.175 66.388 ;
			RECT	177.311 66.324 177.343 66.388 ;
			RECT	177.479 66.324 177.511 66.388 ;
			RECT	177.647 66.324 177.679 66.388 ;
			RECT	177.815 66.324 177.847 66.388 ;
			RECT	177.983 66.324 178.015 66.388 ;
			RECT	178.151 66.324 178.183 66.388 ;
			RECT	178.319 66.324 178.351 66.388 ;
			RECT	178.487 66.324 178.519 66.388 ;
			RECT	178.655 66.324 178.687 66.388 ;
			RECT	178.823 66.324 178.855 66.388 ;
			RECT	178.991 66.324 179.023 66.388 ;
			RECT	179.159 66.324 179.191 66.388 ;
			RECT	179.327 66.324 179.359 66.388 ;
			RECT	179.495 66.324 179.527 66.388 ;
			RECT	179.663 66.324 179.695 66.388 ;
			RECT	179.831 66.324 179.863 66.388 ;
			RECT	179.999 66.324 180.031 66.388 ;
			RECT	180.167 66.324 180.199 66.388 ;
			RECT	180.335 66.324 180.367 66.388 ;
			RECT	180.503 66.324 180.535 66.388 ;
			RECT	180.671 66.324 180.703 66.388 ;
			RECT	180.839 66.324 180.871 66.388 ;
			RECT	181.007 66.324 181.039 66.388 ;
			RECT	181.175 66.324 181.207 66.388 ;
			RECT	181.343 66.324 181.375 66.388 ;
			RECT	181.511 66.324 181.543 66.388 ;
			RECT	181.679 66.324 181.711 66.388 ;
			RECT	181.847 66.324 181.879 66.388 ;
			RECT	182.015 66.324 182.047 66.388 ;
			RECT	182.183 66.324 182.215 66.388 ;
			RECT	182.351 66.324 182.383 66.388 ;
			RECT	182.519 66.324 182.551 66.388 ;
			RECT	182.687 66.324 182.719 66.388 ;
			RECT	182.855 66.324 182.887 66.388 ;
			RECT	183.023 66.324 183.055 66.388 ;
			RECT	183.191 66.324 183.223 66.388 ;
			RECT	183.359 66.324 183.391 66.388 ;
			RECT	183.527 66.324 183.559 66.388 ;
			RECT	183.695 66.324 183.727 66.388 ;
			RECT	183.863 66.324 183.895 66.388 ;
			RECT	184.031 66.324 184.063 66.388 ;
			RECT	184.199 66.324 184.231 66.388 ;
			RECT	184.367 66.324 184.399 66.388 ;
			RECT	184.535 66.324 184.567 66.388 ;
			RECT	184.703 66.324 184.735 66.388 ;
			RECT	184.871 66.324 184.903 66.388 ;
			RECT	185.039 66.324 185.071 66.388 ;
			RECT	185.207 66.324 185.239 66.388 ;
			RECT	185.375 66.324 185.407 66.388 ;
			RECT	185.543 66.324 185.575 66.388 ;
			RECT	185.711 66.324 185.743 66.388 ;
			RECT	185.879 66.324 185.911 66.388 ;
			RECT	186.047 66.324 186.079 66.388 ;
			RECT	186.215 66.324 186.247 66.388 ;
			RECT	186.383 66.324 186.415 66.388 ;
			RECT	186.551 66.324 186.583 66.388 ;
			RECT	186.719 66.324 186.751 66.388 ;
			RECT	186.887 66.324 186.919 66.388 ;
			RECT	187.055 66.324 187.087 66.388 ;
			RECT	187.223 66.324 187.255 66.388 ;
			RECT	187.391 66.324 187.423 66.388 ;
			RECT	187.559 66.324 187.591 66.388 ;
			RECT	187.727 66.324 187.759 66.388 ;
			RECT	187.895 66.324 187.927 66.388 ;
			RECT	188.063 66.324 188.095 66.388 ;
			RECT	188.231 66.324 188.263 66.388 ;
			RECT	188.399 66.324 188.431 66.388 ;
			RECT	188.567 66.324 188.599 66.388 ;
			RECT	188.735 66.324 188.767 66.388 ;
			RECT	188.903 66.324 188.935 66.388 ;
			RECT	189.071 66.324 189.103 66.388 ;
			RECT	189.239 66.324 189.271 66.388 ;
			RECT	189.407 66.324 189.439 66.388 ;
			RECT	189.575 66.324 189.607 66.388 ;
			RECT	189.743 66.324 189.775 66.388 ;
			RECT	189.911 66.324 189.943 66.388 ;
			RECT	190.079 66.324 190.111 66.388 ;
			RECT	190.247 66.324 190.279 66.388 ;
			RECT	190.415 66.324 190.447 66.388 ;
			RECT	190.583 66.324 190.615 66.388 ;
			RECT	190.751 66.324 190.783 66.388 ;
			RECT	190.919 66.324 190.951 66.388 ;
			RECT	191.087 66.324 191.119 66.388 ;
			RECT	191.255 66.324 191.287 66.388 ;
			RECT	191.423 66.324 191.455 66.388 ;
			RECT	191.591 66.324 191.623 66.388 ;
			RECT	191.759 66.324 191.791 66.388 ;
			RECT	191.927 66.324 191.959 66.388 ;
			RECT	192.095 66.324 192.127 66.388 ;
			RECT	192.263 66.324 192.295 66.388 ;
			RECT	192.431 66.324 192.463 66.388 ;
			RECT	192.599 66.324 192.631 66.388 ;
			RECT	192.767 66.324 192.799 66.388 ;
			RECT	192.935 66.324 192.967 66.388 ;
			RECT	193.103 66.324 193.135 66.388 ;
			RECT	193.271 66.324 193.303 66.388 ;
			RECT	193.439 66.324 193.471 66.388 ;
			RECT	193.607 66.324 193.639 66.388 ;
			RECT	193.775 66.324 193.807 66.388 ;
			RECT	193.943 66.324 193.975 66.388 ;
			RECT	194.111 66.324 194.143 66.388 ;
			RECT	194.279 66.324 194.311 66.388 ;
			RECT	194.447 66.324 194.479 66.388 ;
			RECT	194.615 66.324 194.647 66.388 ;
			RECT	194.783 66.324 194.815 66.388 ;
			RECT	194.951 66.324 194.983 66.388 ;
			RECT	195.119 66.324 195.151 66.388 ;
			RECT	195.287 66.324 195.319 66.388 ;
			RECT	195.455 66.324 195.487 66.388 ;
			RECT	195.623 66.324 195.655 66.388 ;
			RECT	195.791 66.324 195.823 66.388 ;
			RECT	195.959 66.324 195.991 66.388 ;
			RECT	196.127 66.324 196.159 66.388 ;
			RECT	196.295 66.324 196.327 66.388 ;
			RECT	196.463 66.324 196.495 66.388 ;
			RECT	196.631 66.324 196.663 66.388 ;
			RECT	196.799 66.324 196.831 66.388 ;
			RECT	196.967 66.324 196.999 66.388 ;
			RECT	197.135 66.324 197.167 66.388 ;
			RECT	197.303 66.324 197.335 66.388 ;
			RECT	197.471 66.324 197.503 66.388 ;
			RECT	197.639 66.324 197.671 66.388 ;
			RECT	197.807 66.324 197.839 66.388 ;
			RECT	197.975 66.324 198.007 66.388 ;
			RECT	198.143 66.324 198.175 66.388 ;
			RECT	198.311 66.324 198.343 66.388 ;
			RECT	198.479 66.324 198.511 66.388 ;
			RECT	198.647 66.324 198.679 66.388 ;
			RECT	198.815 66.324 198.847 66.388 ;
			RECT	198.983 66.324 199.015 66.388 ;
			RECT	199.151 66.324 199.183 66.388 ;
			RECT	199.319 66.324 199.351 66.388 ;
			RECT	199.487 66.324 199.519 66.388 ;
			RECT	199.655 66.324 199.687 66.388 ;
			RECT	199.823 66.324 199.855 66.388 ;
			RECT	199.991 66.324 200.023 66.388 ;
			RECT	200.121 66.34 200.153 66.372 ;
			RECT	200.243 66.335 200.275 66.367 ;
			RECT	200.373 66.324 200.405 66.388 ;
			RECT	200.9 66.324 200.932 66.388 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 64.376 201.665 64.496 ;
			LAYER	J3 ;
			RECT	0.755 64.404 0.787 64.468 ;
			RECT	1.645 64.404 1.709 64.468 ;
			RECT	2.323 64.404 2.387 64.468 ;
			RECT	3.438 64.404 3.47 64.468 ;
			RECT	3.585 64.404 3.617 64.468 ;
			RECT	4.195 64.404 4.227 64.468 ;
			RECT	4.72 64.404 4.752 64.468 ;
			RECT	4.944 64.404 5.008 64.468 ;
			RECT	5.267 64.404 5.299 64.468 ;
			RECT	5.797 64.404 5.829 64.468 ;
			RECT	5.927 64.415 5.959 64.447 ;
			RECT	6.049 64.42 6.081 64.452 ;
			RECT	6.179 64.404 6.211 64.468 ;
			RECT	6.347 64.404 6.379 64.468 ;
			RECT	6.515 64.404 6.547 64.468 ;
			RECT	6.683 64.404 6.715 64.468 ;
			RECT	6.851 64.404 6.883 64.468 ;
			RECT	7.019 64.404 7.051 64.468 ;
			RECT	7.187 64.404 7.219 64.468 ;
			RECT	7.355 64.404 7.387 64.468 ;
			RECT	7.523 64.404 7.555 64.468 ;
			RECT	7.691 64.404 7.723 64.468 ;
			RECT	7.859 64.404 7.891 64.468 ;
			RECT	8.027 64.404 8.059 64.468 ;
			RECT	8.195 64.404 8.227 64.468 ;
			RECT	8.363 64.404 8.395 64.468 ;
			RECT	8.531 64.404 8.563 64.468 ;
			RECT	8.699 64.404 8.731 64.468 ;
			RECT	8.867 64.404 8.899 64.468 ;
			RECT	9.035 64.404 9.067 64.468 ;
			RECT	9.203 64.404 9.235 64.468 ;
			RECT	9.371 64.404 9.403 64.468 ;
			RECT	9.539 64.404 9.571 64.468 ;
			RECT	9.707 64.404 9.739 64.468 ;
			RECT	9.875 64.404 9.907 64.468 ;
			RECT	10.043 64.404 10.075 64.468 ;
			RECT	10.211 64.404 10.243 64.468 ;
			RECT	10.379 64.404 10.411 64.468 ;
			RECT	10.547 64.404 10.579 64.468 ;
			RECT	10.715 64.404 10.747 64.468 ;
			RECT	10.883 64.404 10.915 64.468 ;
			RECT	11.051 64.404 11.083 64.468 ;
			RECT	11.219 64.404 11.251 64.468 ;
			RECT	11.387 64.404 11.419 64.468 ;
			RECT	11.555 64.404 11.587 64.468 ;
			RECT	11.723 64.404 11.755 64.468 ;
			RECT	11.891 64.404 11.923 64.468 ;
			RECT	12.059 64.404 12.091 64.468 ;
			RECT	12.227 64.404 12.259 64.468 ;
			RECT	12.395 64.404 12.427 64.468 ;
			RECT	12.563 64.404 12.595 64.468 ;
			RECT	12.731 64.404 12.763 64.468 ;
			RECT	12.899 64.404 12.931 64.468 ;
			RECT	13.067 64.404 13.099 64.468 ;
			RECT	13.235 64.404 13.267 64.468 ;
			RECT	13.403 64.404 13.435 64.468 ;
			RECT	13.571 64.404 13.603 64.468 ;
			RECT	13.739 64.404 13.771 64.468 ;
			RECT	13.907 64.404 13.939 64.468 ;
			RECT	14.075 64.404 14.107 64.468 ;
			RECT	14.243 64.404 14.275 64.468 ;
			RECT	14.411 64.404 14.443 64.468 ;
			RECT	14.579 64.404 14.611 64.468 ;
			RECT	14.747 64.404 14.779 64.468 ;
			RECT	14.915 64.404 14.947 64.468 ;
			RECT	15.083 64.404 15.115 64.468 ;
			RECT	15.251 64.404 15.283 64.468 ;
			RECT	15.419 64.404 15.451 64.468 ;
			RECT	15.587 64.404 15.619 64.468 ;
			RECT	15.755 64.404 15.787 64.468 ;
			RECT	15.923 64.404 15.955 64.468 ;
			RECT	16.091 64.404 16.123 64.468 ;
			RECT	16.259 64.404 16.291 64.468 ;
			RECT	16.427 64.404 16.459 64.468 ;
			RECT	16.595 64.404 16.627 64.468 ;
			RECT	16.763 64.404 16.795 64.468 ;
			RECT	16.931 64.404 16.963 64.468 ;
			RECT	17.099 64.404 17.131 64.468 ;
			RECT	17.267 64.404 17.299 64.468 ;
			RECT	17.435 64.404 17.467 64.468 ;
			RECT	17.603 64.404 17.635 64.468 ;
			RECT	17.771 64.404 17.803 64.468 ;
			RECT	17.939 64.404 17.971 64.468 ;
			RECT	18.107 64.404 18.139 64.468 ;
			RECT	18.275 64.404 18.307 64.468 ;
			RECT	18.443 64.404 18.475 64.468 ;
			RECT	18.611 64.404 18.643 64.468 ;
			RECT	18.779 64.404 18.811 64.468 ;
			RECT	18.947 64.404 18.979 64.468 ;
			RECT	19.115 64.404 19.147 64.468 ;
			RECT	19.283 64.404 19.315 64.468 ;
			RECT	19.451 64.404 19.483 64.468 ;
			RECT	19.619 64.404 19.651 64.468 ;
			RECT	19.787 64.404 19.819 64.468 ;
			RECT	19.955 64.404 19.987 64.468 ;
			RECT	20.123 64.404 20.155 64.468 ;
			RECT	20.291 64.404 20.323 64.468 ;
			RECT	20.459 64.404 20.491 64.468 ;
			RECT	20.627 64.404 20.659 64.468 ;
			RECT	20.795 64.404 20.827 64.468 ;
			RECT	20.963 64.404 20.995 64.468 ;
			RECT	21.131 64.404 21.163 64.468 ;
			RECT	21.299 64.404 21.331 64.468 ;
			RECT	21.467 64.404 21.499 64.468 ;
			RECT	21.635 64.404 21.667 64.468 ;
			RECT	21.803 64.404 21.835 64.468 ;
			RECT	21.971 64.404 22.003 64.468 ;
			RECT	22.139 64.404 22.171 64.468 ;
			RECT	22.307 64.404 22.339 64.468 ;
			RECT	22.475 64.404 22.507 64.468 ;
			RECT	22.643 64.404 22.675 64.468 ;
			RECT	22.811 64.404 22.843 64.468 ;
			RECT	22.979 64.404 23.011 64.468 ;
			RECT	23.147 64.404 23.179 64.468 ;
			RECT	23.315 64.404 23.347 64.468 ;
			RECT	23.483 64.404 23.515 64.468 ;
			RECT	23.651 64.404 23.683 64.468 ;
			RECT	23.819 64.404 23.851 64.468 ;
			RECT	23.987 64.404 24.019 64.468 ;
			RECT	24.155 64.404 24.187 64.468 ;
			RECT	24.323 64.404 24.355 64.468 ;
			RECT	24.491 64.404 24.523 64.468 ;
			RECT	24.659 64.404 24.691 64.468 ;
			RECT	24.827 64.404 24.859 64.468 ;
			RECT	24.995 64.404 25.027 64.468 ;
			RECT	25.163 64.404 25.195 64.468 ;
			RECT	25.331 64.404 25.363 64.468 ;
			RECT	25.499 64.404 25.531 64.468 ;
			RECT	25.667 64.404 25.699 64.468 ;
			RECT	25.835 64.404 25.867 64.468 ;
			RECT	26.003 64.404 26.035 64.468 ;
			RECT	26.171 64.404 26.203 64.468 ;
			RECT	26.339 64.404 26.371 64.468 ;
			RECT	26.507 64.404 26.539 64.468 ;
			RECT	26.675 64.404 26.707 64.468 ;
			RECT	26.843 64.404 26.875 64.468 ;
			RECT	27.011 64.404 27.043 64.468 ;
			RECT	27.179 64.404 27.211 64.468 ;
			RECT	27.347 64.404 27.379 64.468 ;
			RECT	27.515 64.404 27.547 64.468 ;
			RECT	27.683 64.404 27.715 64.468 ;
			RECT	27.851 64.404 27.883 64.468 ;
			RECT	28.019 64.404 28.051 64.468 ;
			RECT	28.187 64.404 28.219 64.468 ;
			RECT	28.355 64.404 28.387 64.468 ;
			RECT	28.523 64.404 28.555 64.468 ;
			RECT	28.691 64.404 28.723 64.468 ;
			RECT	28.859 64.404 28.891 64.468 ;
			RECT	29.027 64.404 29.059 64.468 ;
			RECT	29.195 64.404 29.227 64.468 ;
			RECT	29.363 64.404 29.395 64.468 ;
			RECT	29.531 64.404 29.563 64.468 ;
			RECT	29.699 64.404 29.731 64.468 ;
			RECT	29.867 64.404 29.899 64.468 ;
			RECT	30.035 64.404 30.067 64.468 ;
			RECT	30.203 64.404 30.235 64.468 ;
			RECT	30.371 64.404 30.403 64.468 ;
			RECT	30.539 64.404 30.571 64.468 ;
			RECT	30.707 64.404 30.739 64.468 ;
			RECT	30.875 64.404 30.907 64.468 ;
			RECT	31.043 64.404 31.075 64.468 ;
			RECT	31.211 64.404 31.243 64.468 ;
			RECT	31.379 64.404 31.411 64.468 ;
			RECT	31.547 64.404 31.579 64.468 ;
			RECT	31.715 64.404 31.747 64.468 ;
			RECT	31.883 64.404 31.915 64.468 ;
			RECT	32.051 64.404 32.083 64.468 ;
			RECT	32.219 64.404 32.251 64.468 ;
			RECT	32.387 64.404 32.419 64.468 ;
			RECT	32.555 64.404 32.587 64.468 ;
			RECT	32.723 64.404 32.755 64.468 ;
			RECT	32.891 64.404 32.923 64.468 ;
			RECT	33.059 64.404 33.091 64.468 ;
			RECT	33.227 64.404 33.259 64.468 ;
			RECT	33.395 64.404 33.427 64.468 ;
			RECT	33.563 64.404 33.595 64.468 ;
			RECT	33.731 64.404 33.763 64.468 ;
			RECT	33.899 64.404 33.931 64.468 ;
			RECT	34.067 64.404 34.099 64.468 ;
			RECT	34.235 64.404 34.267 64.468 ;
			RECT	34.403 64.404 34.435 64.468 ;
			RECT	34.571 64.404 34.603 64.468 ;
			RECT	34.739 64.404 34.771 64.468 ;
			RECT	34.907 64.404 34.939 64.468 ;
			RECT	35.075 64.404 35.107 64.468 ;
			RECT	35.243 64.404 35.275 64.468 ;
			RECT	35.411 64.404 35.443 64.468 ;
			RECT	35.579 64.404 35.611 64.468 ;
			RECT	35.747 64.404 35.779 64.468 ;
			RECT	35.915 64.404 35.947 64.468 ;
			RECT	36.083 64.404 36.115 64.468 ;
			RECT	36.251 64.404 36.283 64.468 ;
			RECT	36.419 64.404 36.451 64.468 ;
			RECT	36.587 64.404 36.619 64.468 ;
			RECT	36.755 64.404 36.787 64.468 ;
			RECT	36.923 64.404 36.955 64.468 ;
			RECT	37.091 64.404 37.123 64.468 ;
			RECT	37.259 64.404 37.291 64.468 ;
			RECT	37.427 64.404 37.459 64.468 ;
			RECT	37.595 64.404 37.627 64.468 ;
			RECT	37.763 64.404 37.795 64.468 ;
			RECT	37.931 64.404 37.963 64.468 ;
			RECT	38.099 64.404 38.131 64.468 ;
			RECT	38.267 64.404 38.299 64.468 ;
			RECT	38.435 64.404 38.467 64.468 ;
			RECT	38.603 64.404 38.635 64.468 ;
			RECT	38.771 64.404 38.803 64.468 ;
			RECT	38.939 64.404 38.971 64.468 ;
			RECT	39.107 64.404 39.139 64.468 ;
			RECT	39.275 64.404 39.307 64.468 ;
			RECT	39.443 64.404 39.475 64.468 ;
			RECT	39.611 64.404 39.643 64.468 ;
			RECT	39.779 64.404 39.811 64.468 ;
			RECT	39.947 64.404 39.979 64.468 ;
			RECT	40.115 64.404 40.147 64.468 ;
			RECT	40.283 64.404 40.315 64.468 ;
			RECT	40.451 64.404 40.483 64.468 ;
			RECT	40.619 64.404 40.651 64.468 ;
			RECT	40.787 64.404 40.819 64.468 ;
			RECT	40.955 64.404 40.987 64.468 ;
			RECT	41.123 64.404 41.155 64.468 ;
			RECT	41.291 64.404 41.323 64.468 ;
			RECT	41.459 64.404 41.491 64.468 ;
			RECT	41.627 64.404 41.659 64.468 ;
			RECT	41.795 64.404 41.827 64.468 ;
			RECT	41.963 64.404 41.995 64.468 ;
			RECT	42.131 64.404 42.163 64.468 ;
			RECT	42.299 64.404 42.331 64.468 ;
			RECT	42.467 64.404 42.499 64.468 ;
			RECT	42.635 64.404 42.667 64.468 ;
			RECT	42.803 64.404 42.835 64.468 ;
			RECT	42.971 64.404 43.003 64.468 ;
			RECT	43.139 64.404 43.171 64.468 ;
			RECT	43.307 64.404 43.339 64.468 ;
			RECT	43.475 64.404 43.507 64.468 ;
			RECT	43.643 64.404 43.675 64.468 ;
			RECT	43.811 64.404 43.843 64.468 ;
			RECT	43.979 64.404 44.011 64.468 ;
			RECT	44.147 64.404 44.179 64.468 ;
			RECT	44.315 64.404 44.347 64.468 ;
			RECT	44.483 64.404 44.515 64.468 ;
			RECT	44.651 64.404 44.683 64.468 ;
			RECT	44.819 64.404 44.851 64.468 ;
			RECT	44.987 64.404 45.019 64.468 ;
			RECT	45.155 64.404 45.187 64.468 ;
			RECT	45.323 64.404 45.355 64.468 ;
			RECT	45.491 64.404 45.523 64.468 ;
			RECT	45.659 64.404 45.691 64.468 ;
			RECT	45.827 64.404 45.859 64.468 ;
			RECT	45.995 64.404 46.027 64.468 ;
			RECT	46.163 64.404 46.195 64.468 ;
			RECT	46.331 64.404 46.363 64.468 ;
			RECT	46.499 64.404 46.531 64.468 ;
			RECT	46.667 64.404 46.699 64.468 ;
			RECT	46.835 64.404 46.867 64.468 ;
			RECT	47.003 64.404 47.035 64.468 ;
			RECT	47.171 64.404 47.203 64.468 ;
			RECT	47.339 64.404 47.371 64.468 ;
			RECT	47.507 64.404 47.539 64.468 ;
			RECT	47.675 64.404 47.707 64.468 ;
			RECT	47.843 64.404 47.875 64.468 ;
			RECT	48.011 64.404 48.043 64.468 ;
			RECT	48.179 64.404 48.211 64.468 ;
			RECT	48.347 64.404 48.379 64.468 ;
			RECT	48.515 64.404 48.547 64.468 ;
			RECT	48.683 64.404 48.715 64.468 ;
			RECT	48.851 64.404 48.883 64.468 ;
			RECT	49.019 64.404 49.051 64.468 ;
			RECT	49.187 64.404 49.219 64.468 ;
			RECT	49.318 64.42 49.35 64.452 ;
			RECT	49.439 64.42 49.471 64.452 ;
			RECT	49.569 64.404 49.601 64.468 ;
			RECT	51.881 64.404 51.913 64.468 ;
			RECT	53.132 64.404 53.196 64.468 ;
			RECT	53.812 64.404 53.844 64.468 ;
			RECT	54.251 64.404 54.283 64.468 ;
			RECT	55.562 64.404 55.626 64.468 ;
			RECT	58.603 64.404 58.635 64.468 ;
			RECT	58.733 64.42 58.765 64.452 ;
			RECT	58.854 64.42 58.886 64.452 ;
			RECT	58.985 64.404 59.017 64.468 ;
			RECT	59.153 64.404 59.185 64.468 ;
			RECT	59.321 64.404 59.353 64.468 ;
			RECT	59.489 64.404 59.521 64.468 ;
			RECT	59.657 64.404 59.689 64.468 ;
			RECT	59.825 64.404 59.857 64.468 ;
			RECT	59.993 64.404 60.025 64.468 ;
			RECT	60.161 64.404 60.193 64.468 ;
			RECT	60.329 64.404 60.361 64.468 ;
			RECT	60.497 64.404 60.529 64.468 ;
			RECT	60.665 64.404 60.697 64.468 ;
			RECT	60.833 64.404 60.865 64.468 ;
			RECT	61.001 64.404 61.033 64.468 ;
			RECT	61.169 64.404 61.201 64.468 ;
			RECT	61.337 64.404 61.369 64.468 ;
			RECT	61.505 64.404 61.537 64.468 ;
			RECT	61.673 64.404 61.705 64.468 ;
			RECT	61.841 64.404 61.873 64.468 ;
			RECT	62.009 64.404 62.041 64.468 ;
			RECT	62.177 64.404 62.209 64.468 ;
			RECT	62.345 64.404 62.377 64.468 ;
			RECT	62.513 64.404 62.545 64.468 ;
			RECT	62.681 64.404 62.713 64.468 ;
			RECT	62.849 64.404 62.881 64.468 ;
			RECT	63.017 64.404 63.049 64.468 ;
			RECT	63.185 64.404 63.217 64.468 ;
			RECT	63.353 64.404 63.385 64.468 ;
			RECT	63.521 64.404 63.553 64.468 ;
			RECT	63.689 64.404 63.721 64.468 ;
			RECT	63.857 64.404 63.889 64.468 ;
			RECT	64.025 64.404 64.057 64.468 ;
			RECT	64.193 64.404 64.225 64.468 ;
			RECT	64.361 64.404 64.393 64.468 ;
			RECT	64.529 64.404 64.561 64.468 ;
			RECT	64.697 64.404 64.729 64.468 ;
			RECT	64.865 64.404 64.897 64.468 ;
			RECT	65.033 64.404 65.065 64.468 ;
			RECT	65.201 64.404 65.233 64.468 ;
			RECT	65.369 64.404 65.401 64.468 ;
			RECT	65.537 64.404 65.569 64.468 ;
			RECT	65.705 64.404 65.737 64.468 ;
			RECT	65.873 64.404 65.905 64.468 ;
			RECT	66.041 64.404 66.073 64.468 ;
			RECT	66.209 64.404 66.241 64.468 ;
			RECT	66.377 64.404 66.409 64.468 ;
			RECT	66.545 64.404 66.577 64.468 ;
			RECT	66.713 64.404 66.745 64.468 ;
			RECT	66.881 64.404 66.913 64.468 ;
			RECT	67.049 64.404 67.081 64.468 ;
			RECT	67.217 64.404 67.249 64.468 ;
			RECT	67.385 64.404 67.417 64.468 ;
			RECT	67.553 64.404 67.585 64.468 ;
			RECT	67.721 64.404 67.753 64.468 ;
			RECT	67.889 64.404 67.921 64.468 ;
			RECT	68.057 64.404 68.089 64.468 ;
			RECT	68.225 64.404 68.257 64.468 ;
			RECT	68.393 64.404 68.425 64.468 ;
			RECT	68.561 64.404 68.593 64.468 ;
			RECT	68.729 64.404 68.761 64.468 ;
			RECT	68.897 64.404 68.929 64.468 ;
			RECT	69.065 64.404 69.097 64.468 ;
			RECT	69.233 64.404 69.265 64.468 ;
			RECT	69.401 64.404 69.433 64.468 ;
			RECT	69.569 64.404 69.601 64.468 ;
			RECT	69.737 64.404 69.769 64.468 ;
			RECT	69.905 64.404 69.937 64.468 ;
			RECT	70.073 64.404 70.105 64.468 ;
			RECT	70.241 64.404 70.273 64.468 ;
			RECT	70.409 64.404 70.441 64.468 ;
			RECT	70.577 64.404 70.609 64.468 ;
			RECT	70.745 64.404 70.777 64.468 ;
			RECT	70.913 64.404 70.945 64.468 ;
			RECT	71.081 64.404 71.113 64.468 ;
			RECT	71.249 64.404 71.281 64.468 ;
			RECT	71.417 64.404 71.449 64.468 ;
			RECT	71.585 64.404 71.617 64.468 ;
			RECT	71.753 64.404 71.785 64.468 ;
			RECT	71.921 64.404 71.953 64.468 ;
			RECT	72.089 64.404 72.121 64.468 ;
			RECT	72.257 64.404 72.289 64.468 ;
			RECT	72.425 64.404 72.457 64.468 ;
			RECT	72.593 64.404 72.625 64.468 ;
			RECT	72.761 64.404 72.793 64.468 ;
			RECT	72.929 64.404 72.961 64.468 ;
			RECT	73.097 64.404 73.129 64.468 ;
			RECT	73.265 64.404 73.297 64.468 ;
			RECT	73.433 64.404 73.465 64.468 ;
			RECT	73.601 64.404 73.633 64.468 ;
			RECT	73.769 64.404 73.801 64.468 ;
			RECT	73.937 64.404 73.969 64.468 ;
			RECT	74.105 64.404 74.137 64.468 ;
			RECT	74.273 64.404 74.305 64.468 ;
			RECT	74.441 64.404 74.473 64.468 ;
			RECT	74.609 64.404 74.641 64.468 ;
			RECT	74.777 64.404 74.809 64.468 ;
			RECT	74.945 64.404 74.977 64.468 ;
			RECT	75.113 64.404 75.145 64.468 ;
			RECT	75.281 64.404 75.313 64.468 ;
			RECT	75.449 64.404 75.481 64.468 ;
			RECT	75.617 64.404 75.649 64.468 ;
			RECT	75.785 64.404 75.817 64.468 ;
			RECT	75.953 64.404 75.985 64.468 ;
			RECT	76.121 64.404 76.153 64.468 ;
			RECT	76.289 64.404 76.321 64.468 ;
			RECT	76.457 64.404 76.489 64.468 ;
			RECT	76.625 64.404 76.657 64.468 ;
			RECT	76.793 64.404 76.825 64.468 ;
			RECT	76.961 64.404 76.993 64.468 ;
			RECT	77.129 64.404 77.161 64.468 ;
			RECT	77.297 64.404 77.329 64.468 ;
			RECT	77.465 64.404 77.497 64.468 ;
			RECT	77.633 64.404 77.665 64.468 ;
			RECT	77.801 64.404 77.833 64.468 ;
			RECT	77.969 64.404 78.001 64.468 ;
			RECT	78.137 64.404 78.169 64.468 ;
			RECT	78.305 64.404 78.337 64.468 ;
			RECT	78.473 64.404 78.505 64.468 ;
			RECT	78.641 64.404 78.673 64.468 ;
			RECT	78.809 64.404 78.841 64.468 ;
			RECT	78.977 64.404 79.009 64.468 ;
			RECT	79.145 64.404 79.177 64.468 ;
			RECT	79.313 64.404 79.345 64.468 ;
			RECT	79.481 64.404 79.513 64.468 ;
			RECT	79.649 64.404 79.681 64.468 ;
			RECT	79.817 64.404 79.849 64.468 ;
			RECT	79.985 64.404 80.017 64.468 ;
			RECT	80.153 64.404 80.185 64.468 ;
			RECT	80.321 64.404 80.353 64.468 ;
			RECT	80.489 64.404 80.521 64.468 ;
			RECT	80.657 64.404 80.689 64.468 ;
			RECT	80.825 64.404 80.857 64.468 ;
			RECT	80.993 64.404 81.025 64.468 ;
			RECT	81.161 64.404 81.193 64.468 ;
			RECT	81.329 64.404 81.361 64.468 ;
			RECT	81.497 64.404 81.529 64.468 ;
			RECT	81.665 64.404 81.697 64.468 ;
			RECT	81.833 64.404 81.865 64.468 ;
			RECT	82.001 64.404 82.033 64.468 ;
			RECT	82.169 64.404 82.201 64.468 ;
			RECT	82.337 64.404 82.369 64.468 ;
			RECT	82.505 64.404 82.537 64.468 ;
			RECT	82.673 64.404 82.705 64.468 ;
			RECT	82.841 64.404 82.873 64.468 ;
			RECT	83.009 64.404 83.041 64.468 ;
			RECT	83.177 64.404 83.209 64.468 ;
			RECT	83.345 64.404 83.377 64.468 ;
			RECT	83.513 64.404 83.545 64.468 ;
			RECT	83.681 64.404 83.713 64.468 ;
			RECT	83.849 64.404 83.881 64.468 ;
			RECT	84.017 64.404 84.049 64.468 ;
			RECT	84.185 64.404 84.217 64.468 ;
			RECT	84.353 64.404 84.385 64.468 ;
			RECT	84.521 64.404 84.553 64.468 ;
			RECT	84.689 64.404 84.721 64.468 ;
			RECT	84.857 64.404 84.889 64.468 ;
			RECT	85.025 64.404 85.057 64.468 ;
			RECT	85.193 64.404 85.225 64.468 ;
			RECT	85.361 64.404 85.393 64.468 ;
			RECT	85.529 64.404 85.561 64.468 ;
			RECT	85.697 64.404 85.729 64.468 ;
			RECT	85.865 64.404 85.897 64.468 ;
			RECT	86.033 64.404 86.065 64.468 ;
			RECT	86.201 64.404 86.233 64.468 ;
			RECT	86.369 64.404 86.401 64.468 ;
			RECT	86.537 64.404 86.569 64.468 ;
			RECT	86.705 64.404 86.737 64.468 ;
			RECT	86.873 64.404 86.905 64.468 ;
			RECT	87.041 64.404 87.073 64.468 ;
			RECT	87.209 64.404 87.241 64.468 ;
			RECT	87.377 64.404 87.409 64.468 ;
			RECT	87.545 64.404 87.577 64.468 ;
			RECT	87.713 64.404 87.745 64.468 ;
			RECT	87.881 64.404 87.913 64.468 ;
			RECT	88.049 64.404 88.081 64.468 ;
			RECT	88.217 64.404 88.249 64.468 ;
			RECT	88.385 64.404 88.417 64.468 ;
			RECT	88.553 64.404 88.585 64.468 ;
			RECT	88.721 64.404 88.753 64.468 ;
			RECT	88.889 64.404 88.921 64.468 ;
			RECT	89.057 64.404 89.089 64.468 ;
			RECT	89.225 64.404 89.257 64.468 ;
			RECT	89.393 64.404 89.425 64.468 ;
			RECT	89.561 64.404 89.593 64.468 ;
			RECT	89.729 64.404 89.761 64.468 ;
			RECT	89.897 64.404 89.929 64.468 ;
			RECT	90.065 64.404 90.097 64.468 ;
			RECT	90.233 64.404 90.265 64.468 ;
			RECT	90.401 64.404 90.433 64.468 ;
			RECT	90.569 64.404 90.601 64.468 ;
			RECT	90.737 64.404 90.769 64.468 ;
			RECT	90.905 64.404 90.937 64.468 ;
			RECT	91.073 64.404 91.105 64.468 ;
			RECT	91.241 64.404 91.273 64.468 ;
			RECT	91.409 64.404 91.441 64.468 ;
			RECT	91.577 64.404 91.609 64.468 ;
			RECT	91.745 64.404 91.777 64.468 ;
			RECT	91.913 64.404 91.945 64.468 ;
			RECT	92.081 64.404 92.113 64.468 ;
			RECT	92.249 64.404 92.281 64.468 ;
			RECT	92.417 64.404 92.449 64.468 ;
			RECT	92.585 64.404 92.617 64.468 ;
			RECT	92.753 64.404 92.785 64.468 ;
			RECT	92.921 64.404 92.953 64.468 ;
			RECT	93.089 64.404 93.121 64.468 ;
			RECT	93.257 64.404 93.289 64.468 ;
			RECT	93.425 64.404 93.457 64.468 ;
			RECT	93.593 64.404 93.625 64.468 ;
			RECT	93.761 64.404 93.793 64.468 ;
			RECT	93.929 64.404 93.961 64.468 ;
			RECT	94.097 64.404 94.129 64.468 ;
			RECT	94.265 64.404 94.297 64.468 ;
			RECT	94.433 64.404 94.465 64.468 ;
			RECT	94.601 64.404 94.633 64.468 ;
			RECT	94.769 64.404 94.801 64.468 ;
			RECT	94.937 64.404 94.969 64.468 ;
			RECT	95.105 64.404 95.137 64.468 ;
			RECT	95.273 64.404 95.305 64.468 ;
			RECT	95.441 64.404 95.473 64.468 ;
			RECT	95.609 64.404 95.641 64.468 ;
			RECT	95.777 64.404 95.809 64.468 ;
			RECT	95.945 64.404 95.977 64.468 ;
			RECT	96.113 64.404 96.145 64.468 ;
			RECT	96.281 64.404 96.313 64.468 ;
			RECT	96.449 64.404 96.481 64.468 ;
			RECT	96.617 64.404 96.649 64.468 ;
			RECT	96.785 64.404 96.817 64.468 ;
			RECT	96.953 64.404 96.985 64.468 ;
			RECT	97.121 64.404 97.153 64.468 ;
			RECT	97.289 64.404 97.321 64.468 ;
			RECT	97.457 64.404 97.489 64.468 ;
			RECT	97.625 64.404 97.657 64.468 ;
			RECT	97.793 64.404 97.825 64.468 ;
			RECT	97.961 64.404 97.993 64.468 ;
			RECT	98.129 64.404 98.161 64.468 ;
			RECT	98.297 64.404 98.329 64.468 ;
			RECT	98.465 64.404 98.497 64.468 ;
			RECT	98.633 64.404 98.665 64.468 ;
			RECT	98.801 64.404 98.833 64.468 ;
			RECT	98.969 64.404 99.001 64.468 ;
			RECT	99.137 64.404 99.169 64.468 ;
			RECT	99.305 64.404 99.337 64.468 ;
			RECT	99.473 64.404 99.505 64.468 ;
			RECT	99.641 64.404 99.673 64.468 ;
			RECT	99.809 64.404 99.841 64.468 ;
			RECT	99.977 64.404 100.009 64.468 ;
			RECT	100.145 64.404 100.177 64.468 ;
			RECT	100.313 64.404 100.345 64.468 ;
			RECT	100.481 64.404 100.513 64.468 ;
			RECT	100.649 64.404 100.681 64.468 ;
			RECT	100.817 64.404 100.849 64.468 ;
			RECT	100.985 64.404 101.017 64.468 ;
			RECT	101.153 64.404 101.185 64.468 ;
			RECT	101.321 64.404 101.353 64.468 ;
			RECT	101.489 64.404 101.521 64.468 ;
			RECT	101.657 64.404 101.689 64.468 ;
			RECT	101.825 64.404 101.857 64.468 ;
			RECT	101.993 64.404 102.025 64.468 ;
			RECT	102.123 64.42 102.155 64.452 ;
			RECT	102.245 64.415 102.277 64.447 ;
			RECT	102.375 64.404 102.407 64.468 ;
			RECT	103.795 64.404 103.827 64.468 ;
			RECT	103.925 64.415 103.957 64.447 ;
			RECT	104.047 64.42 104.079 64.452 ;
			RECT	104.177 64.404 104.209 64.468 ;
			RECT	104.345 64.404 104.377 64.468 ;
			RECT	104.513 64.404 104.545 64.468 ;
			RECT	104.681 64.404 104.713 64.468 ;
			RECT	104.849 64.404 104.881 64.468 ;
			RECT	105.017 64.404 105.049 64.468 ;
			RECT	105.185 64.404 105.217 64.468 ;
			RECT	105.353 64.404 105.385 64.468 ;
			RECT	105.521 64.404 105.553 64.468 ;
			RECT	105.689 64.404 105.721 64.468 ;
			RECT	105.857 64.404 105.889 64.468 ;
			RECT	106.025 64.404 106.057 64.468 ;
			RECT	106.193 64.404 106.225 64.468 ;
			RECT	106.361 64.404 106.393 64.468 ;
			RECT	106.529 64.404 106.561 64.468 ;
			RECT	106.697 64.404 106.729 64.468 ;
			RECT	106.865 64.404 106.897 64.468 ;
			RECT	107.033 64.404 107.065 64.468 ;
			RECT	107.201 64.404 107.233 64.468 ;
			RECT	107.369 64.404 107.401 64.468 ;
			RECT	107.537 64.404 107.569 64.468 ;
			RECT	107.705 64.404 107.737 64.468 ;
			RECT	107.873 64.404 107.905 64.468 ;
			RECT	108.041 64.404 108.073 64.468 ;
			RECT	108.209 64.404 108.241 64.468 ;
			RECT	108.377 64.404 108.409 64.468 ;
			RECT	108.545 64.404 108.577 64.468 ;
			RECT	108.713 64.404 108.745 64.468 ;
			RECT	108.881 64.404 108.913 64.468 ;
			RECT	109.049 64.404 109.081 64.468 ;
			RECT	109.217 64.404 109.249 64.468 ;
			RECT	109.385 64.404 109.417 64.468 ;
			RECT	109.553 64.404 109.585 64.468 ;
			RECT	109.721 64.404 109.753 64.468 ;
			RECT	109.889 64.404 109.921 64.468 ;
			RECT	110.057 64.404 110.089 64.468 ;
			RECT	110.225 64.404 110.257 64.468 ;
			RECT	110.393 64.404 110.425 64.468 ;
			RECT	110.561 64.404 110.593 64.468 ;
			RECT	110.729 64.404 110.761 64.468 ;
			RECT	110.897 64.404 110.929 64.468 ;
			RECT	111.065 64.404 111.097 64.468 ;
			RECT	111.233 64.404 111.265 64.468 ;
			RECT	111.401 64.404 111.433 64.468 ;
			RECT	111.569 64.404 111.601 64.468 ;
			RECT	111.737 64.404 111.769 64.468 ;
			RECT	111.905 64.404 111.937 64.468 ;
			RECT	112.073 64.404 112.105 64.468 ;
			RECT	112.241 64.404 112.273 64.468 ;
			RECT	112.409 64.404 112.441 64.468 ;
			RECT	112.577 64.404 112.609 64.468 ;
			RECT	112.745 64.404 112.777 64.468 ;
			RECT	112.913 64.404 112.945 64.468 ;
			RECT	113.081 64.404 113.113 64.468 ;
			RECT	113.249 64.404 113.281 64.468 ;
			RECT	113.417 64.404 113.449 64.468 ;
			RECT	113.585 64.404 113.617 64.468 ;
			RECT	113.753 64.404 113.785 64.468 ;
			RECT	113.921 64.404 113.953 64.468 ;
			RECT	114.089 64.404 114.121 64.468 ;
			RECT	114.257 64.404 114.289 64.468 ;
			RECT	114.425 64.404 114.457 64.468 ;
			RECT	114.593 64.404 114.625 64.468 ;
			RECT	114.761 64.404 114.793 64.468 ;
			RECT	114.929 64.404 114.961 64.468 ;
			RECT	115.097 64.404 115.129 64.468 ;
			RECT	115.265 64.404 115.297 64.468 ;
			RECT	115.433 64.404 115.465 64.468 ;
			RECT	115.601 64.404 115.633 64.468 ;
			RECT	115.769 64.404 115.801 64.468 ;
			RECT	115.937 64.404 115.969 64.468 ;
			RECT	116.105 64.404 116.137 64.468 ;
			RECT	116.273 64.404 116.305 64.468 ;
			RECT	116.441 64.404 116.473 64.468 ;
			RECT	116.609 64.404 116.641 64.468 ;
			RECT	116.777 64.404 116.809 64.468 ;
			RECT	116.945 64.404 116.977 64.468 ;
			RECT	117.113 64.404 117.145 64.468 ;
			RECT	117.281 64.404 117.313 64.468 ;
			RECT	117.449 64.404 117.481 64.468 ;
			RECT	117.617 64.404 117.649 64.468 ;
			RECT	117.785 64.404 117.817 64.468 ;
			RECT	117.953 64.404 117.985 64.468 ;
			RECT	118.121 64.404 118.153 64.468 ;
			RECT	118.289 64.404 118.321 64.468 ;
			RECT	118.457 64.404 118.489 64.468 ;
			RECT	118.625 64.404 118.657 64.468 ;
			RECT	118.793 64.404 118.825 64.468 ;
			RECT	118.961 64.404 118.993 64.468 ;
			RECT	119.129 64.404 119.161 64.468 ;
			RECT	119.297 64.404 119.329 64.468 ;
			RECT	119.465 64.404 119.497 64.468 ;
			RECT	119.633 64.404 119.665 64.468 ;
			RECT	119.801 64.404 119.833 64.468 ;
			RECT	119.969 64.404 120.001 64.468 ;
			RECT	120.137 64.404 120.169 64.468 ;
			RECT	120.305 64.404 120.337 64.468 ;
			RECT	120.473 64.404 120.505 64.468 ;
			RECT	120.641 64.404 120.673 64.468 ;
			RECT	120.809 64.404 120.841 64.468 ;
			RECT	120.977 64.404 121.009 64.468 ;
			RECT	121.145 64.404 121.177 64.468 ;
			RECT	121.313 64.404 121.345 64.468 ;
			RECT	121.481 64.404 121.513 64.468 ;
			RECT	121.649 64.404 121.681 64.468 ;
			RECT	121.817 64.404 121.849 64.468 ;
			RECT	121.985 64.404 122.017 64.468 ;
			RECT	122.153 64.404 122.185 64.468 ;
			RECT	122.321 64.404 122.353 64.468 ;
			RECT	122.489 64.404 122.521 64.468 ;
			RECT	122.657 64.404 122.689 64.468 ;
			RECT	122.825 64.404 122.857 64.468 ;
			RECT	122.993 64.404 123.025 64.468 ;
			RECT	123.161 64.404 123.193 64.468 ;
			RECT	123.329 64.404 123.361 64.468 ;
			RECT	123.497 64.404 123.529 64.468 ;
			RECT	123.665 64.404 123.697 64.468 ;
			RECT	123.833 64.404 123.865 64.468 ;
			RECT	124.001 64.404 124.033 64.468 ;
			RECT	124.169 64.404 124.201 64.468 ;
			RECT	124.337 64.404 124.369 64.468 ;
			RECT	124.505 64.404 124.537 64.468 ;
			RECT	124.673 64.404 124.705 64.468 ;
			RECT	124.841 64.404 124.873 64.468 ;
			RECT	125.009 64.404 125.041 64.468 ;
			RECT	125.177 64.404 125.209 64.468 ;
			RECT	125.345 64.404 125.377 64.468 ;
			RECT	125.513 64.404 125.545 64.468 ;
			RECT	125.681 64.404 125.713 64.468 ;
			RECT	125.849 64.404 125.881 64.468 ;
			RECT	126.017 64.404 126.049 64.468 ;
			RECT	126.185 64.404 126.217 64.468 ;
			RECT	126.353 64.404 126.385 64.468 ;
			RECT	126.521 64.404 126.553 64.468 ;
			RECT	126.689 64.404 126.721 64.468 ;
			RECT	126.857 64.404 126.889 64.468 ;
			RECT	127.025 64.404 127.057 64.468 ;
			RECT	127.193 64.404 127.225 64.468 ;
			RECT	127.361 64.404 127.393 64.468 ;
			RECT	127.529 64.404 127.561 64.468 ;
			RECT	127.697 64.404 127.729 64.468 ;
			RECT	127.865 64.404 127.897 64.468 ;
			RECT	128.033 64.404 128.065 64.468 ;
			RECT	128.201 64.404 128.233 64.468 ;
			RECT	128.369 64.404 128.401 64.468 ;
			RECT	128.537 64.404 128.569 64.468 ;
			RECT	128.705 64.404 128.737 64.468 ;
			RECT	128.873 64.404 128.905 64.468 ;
			RECT	129.041 64.404 129.073 64.468 ;
			RECT	129.209 64.404 129.241 64.468 ;
			RECT	129.377 64.404 129.409 64.468 ;
			RECT	129.545 64.404 129.577 64.468 ;
			RECT	129.713 64.404 129.745 64.468 ;
			RECT	129.881 64.404 129.913 64.468 ;
			RECT	130.049 64.404 130.081 64.468 ;
			RECT	130.217 64.404 130.249 64.468 ;
			RECT	130.385 64.404 130.417 64.468 ;
			RECT	130.553 64.404 130.585 64.468 ;
			RECT	130.721 64.404 130.753 64.468 ;
			RECT	130.889 64.404 130.921 64.468 ;
			RECT	131.057 64.404 131.089 64.468 ;
			RECT	131.225 64.404 131.257 64.468 ;
			RECT	131.393 64.404 131.425 64.468 ;
			RECT	131.561 64.404 131.593 64.468 ;
			RECT	131.729 64.404 131.761 64.468 ;
			RECT	131.897 64.404 131.929 64.468 ;
			RECT	132.065 64.404 132.097 64.468 ;
			RECT	132.233 64.404 132.265 64.468 ;
			RECT	132.401 64.404 132.433 64.468 ;
			RECT	132.569 64.404 132.601 64.468 ;
			RECT	132.737 64.404 132.769 64.468 ;
			RECT	132.905 64.404 132.937 64.468 ;
			RECT	133.073 64.404 133.105 64.468 ;
			RECT	133.241 64.404 133.273 64.468 ;
			RECT	133.409 64.404 133.441 64.468 ;
			RECT	133.577 64.404 133.609 64.468 ;
			RECT	133.745 64.404 133.777 64.468 ;
			RECT	133.913 64.404 133.945 64.468 ;
			RECT	134.081 64.404 134.113 64.468 ;
			RECT	134.249 64.404 134.281 64.468 ;
			RECT	134.417 64.404 134.449 64.468 ;
			RECT	134.585 64.404 134.617 64.468 ;
			RECT	134.753 64.404 134.785 64.468 ;
			RECT	134.921 64.404 134.953 64.468 ;
			RECT	135.089 64.404 135.121 64.468 ;
			RECT	135.257 64.404 135.289 64.468 ;
			RECT	135.425 64.404 135.457 64.468 ;
			RECT	135.593 64.404 135.625 64.468 ;
			RECT	135.761 64.404 135.793 64.468 ;
			RECT	135.929 64.404 135.961 64.468 ;
			RECT	136.097 64.404 136.129 64.468 ;
			RECT	136.265 64.404 136.297 64.468 ;
			RECT	136.433 64.404 136.465 64.468 ;
			RECT	136.601 64.404 136.633 64.468 ;
			RECT	136.769 64.404 136.801 64.468 ;
			RECT	136.937 64.404 136.969 64.468 ;
			RECT	137.105 64.404 137.137 64.468 ;
			RECT	137.273 64.404 137.305 64.468 ;
			RECT	137.441 64.404 137.473 64.468 ;
			RECT	137.609 64.404 137.641 64.468 ;
			RECT	137.777 64.404 137.809 64.468 ;
			RECT	137.945 64.404 137.977 64.468 ;
			RECT	138.113 64.404 138.145 64.468 ;
			RECT	138.281 64.404 138.313 64.468 ;
			RECT	138.449 64.404 138.481 64.468 ;
			RECT	138.617 64.404 138.649 64.468 ;
			RECT	138.785 64.404 138.817 64.468 ;
			RECT	138.953 64.404 138.985 64.468 ;
			RECT	139.121 64.404 139.153 64.468 ;
			RECT	139.289 64.404 139.321 64.468 ;
			RECT	139.457 64.404 139.489 64.468 ;
			RECT	139.625 64.404 139.657 64.468 ;
			RECT	139.793 64.404 139.825 64.468 ;
			RECT	139.961 64.404 139.993 64.468 ;
			RECT	140.129 64.404 140.161 64.468 ;
			RECT	140.297 64.404 140.329 64.468 ;
			RECT	140.465 64.404 140.497 64.468 ;
			RECT	140.633 64.404 140.665 64.468 ;
			RECT	140.801 64.404 140.833 64.468 ;
			RECT	140.969 64.404 141.001 64.468 ;
			RECT	141.137 64.404 141.169 64.468 ;
			RECT	141.305 64.404 141.337 64.468 ;
			RECT	141.473 64.404 141.505 64.468 ;
			RECT	141.641 64.404 141.673 64.468 ;
			RECT	141.809 64.404 141.841 64.468 ;
			RECT	141.977 64.404 142.009 64.468 ;
			RECT	142.145 64.404 142.177 64.468 ;
			RECT	142.313 64.404 142.345 64.468 ;
			RECT	142.481 64.404 142.513 64.468 ;
			RECT	142.649 64.404 142.681 64.468 ;
			RECT	142.817 64.404 142.849 64.468 ;
			RECT	142.985 64.404 143.017 64.468 ;
			RECT	143.153 64.404 143.185 64.468 ;
			RECT	143.321 64.404 143.353 64.468 ;
			RECT	143.489 64.404 143.521 64.468 ;
			RECT	143.657 64.404 143.689 64.468 ;
			RECT	143.825 64.404 143.857 64.468 ;
			RECT	143.993 64.404 144.025 64.468 ;
			RECT	144.161 64.404 144.193 64.468 ;
			RECT	144.329 64.404 144.361 64.468 ;
			RECT	144.497 64.404 144.529 64.468 ;
			RECT	144.665 64.404 144.697 64.468 ;
			RECT	144.833 64.404 144.865 64.468 ;
			RECT	145.001 64.404 145.033 64.468 ;
			RECT	145.169 64.404 145.201 64.468 ;
			RECT	145.337 64.404 145.369 64.468 ;
			RECT	145.505 64.404 145.537 64.468 ;
			RECT	145.673 64.404 145.705 64.468 ;
			RECT	145.841 64.404 145.873 64.468 ;
			RECT	146.009 64.404 146.041 64.468 ;
			RECT	146.177 64.404 146.209 64.468 ;
			RECT	146.345 64.404 146.377 64.468 ;
			RECT	146.513 64.404 146.545 64.468 ;
			RECT	146.681 64.404 146.713 64.468 ;
			RECT	146.849 64.404 146.881 64.468 ;
			RECT	147.017 64.404 147.049 64.468 ;
			RECT	147.185 64.404 147.217 64.468 ;
			RECT	147.316 64.42 147.348 64.452 ;
			RECT	147.437 64.42 147.469 64.452 ;
			RECT	147.567 64.404 147.599 64.468 ;
			RECT	149.879 64.404 149.911 64.468 ;
			RECT	151.13 64.404 151.194 64.468 ;
			RECT	151.81 64.404 151.842 64.468 ;
			RECT	152.249 64.404 152.281 64.468 ;
			RECT	153.56 64.404 153.624 64.468 ;
			RECT	156.601 64.404 156.633 64.468 ;
			RECT	156.731 64.42 156.763 64.452 ;
			RECT	156.852 64.42 156.884 64.452 ;
			RECT	156.983 64.404 157.015 64.468 ;
			RECT	157.151 64.404 157.183 64.468 ;
			RECT	157.319 64.404 157.351 64.468 ;
			RECT	157.487 64.404 157.519 64.468 ;
			RECT	157.655 64.404 157.687 64.468 ;
			RECT	157.823 64.404 157.855 64.468 ;
			RECT	157.991 64.404 158.023 64.468 ;
			RECT	158.159 64.404 158.191 64.468 ;
			RECT	158.327 64.404 158.359 64.468 ;
			RECT	158.495 64.404 158.527 64.468 ;
			RECT	158.663 64.404 158.695 64.468 ;
			RECT	158.831 64.404 158.863 64.468 ;
			RECT	158.999 64.404 159.031 64.468 ;
			RECT	159.167 64.404 159.199 64.468 ;
			RECT	159.335 64.404 159.367 64.468 ;
			RECT	159.503 64.404 159.535 64.468 ;
			RECT	159.671 64.404 159.703 64.468 ;
			RECT	159.839 64.404 159.871 64.468 ;
			RECT	160.007 64.404 160.039 64.468 ;
			RECT	160.175 64.404 160.207 64.468 ;
			RECT	160.343 64.404 160.375 64.468 ;
			RECT	160.511 64.404 160.543 64.468 ;
			RECT	160.679 64.404 160.711 64.468 ;
			RECT	160.847 64.404 160.879 64.468 ;
			RECT	161.015 64.404 161.047 64.468 ;
			RECT	161.183 64.404 161.215 64.468 ;
			RECT	161.351 64.404 161.383 64.468 ;
			RECT	161.519 64.404 161.551 64.468 ;
			RECT	161.687 64.404 161.719 64.468 ;
			RECT	161.855 64.404 161.887 64.468 ;
			RECT	162.023 64.404 162.055 64.468 ;
			RECT	162.191 64.404 162.223 64.468 ;
			RECT	162.359 64.404 162.391 64.468 ;
			RECT	162.527 64.404 162.559 64.468 ;
			RECT	162.695 64.404 162.727 64.468 ;
			RECT	162.863 64.404 162.895 64.468 ;
			RECT	163.031 64.404 163.063 64.468 ;
			RECT	163.199 64.404 163.231 64.468 ;
			RECT	163.367 64.404 163.399 64.468 ;
			RECT	163.535 64.404 163.567 64.468 ;
			RECT	163.703 64.404 163.735 64.468 ;
			RECT	163.871 64.404 163.903 64.468 ;
			RECT	164.039 64.404 164.071 64.468 ;
			RECT	164.207 64.404 164.239 64.468 ;
			RECT	164.375 64.404 164.407 64.468 ;
			RECT	164.543 64.404 164.575 64.468 ;
			RECT	164.711 64.404 164.743 64.468 ;
			RECT	164.879 64.404 164.911 64.468 ;
			RECT	165.047 64.404 165.079 64.468 ;
			RECT	165.215 64.404 165.247 64.468 ;
			RECT	165.383 64.404 165.415 64.468 ;
			RECT	165.551 64.404 165.583 64.468 ;
			RECT	165.719 64.404 165.751 64.468 ;
			RECT	165.887 64.404 165.919 64.468 ;
			RECT	166.055 64.404 166.087 64.468 ;
			RECT	166.223 64.404 166.255 64.468 ;
			RECT	166.391 64.404 166.423 64.468 ;
			RECT	166.559 64.404 166.591 64.468 ;
			RECT	166.727 64.404 166.759 64.468 ;
			RECT	166.895 64.404 166.927 64.468 ;
			RECT	167.063 64.404 167.095 64.468 ;
			RECT	167.231 64.404 167.263 64.468 ;
			RECT	167.399 64.404 167.431 64.468 ;
			RECT	167.567 64.404 167.599 64.468 ;
			RECT	167.735 64.404 167.767 64.468 ;
			RECT	167.903 64.404 167.935 64.468 ;
			RECT	168.071 64.404 168.103 64.468 ;
			RECT	168.239 64.404 168.271 64.468 ;
			RECT	168.407 64.404 168.439 64.468 ;
			RECT	168.575 64.404 168.607 64.468 ;
			RECT	168.743 64.404 168.775 64.468 ;
			RECT	168.911 64.404 168.943 64.468 ;
			RECT	169.079 64.404 169.111 64.468 ;
			RECT	169.247 64.404 169.279 64.468 ;
			RECT	169.415 64.404 169.447 64.468 ;
			RECT	169.583 64.404 169.615 64.468 ;
			RECT	169.751 64.404 169.783 64.468 ;
			RECT	169.919 64.404 169.951 64.468 ;
			RECT	170.087 64.404 170.119 64.468 ;
			RECT	170.255 64.404 170.287 64.468 ;
			RECT	170.423 64.404 170.455 64.468 ;
			RECT	170.591 64.404 170.623 64.468 ;
			RECT	170.759 64.404 170.791 64.468 ;
			RECT	170.927 64.404 170.959 64.468 ;
			RECT	171.095 64.404 171.127 64.468 ;
			RECT	171.263 64.404 171.295 64.468 ;
			RECT	171.431 64.404 171.463 64.468 ;
			RECT	171.599 64.404 171.631 64.468 ;
			RECT	171.767 64.404 171.799 64.468 ;
			RECT	171.935 64.404 171.967 64.468 ;
			RECT	172.103 64.404 172.135 64.468 ;
			RECT	172.271 64.404 172.303 64.468 ;
			RECT	172.439 64.404 172.471 64.468 ;
			RECT	172.607 64.404 172.639 64.468 ;
			RECT	172.775 64.404 172.807 64.468 ;
			RECT	172.943 64.404 172.975 64.468 ;
			RECT	173.111 64.404 173.143 64.468 ;
			RECT	173.279 64.404 173.311 64.468 ;
			RECT	173.447 64.404 173.479 64.468 ;
			RECT	173.615 64.404 173.647 64.468 ;
			RECT	173.783 64.404 173.815 64.468 ;
			RECT	173.951 64.404 173.983 64.468 ;
			RECT	174.119 64.404 174.151 64.468 ;
			RECT	174.287 64.404 174.319 64.468 ;
			RECT	174.455 64.404 174.487 64.468 ;
			RECT	174.623 64.404 174.655 64.468 ;
			RECT	174.791 64.404 174.823 64.468 ;
			RECT	174.959 64.404 174.991 64.468 ;
			RECT	175.127 64.404 175.159 64.468 ;
			RECT	175.295 64.404 175.327 64.468 ;
			RECT	175.463 64.404 175.495 64.468 ;
			RECT	175.631 64.404 175.663 64.468 ;
			RECT	175.799 64.404 175.831 64.468 ;
			RECT	175.967 64.404 175.999 64.468 ;
			RECT	176.135 64.404 176.167 64.468 ;
			RECT	176.303 64.404 176.335 64.468 ;
			RECT	176.471 64.404 176.503 64.468 ;
			RECT	176.639 64.404 176.671 64.468 ;
			RECT	176.807 64.404 176.839 64.468 ;
			RECT	176.975 64.404 177.007 64.468 ;
			RECT	177.143 64.404 177.175 64.468 ;
			RECT	177.311 64.404 177.343 64.468 ;
			RECT	177.479 64.404 177.511 64.468 ;
			RECT	177.647 64.404 177.679 64.468 ;
			RECT	177.815 64.404 177.847 64.468 ;
			RECT	177.983 64.404 178.015 64.468 ;
			RECT	178.151 64.404 178.183 64.468 ;
			RECT	178.319 64.404 178.351 64.468 ;
			RECT	178.487 64.404 178.519 64.468 ;
			RECT	178.655 64.404 178.687 64.468 ;
			RECT	178.823 64.404 178.855 64.468 ;
			RECT	178.991 64.404 179.023 64.468 ;
			RECT	179.159 64.404 179.191 64.468 ;
			RECT	179.327 64.404 179.359 64.468 ;
			RECT	179.495 64.404 179.527 64.468 ;
			RECT	179.663 64.404 179.695 64.468 ;
			RECT	179.831 64.404 179.863 64.468 ;
			RECT	179.999 64.404 180.031 64.468 ;
			RECT	180.167 64.404 180.199 64.468 ;
			RECT	180.335 64.404 180.367 64.468 ;
			RECT	180.503 64.404 180.535 64.468 ;
			RECT	180.671 64.404 180.703 64.468 ;
			RECT	180.839 64.404 180.871 64.468 ;
			RECT	181.007 64.404 181.039 64.468 ;
			RECT	181.175 64.404 181.207 64.468 ;
			RECT	181.343 64.404 181.375 64.468 ;
			RECT	181.511 64.404 181.543 64.468 ;
			RECT	181.679 64.404 181.711 64.468 ;
			RECT	181.847 64.404 181.879 64.468 ;
			RECT	182.015 64.404 182.047 64.468 ;
			RECT	182.183 64.404 182.215 64.468 ;
			RECT	182.351 64.404 182.383 64.468 ;
			RECT	182.519 64.404 182.551 64.468 ;
			RECT	182.687 64.404 182.719 64.468 ;
			RECT	182.855 64.404 182.887 64.468 ;
			RECT	183.023 64.404 183.055 64.468 ;
			RECT	183.191 64.404 183.223 64.468 ;
			RECT	183.359 64.404 183.391 64.468 ;
			RECT	183.527 64.404 183.559 64.468 ;
			RECT	183.695 64.404 183.727 64.468 ;
			RECT	183.863 64.404 183.895 64.468 ;
			RECT	184.031 64.404 184.063 64.468 ;
			RECT	184.199 64.404 184.231 64.468 ;
			RECT	184.367 64.404 184.399 64.468 ;
			RECT	184.535 64.404 184.567 64.468 ;
			RECT	184.703 64.404 184.735 64.468 ;
			RECT	184.871 64.404 184.903 64.468 ;
			RECT	185.039 64.404 185.071 64.468 ;
			RECT	185.207 64.404 185.239 64.468 ;
			RECT	185.375 64.404 185.407 64.468 ;
			RECT	185.543 64.404 185.575 64.468 ;
			RECT	185.711 64.404 185.743 64.468 ;
			RECT	185.879 64.404 185.911 64.468 ;
			RECT	186.047 64.404 186.079 64.468 ;
			RECT	186.215 64.404 186.247 64.468 ;
			RECT	186.383 64.404 186.415 64.468 ;
			RECT	186.551 64.404 186.583 64.468 ;
			RECT	186.719 64.404 186.751 64.468 ;
			RECT	186.887 64.404 186.919 64.468 ;
			RECT	187.055 64.404 187.087 64.468 ;
			RECT	187.223 64.404 187.255 64.468 ;
			RECT	187.391 64.404 187.423 64.468 ;
			RECT	187.559 64.404 187.591 64.468 ;
			RECT	187.727 64.404 187.759 64.468 ;
			RECT	187.895 64.404 187.927 64.468 ;
			RECT	188.063 64.404 188.095 64.468 ;
			RECT	188.231 64.404 188.263 64.468 ;
			RECT	188.399 64.404 188.431 64.468 ;
			RECT	188.567 64.404 188.599 64.468 ;
			RECT	188.735 64.404 188.767 64.468 ;
			RECT	188.903 64.404 188.935 64.468 ;
			RECT	189.071 64.404 189.103 64.468 ;
			RECT	189.239 64.404 189.271 64.468 ;
			RECT	189.407 64.404 189.439 64.468 ;
			RECT	189.575 64.404 189.607 64.468 ;
			RECT	189.743 64.404 189.775 64.468 ;
			RECT	189.911 64.404 189.943 64.468 ;
			RECT	190.079 64.404 190.111 64.468 ;
			RECT	190.247 64.404 190.279 64.468 ;
			RECT	190.415 64.404 190.447 64.468 ;
			RECT	190.583 64.404 190.615 64.468 ;
			RECT	190.751 64.404 190.783 64.468 ;
			RECT	190.919 64.404 190.951 64.468 ;
			RECT	191.087 64.404 191.119 64.468 ;
			RECT	191.255 64.404 191.287 64.468 ;
			RECT	191.423 64.404 191.455 64.468 ;
			RECT	191.591 64.404 191.623 64.468 ;
			RECT	191.759 64.404 191.791 64.468 ;
			RECT	191.927 64.404 191.959 64.468 ;
			RECT	192.095 64.404 192.127 64.468 ;
			RECT	192.263 64.404 192.295 64.468 ;
			RECT	192.431 64.404 192.463 64.468 ;
			RECT	192.599 64.404 192.631 64.468 ;
			RECT	192.767 64.404 192.799 64.468 ;
			RECT	192.935 64.404 192.967 64.468 ;
			RECT	193.103 64.404 193.135 64.468 ;
			RECT	193.271 64.404 193.303 64.468 ;
			RECT	193.439 64.404 193.471 64.468 ;
			RECT	193.607 64.404 193.639 64.468 ;
			RECT	193.775 64.404 193.807 64.468 ;
			RECT	193.943 64.404 193.975 64.468 ;
			RECT	194.111 64.404 194.143 64.468 ;
			RECT	194.279 64.404 194.311 64.468 ;
			RECT	194.447 64.404 194.479 64.468 ;
			RECT	194.615 64.404 194.647 64.468 ;
			RECT	194.783 64.404 194.815 64.468 ;
			RECT	194.951 64.404 194.983 64.468 ;
			RECT	195.119 64.404 195.151 64.468 ;
			RECT	195.287 64.404 195.319 64.468 ;
			RECT	195.455 64.404 195.487 64.468 ;
			RECT	195.623 64.404 195.655 64.468 ;
			RECT	195.791 64.404 195.823 64.468 ;
			RECT	195.959 64.404 195.991 64.468 ;
			RECT	196.127 64.404 196.159 64.468 ;
			RECT	196.295 64.404 196.327 64.468 ;
			RECT	196.463 64.404 196.495 64.468 ;
			RECT	196.631 64.404 196.663 64.468 ;
			RECT	196.799 64.404 196.831 64.468 ;
			RECT	196.967 64.404 196.999 64.468 ;
			RECT	197.135 64.404 197.167 64.468 ;
			RECT	197.303 64.404 197.335 64.468 ;
			RECT	197.471 64.404 197.503 64.468 ;
			RECT	197.639 64.404 197.671 64.468 ;
			RECT	197.807 64.404 197.839 64.468 ;
			RECT	197.975 64.404 198.007 64.468 ;
			RECT	198.143 64.404 198.175 64.468 ;
			RECT	198.311 64.404 198.343 64.468 ;
			RECT	198.479 64.404 198.511 64.468 ;
			RECT	198.647 64.404 198.679 64.468 ;
			RECT	198.815 64.404 198.847 64.468 ;
			RECT	198.983 64.404 199.015 64.468 ;
			RECT	199.151 64.404 199.183 64.468 ;
			RECT	199.319 64.404 199.351 64.468 ;
			RECT	199.487 64.404 199.519 64.468 ;
			RECT	199.655 64.404 199.687 64.468 ;
			RECT	199.823 64.404 199.855 64.468 ;
			RECT	199.991 64.404 200.023 64.468 ;
			RECT	200.121 64.42 200.153 64.452 ;
			RECT	200.243 64.415 200.275 64.447 ;
			RECT	200.373 64.404 200.405 64.468 ;
			RECT	200.9 64.404 200.932 64.468 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 62.456 201.665 62.576 ;
			LAYER	J3 ;
			RECT	0.755 62.484 0.787 62.548 ;
			RECT	1.645 62.484 1.709 62.548 ;
			RECT	2.323 62.484 2.387 62.548 ;
			RECT	3.438 62.484 3.47 62.548 ;
			RECT	3.585 62.484 3.617 62.548 ;
			RECT	4.195 62.484 4.227 62.548 ;
			RECT	4.72 62.484 4.752 62.548 ;
			RECT	4.944 62.484 5.008 62.548 ;
			RECT	5.267 62.484 5.299 62.548 ;
			RECT	5.797 62.484 5.829 62.548 ;
			RECT	5.927 62.495 5.959 62.527 ;
			RECT	6.049 62.5 6.081 62.532 ;
			RECT	6.179 62.484 6.211 62.548 ;
			RECT	6.347 62.484 6.379 62.548 ;
			RECT	6.515 62.484 6.547 62.548 ;
			RECT	6.683 62.484 6.715 62.548 ;
			RECT	6.851 62.484 6.883 62.548 ;
			RECT	7.019 62.484 7.051 62.548 ;
			RECT	7.187 62.484 7.219 62.548 ;
			RECT	7.355 62.484 7.387 62.548 ;
			RECT	7.523 62.484 7.555 62.548 ;
			RECT	7.691 62.484 7.723 62.548 ;
			RECT	7.859 62.484 7.891 62.548 ;
			RECT	8.027 62.484 8.059 62.548 ;
			RECT	8.195 62.484 8.227 62.548 ;
			RECT	8.363 62.484 8.395 62.548 ;
			RECT	8.531 62.484 8.563 62.548 ;
			RECT	8.699 62.484 8.731 62.548 ;
			RECT	8.867 62.484 8.899 62.548 ;
			RECT	9.035 62.484 9.067 62.548 ;
			RECT	9.203 62.484 9.235 62.548 ;
			RECT	9.371 62.484 9.403 62.548 ;
			RECT	9.539 62.484 9.571 62.548 ;
			RECT	9.707 62.484 9.739 62.548 ;
			RECT	9.875 62.484 9.907 62.548 ;
			RECT	10.043 62.484 10.075 62.548 ;
			RECT	10.211 62.484 10.243 62.548 ;
			RECT	10.379 62.484 10.411 62.548 ;
			RECT	10.547 62.484 10.579 62.548 ;
			RECT	10.715 62.484 10.747 62.548 ;
			RECT	10.883 62.484 10.915 62.548 ;
			RECT	11.051 62.484 11.083 62.548 ;
			RECT	11.219 62.484 11.251 62.548 ;
			RECT	11.387 62.484 11.419 62.548 ;
			RECT	11.555 62.484 11.587 62.548 ;
			RECT	11.723 62.484 11.755 62.548 ;
			RECT	11.891 62.484 11.923 62.548 ;
			RECT	12.059 62.484 12.091 62.548 ;
			RECT	12.227 62.484 12.259 62.548 ;
			RECT	12.395 62.484 12.427 62.548 ;
			RECT	12.563 62.484 12.595 62.548 ;
			RECT	12.731 62.484 12.763 62.548 ;
			RECT	12.899 62.484 12.931 62.548 ;
			RECT	13.067 62.484 13.099 62.548 ;
			RECT	13.235 62.484 13.267 62.548 ;
			RECT	13.403 62.484 13.435 62.548 ;
			RECT	13.571 62.484 13.603 62.548 ;
			RECT	13.739 62.484 13.771 62.548 ;
			RECT	13.907 62.484 13.939 62.548 ;
			RECT	14.075 62.484 14.107 62.548 ;
			RECT	14.243 62.484 14.275 62.548 ;
			RECT	14.411 62.484 14.443 62.548 ;
			RECT	14.579 62.484 14.611 62.548 ;
			RECT	14.747 62.484 14.779 62.548 ;
			RECT	14.915 62.484 14.947 62.548 ;
			RECT	15.083 62.484 15.115 62.548 ;
			RECT	15.251 62.484 15.283 62.548 ;
			RECT	15.419 62.484 15.451 62.548 ;
			RECT	15.587 62.484 15.619 62.548 ;
			RECT	15.755 62.484 15.787 62.548 ;
			RECT	15.923 62.484 15.955 62.548 ;
			RECT	16.091 62.484 16.123 62.548 ;
			RECT	16.259 62.484 16.291 62.548 ;
			RECT	16.427 62.484 16.459 62.548 ;
			RECT	16.595 62.484 16.627 62.548 ;
			RECT	16.763 62.484 16.795 62.548 ;
			RECT	16.931 62.484 16.963 62.548 ;
			RECT	17.099 62.484 17.131 62.548 ;
			RECT	17.267 62.484 17.299 62.548 ;
			RECT	17.435 62.484 17.467 62.548 ;
			RECT	17.603 62.484 17.635 62.548 ;
			RECT	17.771 62.484 17.803 62.548 ;
			RECT	17.939 62.484 17.971 62.548 ;
			RECT	18.107 62.484 18.139 62.548 ;
			RECT	18.275 62.484 18.307 62.548 ;
			RECT	18.443 62.484 18.475 62.548 ;
			RECT	18.611 62.484 18.643 62.548 ;
			RECT	18.779 62.484 18.811 62.548 ;
			RECT	18.947 62.484 18.979 62.548 ;
			RECT	19.115 62.484 19.147 62.548 ;
			RECT	19.283 62.484 19.315 62.548 ;
			RECT	19.451 62.484 19.483 62.548 ;
			RECT	19.619 62.484 19.651 62.548 ;
			RECT	19.787 62.484 19.819 62.548 ;
			RECT	19.955 62.484 19.987 62.548 ;
			RECT	20.123 62.484 20.155 62.548 ;
			RECT	20.291 62.484 20.323 62.548 ;
			RECT	20.459 62.484 20.491 62.548 ;
			RECT	20.627 62.484 20.659 62.548 ;
			RECT	20.795 62.484 20.827 62.548 ;
			RECT	20.963 62.484 20.995 62.548 ;
			RECT	21.131 62.484 21.163 62.548 ;
			RECT	21.299 62.484 21.331 62.548 ;
			RECT	21.467 62.484 21.499 62.548 ;
			RECT	21.635 62.484 21.667 62.548 ;
			RECT	21.803 62.484 21.835 62.548 ;
			RECT	21.971 62.484 22.003 62.548 ;
			RECT	22.139 62.484 22.171 62.548 ;
			RECT	22.307 62.484 22.339 62.548 ;
			RECT	22.475 62.484 22.507 62.548 ;
			RECT	22.643 62.484 22.675 62.548 ;
			RECT	22.811 62.484 22.843 62.548 ;
			RECT	22.979 62.484 23.011 62.548 ;
			RECT	23.147 62.484 23.179 62.548 ;
			RECT	23.315 62.484 23.347 62.548 ;
			RECT	23.483 62.484 23.515 62.548 ;
			RECT	23.651 62.484 23.683 62.548 ;
			RECT	23.819 62.484 23.851 62.548 ;
			RECT	23.987 62.484 24.019 62.548 ;
			RECT	24.155 62.484 24.187 62.548 ;
			RECT	24.323 62.484 24.355 62.548 ;
			RECT	24.491 62.484 24.523 62.548 ;
			RECT	24.659 62.484 24.691 62.548 ;
			RECT	24.827 62.484 24.859 62.548 ;
			RECT	24.995 62.484 25.027 62.548 ;
			RECT	25.163 62.484 25.195 62.548 ;
			RECT	25.331 62.484 25.363 62.548 ;
			RECT	25.499 62.484 25.531 62.548 ;
			RECT	25.667 62.484 25.699 62.548 ;
			RECT	25.835 62.484 25.867 62.548 ;
			RECT	26.003 62.484 26.035 62.548 ;
			RECT	26.171 62.484 26.203 62.548 ;
			RECT	26.339 62.484 26.371 62.548 ;
			RECT	26.507 62.484 26.539 62.548 ;
			RECT	26.675 62.484 26.707 62.548 ;
			RECT	26.843 62.484 26.875 62.548 ;
			RECT	27.011 62.484 27.043 62.548 ;
			RECT	27.179 62.484 27.211 62.548 ;
			RECT	27.347 62.484 27.379 62.548 ;
			RECT	27.515 62.484 27.547 62.548 ;
			RECT	27.683 62.484 27.715 62.548 ;
			RECT	27.851 62.484 27.883 62.548 ;
			RECT	28.019 62.484 28.051 62.548 ;
			RECT	28.187 62.484 28.219 62.548 ;
			RECT	28.355 62.484 28.387 62.548 ;
			RECT	28.523 62.484 28.555 62.548 ;
			RECT	28.691 62.484 28.723 62.548 ;
			RECT	28.859 62.484 28.891 62.548 ;
			RECT	29.027 62.484 29.059 62.548 ;
			RECT	29.195 62.484 29.227 62.548 ;
			RECT	29.363 62.484 29.395 62.548 ;
			RECT	29.531 62.484 29.563 62.548 ;
			RECT	29.699 62.484 29.731 62.548 ;
			RECT	29.867 62.484 29.899 62.548 ;
			RECT	30.035 62.484 30.067 62.548 ;
			RECT	30.203 62.484 30.235 62.548 ;
			RECT	30.371 62.484 30.403 62.548 ;
			RECT	30.539 62.484 30.571 62.548 ;
			RECT	30.707 62.484 30.739 62.548 ;
			RECT	30.875 62.484 30.907 62.548 ;
			RECT	31.043 62.484 31.075 62.548 ;
			RECT	31.211 62.484 31.243 62.548 ;
			RECT	31.379 62.484 31.411 62.548 ;
			RECT	31.547 62.484 31.579 62.548 ;
			RECT	31.715 62.484 31.747 62.548 ;
			RECT	31.883 62.484 31.915 62.548 ;
			RECT	32.051 62.484 32.083 62.548 ;
			RECT	32.219 62.484 32.251 62.548 ;
			RECT	32.387 62.484 32.419 62.548 ;
			RECT	32.555 62.484 32.587 62.548 ;
			RECT	32.723 62.484 32.755 62.548 ;
			RECT	32.891 62.484 32.923 62.548 ;
			RECT	33.059 62.484 33.091 62.548 ;
			RECT	33.227 62.484 33.259 62.548 ;
			RECT	33.395 62.484 33.427 62.548 ;
			RECT	33.563 62.484 33.595 62.548 ;
			RECT	33.731 62.484 33.763 62.548 ;
			RECT	33.899 62.484 33.931 62.548 ;
			RECT	34.067 62.484 34.099 62.548 ;
			RECT	34.235 62.484 34.267 62.548 ;
			RECT	34.403 62.484 34.435 62.548 ;
			RECT	34.571 62.484 34.603 62.548 ;
			RECT	34.739 62.484 34.771 62.548 ;
			RECT	34.907 62.484 34.939 62.548 ;
			RECT	35.075 62.484 35.107 62.548 ;
			RECT	35.243 62.484 35.275 62.548 ;
			RECT	35.411 62.484 35.443 62.548 ;
			RECT	35.579 62.484 35.611 62.548 ;
			RECT	35.747 62.484 35.779 62.548 ;
			RECT	35.915 62.484 35.947 62.548 ;
			RECT	36.083 62.484 36.115 62.548 ;
			RECT	36.251 62.484 36.283 62.548 ;
			RECT	36.419 62.484 36.451 62.548 ;
			RECT	36.587 62.484 36.619 62.548 ;
			RECT	36.755 62.484 36.787 62.548 ;
			RECT	36.923 62.484 36.955 62.548 ;
			RECT	37.091 62.484 37.123 62.548 ;
			RECT	37.259 62.484 37.291 62.548 ;
			RECT	37.427 62.484 37.459 62.548 ;
			RECT	37.595 62.484 37.627 62.548 ;
			RECT	37.763 62.484 37.795 62.548 ;
			RECT	37.931 62.484 37.963 62.548 ;
			RECT	38.099 62.484 38.131 62.548 ;
			RECT	38.267 62.484 38.299 62.548 ;
			RECT	38.435 62.484 38.467 62.548 ;
			RECT	38.603 62.484 38.635 62.548 ;
			RECT	38.771 62.484 38.803 62.548 ;
			RECT	38.939 62.484 38.971 62.548 ;
			RECT	39.107 62.484 39.139 62.548 ;
			RECT	39.275 62.484 39.307 62.548 ;
			RECT	39.443 62.484 39.475 62.548 ;
			RECT	39.611 62.484 39.643 62.548 ;
			RECT	39.779 62.484 39.811 62.548 ;
			RECT	39.947 62.484 39.979 62.548 ;
			RECT	40.115 62.484 40.147 62.548 ;
			RECT	40.283 62.484 40.315 62.548 ;
			RECT	40.451 62.484 40.483 62.548 ;
			RECT	40.619 62.484 40.651 62.548 ;
			RECT	40.787 62.484 40.819 62.548 ;
			RECT	40.955 62.484 40.987 62.548 ;
			RECT	41.123 62.484 41.155 62.548 ;
			RECT	41.291 62.484 41.323 62.548 ;
			RECT	41.459 62.484 41.491 62.548 ;
			RECT	41.627 62.484 41.659 62.548 ;
			RECT	41.795 62.484 41.827 62.548 ;
			RECT	41.963 62.484 41.995 62.548 ;
			RECT	42.131 62.484 42.163 62.548 ;
			RECT	42.299 62.484 42.331 62.548 ;
			RECT	42.467 62.484 42.499 62.548 ;
			RECT	42.635 62.484 42.667 62.548 ;
			RECT	42.803 62.484 42.835 62.548 ;
			RECT	42.971 62.484 43.003 62.548 ;
			RECT	43.139 62.484 43.171 62.548 ;
			RECT	43.307 62.484 43.339 62.548 ;
			RECT	43.475 62.484 43.507 62.548 ;
			RECT	43.643 62.484 43.675 62.548 ;
			RECT	43.811 62.484 43.843 62.548 ;
			RECT	43.979 62.484 44.011 62.548 ;
			RECT	44.147 62.484 44.179 62.548 ;
			RECT	44.315 62.484 44.347 62.548 ;
			RECT	44.483 62.484 44.515 62.548 ;
			RECT	44.651 62.484 44.683 62.548 ;
			RECT	44.819 62.484 44.851 62.548 ;
			RECT	44.987 62.484 45.019 62.548 ;
			RECT	45.155 62.484 45.187 62.548 ;
			RECT	45.323 62.484 45.355 62.548 ;
			RECT	45.491 62.484 45.523 62.548 ;
			RECT	45.659 62.484 45.691 62.548 ;
			RECT	45.827 62.484 45.859 62.548 ;
			RECT	45.995 62.484 46.027 62.548 ;
			RECT	46.163 62.484 46.195 62.548 ;
			RECT	46.331 62.484 46.363 62.548 ;
			RECT	46.499 62.484 46.531 62.548 ;
			RECT	46.667 62.484 46.699 62.548 ;
			RECT	46.835 62.484 46.867 62.548 ;
			RECT	47.003 62.484 47.035 62.548 ;
			RECT	47.171 62.484 47.203 62.548 ;
			RECT	47.339 62.484 47.371 62.548 ;
			RECT	47.507 62.484 47.539 62.548 ;
			RECT	47.675 62.484 47.707 62.548 ;
			RECT	47.843 62.484 47.875 62.548 ;
			RECT	48.011 62.484 48.043 62.548 ;
			RECT	48.179 62.484 48.211 62.548 ;
			RECT	48.347 62.484 48.379 62.548 ;
			RECT	48.515 62.484 48.547 62.548 ;
			RECT	48.683 62.484 48.715 62.548 ;
			RECT	48.851 62.484 48.883 62.548 ;
			RECT	49.019 62.484 49.051 62.548 ;
			RECT	49.187 62.484 49.219 62.548 ;
			RECT	49.318 62.5 49.35 62.532 ;
			RECT	49.439 62.5 49.471 62.532 ;
			RECT	49.569 62.484 49.601 62.548 ;
			RECT	51.881 62.484 51.913 62.548 ;
			RECT	53.132 62.484 53.196 62.548 ;
			RECT	53.812 62.484 53.844 62.548 ;
			RECT	54.251 62.484 54.283 62.548 ;
			RECT	55.562 62.484 55.626 62.548 ;
			RECT	58.603 62.484 58.635 62.548 ;
			RECT	58.733 62.5 58.765 62.532 ;
			RECT	58.854 62.5 58.886 62.532 ;
			RECT	58.985 62.484 59.017 62.548 ;
			RECT	59.153 62.484 59.185 62.548 ;
			RECT	59.321 62.484 59.353 62.548 ;
			RECT	59.489 62.484 59.521 62.548 ;
			RECT	59.657 62.484 59.689 62.548 ;
			RECT	59.825 62.484 59.857 62.548 ;
			RECT	59.993 62.484 60.025 62.548 ;
			RECT	60.161 62.484 60.193 62.548 ;
			RECT	60.329 62.484 60.361 62.548 ;
			RECT	60.497 62.484 60.529 62.548 ;
			RECT	60.665 62.484 60.697 62.548 ;
			RECT	60.833 62.484 60.865 62.548 ;
			RECT	61.001 62.484 61.033 62.548 ;
			RECT	61.169 62.484 61.201 62.548 ;
			RECT	61.337 62.484 61.369 62.548 ;
			RECT	61.505 62.484 61.537 62.548 ;
			RECT	61.673 62.484 61.705 62.548 ;
			RECT	61.841 62.484 61.873 62.548 ;
			RECT	62.009 62.484 62.041 62.548 ;
			RECT	62.177 62.484 62.209 62.548 ;
			RECT	62.345 62.484 62.377 62.548 ;
			RECT	62.513 62.484 62.545 62.548 ;
			RECT	62.681 62.484 62.713 62.548 ;
			RECT	62.849 62.484 62.881 62.548 ;
			RECT	63.017 62.484 63.049 62.548 ;
			RECT	63.185 62.484 63.217 62.548 ;
			RECT	63.353 62.484 63.385 62.548 ;
			RECT	63.521 62.484 63.553 62.548 ;
			RECT	63.689 62.484 63.721 62.548 ;
			RECT	63.857 62.484 63.889 62.548 ;
			RECT	64.025 62.484 64.057 62.548 ;
			RECT	64.193 62.484 64.225 62.548 ;
			RECT	64.361 62.484 64.393 62.548 ;
			RECT	64.529 62.484 64.561 62.548 ;
			RECT	64.697 62.484 64.729 62.548 ;
			RECT	64.865 62.484 64.897 62.548 ;
			RECT	65.033 62.484 65.065 62.548 ;
			RECT	65.201 62.484 65.233 62.548 ;
			RECT	65.369 62.484 65.401 62.548 ;
			RECT	65.537 62.484 65.569 62.548 ;
			RECT	65.705 62.484 65.737 62.548 ;
			RECT	65.873 62.484 65.905 62.548 ;
			RECT	66.041 62.484 66.073 62.548 ;
			RECT	66.209 62.484 66.241 62.548 ;
			RECT	66.377 62.484 66.409 62.548 ;
			RECT	66.545 62.484 66.577 62.548 ;
			RECT	66.713 62.484 66.745 62.548 ;
			RECT	66.881 62.484 66.913 62.548 ;
			RECT	67.049 62.484 67.081 62.548 ;
			RECT	67.217 62.484 67.249 62.548 ;
			RECT	67.385 62.484 67.417 62.548 ;
			RECT	67.553 62.484 67.585 62.548 ;
			RECT	67.721 62.484 67.753 62.548 ;
			RECT	67.889 62.484 67.921 62.548 ;
			RECT	68.057 62.484 68.089 62.548 ;
			RECT	68.225 62.484 68.257 62.548 ;
			RECT	68.393 62.484 68.425 62.548 ;
			RECT	68.561 62.484 68.593 62.548 ;
			RECT	68.729 62.484 68.761 62.548 ;
			RECT	68.897 62.484 68.929 62.548 ;
			RECT	69.065 62.484 69.097 62.548 ;
			RECT	69.233 62.484 69.265 62.548 ;
			RECT	69.401 62.484 69.433 62.548 ;
			RECT	69.569 62.484 69.601 62.548 ;
			RECT	69.737 62.484 69.769 62.548 ;
			RECT	69.905 62.484 69.937 62.548 ;
			RECT	70.073 62.484 70.105 62.548 ;
			RECT	70.241 62.484 70.273 62.548 ;
			RECT	70.409 62.484 70.441 62.548 ;
			RECT	70.577 62.484 70.609 62.548 ;
			RECT	70.745 62.484 70.777 62.548 ;
			RECT	70.913 62.484 70.945 62.548 ;
			RECT	71.081 62.484 71.113 62.548 ;
			RECT	71.249 62.484 71.281 62.548 ;
			RECT	71.417 62.484 71.449 62.548 ;
			RECT	71.585 62.484 71.617 62.548 ;
			RECT	71.753 62.484 71.785 62.548 ;
			RECT	71.921 62.484 71.953 62.548 ;
			RECT	72.089 62.484 72.121 62.548 ;
			RECT	72.257 62.484 72.289 62.548 ;
			RECT	72.425 62.484 72.457 62.548 ;
			RECT	72.593 62.484 72.625 62.548 ;
			RECT	72.761 62.484 72.793 62.548 ;
			RECT	72.929 62.484 72.961 62.548 ;
			RECT	73.097 62.484 73.129 62.548 ;
			RECT	73.265 62.484 73.297 62.548 ;
			RECT	73.433 62.484 73.465 62.548 ;
			RECT	73.601 62.484 73.633 62.548 ;
			RECT	73.769 62.484 73.801 62.548 ;
			RECT	73.937 62.484 73.969 62.548 ;
			RECT	74.105 62.484 74.137 62.548 ;
			RECT	74.273 62.484 74.305 62.548 ;
			RECT	74.441 62.484 74.473 62.548 ;
			RECT	74.609 62.484 74.641 62.548 ;
			RECT	74.777 62.484 74.809 62.548 ;
			RECT	74.945 62.484 74.977 62.548 ;
			RECT	75.113 62.484 75.145 62.548 ;
			RECT	75.281 62.484 75.313 62.548 ;
			RECT	75.449 62.484 75.481 62.548 ;
			RECT	75.617 62.484 75.649 62.548 ;
			RECT	75.785 62.484 75.817 62.548 ;
			RECT	75.953 62.484 75.985 62.548 ;
			RECT	76.121 62.484 76.153 62.548 ;
			RECT	76.289 62.484 76.321 62.548 ;
			RECT	76.457 62.484 76.489 62.548 ;
			RECT	76.625 62.484 76.657 62.548 ;
			RECT	76.793 62.484 76.825 62.548 ;
			RECT	76.961 62.484 76.993 62.548 ;
			RECT	77.129 62.484 77.161 62.548 ;
			RECT	77.297 62.484 77.329 62.548 ;
			RECT	77.465 62.484 77.497 62.548 ;
			RECT	77.633 62.484 77.665 62.548 ;
			RECT	77.801 62.484 77.833 62.548 ;
			RECT	77.969 62.484 78.001 62.548 ;
			RECT	78.137 62.484 78.169 62.548 ;
			RECT	78.305 62.484 78.337 62.548 ;
			RECT	78.473 62.484 78.505 62.548 ;
			RECT	78.641 62.484 78.673 62.548 ;
			RECT	78.809 62.484 78.841 62.548 ;
			RECT	78.977 62.484 79.009 62.548 ;
			RECT	79.145 62.484 79.177 62.548 ;
			RECT	79.313 62.484 79.345 62.548 ;
			RECT	79.481 62.484 79.513 62.548 ;
			RECT	79.649 62.484 79.681 62.548 ;
			RECT	79.817 62.484 79.849 62.548 ;
			RECT	79.985 62.484 80.017 62.548 ;
			RECT	80.153 62.484 80.185 62.548 ;
			RECT	80.321 62.484 80.353 62.548 ;
			RECT	80.489 62.484 80.521 62.548 ;
			RECT	80.657 62.484 80.689 62.548 ;
			RECT	80.825 62.484 80.857 62.548 ;
			RECT	80.993 62.484 81.025 62.548 ;
			RECT	81.161 62.484 81.193 62.548 ;
			RECT	81.329 62.484 81.361 62.548 ;
			RECT	81.497 62.484 81.529 62.548 ;
			RECT	81.665 62.484 81.697 62.548 ;
			RECT	81.833 62.484 81.865 62.548 ;
			RECT	82.001 62.484 82.033 62.548 ;
			RECT	82.169 62.484 82.201 62.548 ;
			RECT	82.337 62.484 82.369 62.548 ;
			RECT	82.505 62.484 82.537 62.548 ;
			RECT	82.673 62.484 82.705 62.548 ;
			RECT	82.841 62.484 82.873 62.548 ;
			RECT	83.009 62.484 83.041 62.548 ;
			RECT	83.177 62.484 83.209 62.548 ;
			RECT	83.345 62.484 83.377 62.548 ;
			RECT	83.513 62.484 83.545 62.548 ;
			RECT	83.681 62.484 83.713 62.548 ;
			RECT	83.849 62.484 83.881 62.548 ;
			RECT	84.017 62.484 84.049 62.548 ;
			RECT	84.185 62.484 84.217 62.548 ;
			RECT	84.353 62.484 84.385 62.548 ;
			RECT	84.521 62.484 84.553 62.548 ;
			RECT	84.689 62.484 84.721 62.548 ;
			RECT	84.857 62.484 84.889 62.548 ;
			RECT	85.025 62.484 85.057 62.548 ;
			RECT	85.193 62.484 85.225 62.548 ;
			RECT	85.361 62.484 85.393 62.548 ;
			RECT	85.529 62.484 85.561 62.548 ;
			RECT	85.697 62.484 85.729 62.548 ;
			RECT	85.865 62.484 85.897 62.548 ;
			RECT	86.033 62.484 86.065 62.548 ;
			RECT	86.201 62.484 86.233 62.548 ;
			RECT	86.369 62.484 86.401 62.548 ;
			RECT	86.537 62.484 86.569 62.548 ;
			RECT	86.705 62.484 86.737 62.548 ;
			RECT	86.873 62.484 86.905 62.548 ;
			RECT	87.041 62.484 87.073 62.548 ;
			RECT	87.209 62.484 87.241 62.548 ;
			RECT	87.377 62.484 87.409 62.548 ;
			RECT	87.545 62.484 87.577 62.548 ;
			RECT	87.713 62.484 87.745 62.548 ;
			RECT	87.881 62.484 87.913 62.548 ;
			RECT	88.049 62.484 88.081 62.548 ;
			RECT	88.217 62.484 88.249 62.548 ;
			RECT	88.385 62.484 88.417 62.548 ;
			RECT	88.553 62.484 88.585 62.548 ;
			RECT	88.721 62.484 88.753 62.548 ;
			RECT	88.889 62.484 88.921 62.548 ;
			RECT	89.057 62.484 89.089 62.548 ;
			RECT	89.225 62.484 89.257 62.548 ;
			RECT	89.393 62.484 89.425 62.548 ;
			RECT	89.561 62.484 89.593 62.548 ;
			RECT	89.729 62.484 89.761 62.548 ;
			RECT	89.897 62.484 89.929 62.548 ;
			RECT	90.065 62.484 90.097 62.548 ;
			RECT	90.233 62.484 90.265 62.548 ;
			RECT	90.401 62.484 90.433 62.548 ;
			RECT	90.569 62.484 90.601 62.548 ;
			RECT	90.737 62.484 90.769 62.548 ;
			RECT	90.905 62.484 90.937 62.548 ;
			RECT	91.073 62.484 91.105 62.548 ;
			RECT	91.241 62.484 91.273 62.548 ;
			RECT	91.409 62.484 91.441 62.548 ;
			RECT	91.577 62.484 91.609 62.548 ;
			RECT	91.745 62.484 91.777 62.548 ;
			RECT	91.913 62.484 91.945 62.548 ;
			RECT	92.081 62.484 92.113 62.548 ;
			RECT	92.249 62.484 92.281 62.548 ;
			RECT	92.417 62.484 92.449 62.548 ;
			RECT	92.585 62.484 92.617 62.548 ;
			RECT	92.753 62.484 92.785 62.548 ;
			RECT	92.921 62.484 92.953 62.548 ;
			RECT	93.089 62.484 93.121 62.548 ;
			RECT	93.257 62.484 93.289 62.548 ;
			RECT	93.425 62.484 93.457 62.548 ;
			RECT	93.593 62.484 93.625 62.548 ;
			RECT	93.761 62.484 93.793 62.548 ;
			RECT	93.929 62.484 93.961 62.548 ;
			RECT	94.097 62.484 94.129 62.548 ;
			RECT	94.265 62.484 94.297 62.548 ;
			RECT	94.433 62.484 94.465 62.548 ;
			RECT	94.601 62.484 94.633 62.548 ;
			RECT	94.769 62.484 94.801 62.548 ;
			RECT	94.937 62.484 94.969 62.548 ;
			RECT	95.105 62.484 95.137 62.548 ;
			RECT	95.273 62.484 95.305 62.548 ;
			RECT	95.441 62.484 95.473 62.548 ;
			RECT	95.609 62.484 95.641 62.548 ;
			RECT	95.777 62.484 95.809 62.548 ;
			RECT	95.945 62.484 95.977 62.548 ;
			RECT	96.113 62.484 96.145 62.548 ;
			RECT	96.281 62.484 96.313 62.548 ;
			RECT	96.449 62.484 96.481 62.548 ;
			RECT	96.617 62.484 96.649 62.548 ;
			RECT	96.785 62.484 96.817 62.548 ;
			RECT	96.953 62.484 96.985 62.548 ;
			RECT	97.121 62.484 97.153 62.548 ;
			RECT	97.289 62.484 97.321 62.548 ;
			RECT	97.457 62.484 97.489 62.548 ;
			RECT	97.625 62.484 97.657 62.548 ;
			RECT	97.793 62.484 97.825 62.548 ;
			RECT	97.961 62.484 97.993 62.548 ;
			RECT	98.129 62.484 98.161 62.548 ;
			RECT	98.297 62.484 98.329 62.548 ;
			RECT	98.465 62.484 98.497 62.548 ;
			RECT	98.633 62.484 98.665 62.548 ;
			RECT	98.801 62.484 98.833 62.548 ;
			RECT	98.969 62.484 99.001 62.548 ;
			RECT	99.137 62.484 99.169 62.548 ;
			RECT	99.305 62.484 99.337 62.548 ;
			RECT	99.473 62.484 99.505 62.548 ;
			RECT	99.641 62.484 99.673 62.548 ;
			RECT	99.809 62.484 99.841 62.548 ;
			RECT	99.977 62.484 100.009 62.548 ;
			RECT	100.145 62.484 100.177 62.548 ;
			RECT	100.313 62.484 100.345 62.548 ;
			RECT	100.481 62.484 100.513 62.548 ;
			RECT	100.649 62.484 100.681 62.548 ;
			RECT	100.817 62.484 100.849 62.548 ;
			RECT	100.985 62.484 101.017 62.548 ;
			RECT	101.153 62.484 101.185 62.548 ;
			RECT	101.321 62.484 101.353 62.548 ;
			RECT	101.489 62.484 101.521 62.548 ;
			RECT	101.657 62.484 101.689 62.548 ;
			RECT	101.825 62.484 101.857 62.548 ;
			RECT	101.993 62.484 102.025 62.548 ;
			RECT	102.123 62.5 102.155 62.532 ;
			RECT	102.245 62.495 102.277 62.527 ;
			RECT	102.375 62.484 102.407 62.548 ;
			RECT	103.795 62.484 103.827 62.548 ;
			RECT	103.925 62.495 103.957 62.527 ;
			RECT	104.047 62.5 104.079 62.532 ;
			RECT	104.177 62.484 104.209 62.548 ;
			RECT	104.345 62.484 104.377 62.548 ;
			RECT	104.513 62.484 104.545 62.548 ;
			RECT	104.681 62.484 104.713 62.548 ;
			RECT	104.849 62.484 104.881 62.548 ;
			RECT	105.017 62.484 105.049 62.548 ;
			RECT	105.185 62.484 105.217 62.548 ;
			RECT	105.353 62.484 105.385 62.548 ;
			RECT	105.521 62.484 105.553 62.548 ;
			RECT	105.689 62.484 105.721 62.548 ;
			RECT	105.857 62.484 105.889 62.548 ;
			RECT	106.025 62.484 106.057 62.548 ;
			RECT	106.193 62.484 106.225 62.548 ;
			RECT	106.361 62.484 106.393 62.548 ;
			RECT	106.529 62.484 106.561 62.548 ;
			RECT	106.697 62.484 106.729 62.548 ;
			RECT	106.865 62.484 106.897 62.548 ;
			RECT	107.033 62.484 107.065 62.548 ;
			RECT	107.201 62.484 107.233 62.548 ;
			RECT	107.369 62.484 107.401 62.548 ;
			RECT	107.537 62.484 107.569 62.548 ;
			RECT	107.705 62.484 107.737 62.548 ;
			RECT	107.873 62.484 107.905 62.548 ;
			RECT	108.041 62.484 108.073 62.548 ;
			RECT	108.209 62.484 108.241 62.548 ;
			RECT	108.377 62.484 108.409 62.548 ;
			RECT	108.545 62.484 108.577 62.548 ;
			RECT	108.713 62.484 108.745 62.548 ;
			RECT	108.881 62.484 108.913 62.548 ;
			RECT	109.049 62.484 109.081 62.548 ;
			RECT	109.217 62.484 109.249 62.548 ;
			RECT	109.385 62.484 109.417 62.548 ;
			RECT	109.553 62.484 109.585 62.548 ;
			RECT	109.721 62.484 109.753 62.548 ;
			RECT	109.889 62.484 109.921 62.548 ;
			RECT	110.057 62.484 110.089 62.548 ;
			RECT	110.225 62.484 110.257 62.548 ;
			RECT	110.393 62.484 110.425 62.548 ;
			RECT	110.561 62.484 110.593 62.548 ;
			RECT	110.729 62.484 110.761 62.548 ;
			RECT	110.897 62.484 110.929 62.548 ;
			RECT	111.065 62.484 111.097 62.548 ;
			RECT	111.233 62.484 111.265 62.548 ;
			RECT	111.401 62.484 111.433 62.548 ;
			RECT	111.569 62.484 111.601 62.548 ;
			RECT	111.737 62.484 111.769 62.548 ;
			RECT	111.905 62.484 111.937 62.548 ;
			RECT	112.073 62.484 112.105 62.548 ;
			RECT	112.241 62.484 112.273 62.548 ;
			RECT	112.409 62.484 112.441 62.548 ;
			RECT	112.577 62.484 112.609 62.548 ;
			RECT	112.745 62.484 112.777 62.548 ;
			RECT	112.913 62.484 112.945 62.548 ;
			RECT	113.081 62.484 113.113 62.548 ;
			RECT	113.249 62.484 113.281 62.548 ;
			RECT	113.417 62.484 113.449 62.548 ;
			RECT	113.585 62.484 113.617 62.548 ;
			RECT	113.753 62.484 113.785 62.548 ;
			RECT	113.921 62.484 113.953 62.548 ;
			RECT	114.089 62.484 114.121 62.548 ;
			RECT	114.257 62.484 114.289 62.548 ;
			RECT	114.425 62.484 114.457 62.548 ;
			RECT	114.593 62.484 114.625 62.548 ;
			RECT	114.761 62.484 114.793 62.548 ;
			RECT	114.929 62.484 114.961 62.548 ;
			RECT	115.097 62.484 115.129 62.548 ;
			RECT	115.265 62.484 115.297 62.548 ;
			RECT	115.433 62.484 115.465 62.548 ;
			RECT	115.601 62.484 115.633 62.548 ;
			RECT	115.769 62.484 115.801 62.548 ;
			RECT	115.937 62.484 115.969 62.548 ;
			RECT	116.105 62.484 116.137 62.548 ;
			RECT	116.273 62.484 116.305 62.548 ;
			RECT	116.441 62.484 116.473 62.548 ;
			RECT	116.609 62.484 116.641 62.548 ;
			RECT	116.777 62.484 116.809 62.548 ;
			RECT	116.945 62.484 116.977 62.548 ;
			RECT	117.113 62.484 117.145 62.548 ;
			RECT	117.281 62.484 117.313 62.548 ;
			RECT	117.449 62.484 117.481 62.548 ;
			RECT	117.617 62.484 117.649 62.548 ;
			RECT	117.785 62.484 117.817 62.548 ;
			RECT	117.953 62.484 117.985 62.548 ;
			RECT	118.121 62.484 118.153 62.548 ;
			RECT	118.289 62.484 118.321 62.548 ;
			RECT	118.457 62.484 118.489 62.548 ;
			RECT	118.625 62.484 118.657 62.548 ;
			RECT	118.793 62.484 118.825 62.548 ;
			RECT	118.961 62.484 118.993 62.548 ;
			RECT	119.129 62.484 119.161 62.548 ;
			RECT	119.297 62.484 119.329 62.548 ;
			RECT	119.465 62.484 119.497 62.548 ;
			RECT	119.633 62.484 119.665 62.548 ;
			RECT	119.801 62.484 119.833 62.548 ;
			RECT	119.969 62.484 120.001 62.548 ;
			RECT	120.137 62.484 120.169 62.548 ;
			RECT	120.305 62.484 120.337 62.548 ;
			RECT	120.473 62.484 120.505 62.548 ;
			RECT	120.641 62.484 120.673 62.548 ;
			RECT	120.809 62.484 120.841 62.548 ;
			RECT	120.977 62.484 121.009 62.548 ;
			RECT	121.145 62.484 121.177 62.548 ;
			RECT	121.313 62.484 121.345 62.548 ;
			RECT	121.481 62.484 121.513 62.548 ;
			RECT	121.649 62.484 121.681 62.548 ;
			RECT	121.817 62.484 121.849 62.548 ;
			RECT	121.985 62.484 122.017 62.548 ;
			RECT	122.153 62.484 122.185 62.548 ;
			RECT	122.321 62.484 122.353 62.548 ;
			RECT	122.489 62.484 122.521 62.548 ;
			RECT	122.657 62.484 122.689 62.548 ;
			RECT	122.825 62.484 122.857 62.548 ;
			RECT	122.993 62.484 123.025 62.548 ;
			RECT	123.161 62.484 123.193 62.548 ;
			RECT	123.329 62.484 123.361 62.548 ;
			RECT	123.497 62.484 123.529 62.548 ;
			RECT	123.665 62.484 123.697 62.548 ;
			RECT	123.833 62.484 123.865 62.548 ;
			RECT	124.001 62.484 124.033 62.548 ;
			RECT	124.169 62.484 124.201 62.548 ;
			RECT	124.337 62.484 124.369 62.548 ;
			RECT	124.505 62.484 124.537 62.548 ;
			RECT	124.673 62.484 124.705 62.548 ;
			RECT	124.841 62.484 124.873 62.548 ;
			RECT	125.009 62.484 125.041 62.548 ;
			RECT	125.177 62.484 125.209 62.548 ;
			RECT	125.345 62.484 125.377 62.548 ;
			RECT	125.513 62.484 125.545 62.548 ;
			RECT	125.681 62.484 125.713 62.548 ;
			RECT	125.849 62.484 125.881 62.548 ;
			RECT	126.017 62.484 126.049 62.548 ;
			RECT	126.185 62.484 126.217 62.548 ;
			RECT	126.353 62.484 126.385 62.548 ;
			RECT	126.521 62.484 126.553 62.548 ;
			RECT	126.689 62.484 126.721 62.548 ;
			RECT	126.857 62.484 126.889 62.548 ;
			RECT	127.025 62.484 127.057 62.548 ;
			RECT	127.193 62.484 127.225 62.548 ;
			RECT	127.361 62.484 127.393 62.548 ;
			RECT	127.529 62.484 127.561 62.548 ;
			RECT	127.697 62.484 127.729 62.548 ;
			RECT	127.865 62.484 127.897 62.548 ;
			RECT	128.033 62.484 128.065 62.548 ;
			RECT	128.201 62.484 128.233 62.548 ;
			RECT	128.369 62.484 128.401 62.548 ;
			RECT	128.537 62.484 128.569 62.548 ;
			RECT	128.705 62.484 128.737 62.548 ;
			RECT	128.873 62.484 128.905 62.548 ;
			RECT	129.041 62.484 129.073 62.548 ;
			RECT	129.209 62.484 129.241 62.548 ;
			RECT	129.377 62.484 129.409 62.548 ;
			RECT	129.545 62.484 129.577 62.548 ;
			RECT	129.713 62.484 129.745 62.548 ;
			RECT	129.881 62.484 129.913 62.548 ;
			RECT	130.049 62.484 130.081 62.548 ;
			RECT	130.217 62.484 130.249 62.548 ;
			RECT	130.385 62.484 130.417 62.548 ;
			RECT	130.553 62.484 130.585 62.548 ;
			RECT	130.721 62.484 130.753 62.548 ;
			RECT	130.889 62.484 130.921 62.548 ;
			RECT	131.057 62.484 131.089 62.548 ;
			RECT	131.225 62.484 131.257 62.548 ;
			RECT	131.393 62.484 131.425 62.548 ;
			RECT	131.561 62.484 131.593 62.548 ;
			RECT	131.729 62.484 131.761 62.548 ;
			RECT	131.897 62.484 131.929 62.548 ;
			RECT	132.065 62.484 132.097 62.548 ;
			RECT	132.233 62.484 132.265 62.548 ;
			RECT	132.401 62.484 132.433 62.548 ;
			RECT	132.569 62.484 132.601 62.548 ;
			RECT	132.737 62.484 132.769 62.548 ;
			RECT	132.905 62.484 132.937 62.548 ;
			RECT	133.073 62.484 133.105 62.548 ;
			RECT	133.241 62.484 133.273 62.548 ;
			RECT	133.409 62.484 133.441 62.548 ;
			RECT	133.577 62.484 133.609 62.548 ;
			RECT	133.745 62.484 133.777 62.548 ;
			RECT	133.913 62.484 133.945 62.548 ;
			RECT	134.081 62.484 134.113 62.548 ;
			RECT	134.249 62.484 134.281 62.548 ;
			RECT	134.417 62.484 134.449 62.548 ;
			RECT	134.585 62.484 134.617 62.548 ;
			RECT	134.753 62.484 134.785 62.548 ;
			RECT	134.921 62.484 134.953 62.548 ;
			RECT	135.089 62.484 135.121 62.548 ;
			RECT	135.257 62.484 135.289 62.548 ;
			RECT	135.425 62.484 135.457 62.548 ;
			RECT	135.593 62.484 135.625 62.548 ;
			RECT	135.761 62.484 135.793 62.548 ;
			RECT	135.929 62.484 135.961 62.548 ;
			RECT	136.097 62.484 136.129 62.548 ;
			RECT	136.265 62.484 136.297 62.548 ;
			RECT	136.433 62.484 136.465 62.548 ;
			RECT	136.601 62.484 136.633 62.548 ;
			RECT	136.769 62.484 136.801 62.548 ;
			RECT	136.937 62.484 136.969 62.548 ;
			RECT	137.105 62.484 137.137 62.548 ;
			RECT	137.273 62.484 137.305 62.548 ;
			RECT	137.441 62.484 137.473 62.548 ;
			RECT	137.609 62.484 137.641 62.548 ;
			RECT	137.777 62.484 137.809 62.548 ;
			RECT	137.945 62.484 137.977 62.548 ;
			RECT	138.113 62.484 138.145 62.548 ;
			RECT	138.281 62.484 138.313 62.548 ;
			RECT	138.449 62.484 138.481 62.548 ;
			RECT	138.617 62.484 138.649 62.548 ;
			RECT	138.785 62.484 138.817 62.548 ;
			RECT	138.953 62.484 138.985 62.548 ;
			RECT	139.121 62.484 139.153 62.548 ;
			RECT	139.289 62.484 139.321 62.548 ;
			RECT	139.457 62.484 139.489 62.548 ;
			RECT	139.625 62.484 139.657 62.548 ;
			RECT	139.793 62.484 139.825 62.548 ;
			RECT	139.961 62.484 139.993 62.548 ;
			RECT	140.129 62.484 140.161 62.548 ;
			RECT	140.297 62.484 140.329 62.548 ;
			RECT	140.465 62.484 140.497 62.548 ;
			RECT	140.633 62.484 140.665 62.548 ;
			RECT	140.801 62.484 140.833 62.548 ;
			RECT	140.969 62.484 141.001 62.548 ;
			RECT	141.137 62.484 141.169 62.548 ;
			RECT	141.305 62.484 141.337 62.548 ;
			RECT	141.473 62.484 141.505 62.548 ;
			RECT	141.641 62.484 141.673 62.548 ;
			RECT	141.809 62.484 141.841 62.548 ;
			RECT	141.977 62.484 142.009 62.548 ;
			RECT	142.145 62.484 142.177 62.548 ;
			RECT	142.313 62.484 142.345 62.548 ;
			RECT	142.481 62.484 142.513 62.548 ;
			RECT	142.649 62.484 142.681 62.548 ;
			RECT	142.817 62.484 142.849 62.548 ;
			RECT	142.985 62.484 143.017 62.548 ;
			RECT	143.153 62.484 143.185 62.548 ;
			RECT	143.321 62.484 143.353 62.548 ;
			RECT	143.489 62.484 143.521 62.548 ;
			RECT	143.657 62.484 143.689 62.548 ;
			RECT	143.825 62.484 143.857 62.548 ;
			RECT	143.993 62.484 144.025 62.548 ;
			RECT	144.161 62.484 144.193 62.548 ;
			RECT	144.329 62.484 144.361 62.548 ;
			RECT	144.497 62.484 144.529 62.548 ;
			RECT	144.665 62.484 144.697 62.548 ;
			RECT	144.833 62.484 144.865 62.548 ;
			RECT	145.001 62.484 145.033 62.548 ;
			RECT	145.169 62.484 145.201 62.548 ;
			RECT	145.337 62.484 145.369 62.548 ;
			RECT	145.505 62.484 145.537 62.548 ;
			RECT	145.673 62.484 145.705 62.548 ;
			RECT	145.841 62.484 145.873 62.548 ;
			RECT	146.009 62.484 146.041 62.548 ;
			RECT	146.177 62.484 146.209 62.548 ;
			RECT	146.345 62.484 146.377 62.548 ;
			RECT	146.513 62.484 146.545 62.548 ;
			RECT	146.681 62.484 146.713 62.548 ;
			RECT	146.849 62.484 146.881 62.548 ;
			RECT	147.017 62.484 147.049 62.548 ;
			RECT	147.185 62.484 147.217 62.548 ;
			RECT	147.316 62.5 147.348 62.532 ;
			RECT	147.437 62.5 147.469 62.532 ;
			RECT	147.567 62.484 147.599 62.548 ;
			RECT	149.879 62.484 149.911 62.548 ;
			RECT	151.13 62.484 151.194 62.548 ;
			RECT	151.81 62.484 151.842 62.548 ;
			RECT	152.249 62.484 152.281 62.548 ;
			RECT	153.56 62.484 153.624 62.548 ;
			RECT	156.601 62.484 156.633 62.548 ;
			RECT	156.731 62.5 156.763 62.532 ;
			RECT	156.852 62.5 156.884 62.532 ;
			RECT	156.983 62.484 157.015 62.548 ;
			RECT	157.151 62.484 157.183 62.548 ;
			RECT	157.319 62.484 157.351 62.548 ;
			RECT	157.487 62.484 157.519 62.548 ;
			RECT	157.655 62.484 157.687 62.548 ;
			RECT	157.823 62.484 157.855 62.548 ;
			RECT	157.991 62.484 158.023 62.548 ;
			RECT	158.159 62.484 158.191 62.548 ;
			RECT	158.327 62.484 158.359 62.548 ;
			RECT	158.495 62.484 158.527 62.548 ;
			RECT	158.663 62.484 158.695 62.548 ;
			RECT	158.831 62.484 158.863 62.548 ;
			RECT	158.999 62.484 159.031 62.548 ;
			RECT	159.167 62.484 159.199 62.548 ;
			RECT	159.335 62.484 159.367 62.548 ;
			RECT	159.503 62.484 159.535 62.548 ;
			RECT	159.671 62.484 159.703 62.548 ;
			RECT	159.839 62.484 159.871 62.548 ;
			RECT	160.007 62.484 160.039 62.548 ;
			RECT	160.175 62.484 160.207 62.548 ;
			RECT	160.343 62.484 160.375 62.548 ;
			RECT	160.511 62.484 160.543 62.548 ;
			RECT	160.679 62.484 160.711 62.548 ;
			RECT	160.847 62.484 160.879 62.548 ;
			RECT	161.015 62.484 161.047 62.548 ;
			RECT	161.183 62.484 161.215 62.548 ;
			RECT	161.351 62.484 161.383 62.548 ;
			RECT	161.519 62.484 161.551 62.548 ;
			RECT	161.687 62.484 161.719 62.548 ;
			RECT	161.855 62.484 161.887 62.548 ;
			RECT	162.023 62.484 162.055 62.548 ;
			RECT	162.191 62.484 162.223 62.548 ;
			RECT	162.359 62.484 162.391 62.548 ;
			RECT	162.527 62.484 162.559 62.548 ;
			RECT	162.695 62.484 162.727 62.548 ;
			RECT	162.863 62.484 162.895 62.548 ;
			RECT	163.031 62.484 163.063 62.548 ;
			RECT	163.199 62.484 163.231 62.548 ;
			RECT	163.367 62.484 163.399 62.548 ;
			RECT	163.535 62.484 163.567 62.548 ;
			RECT	163.703 62.484 163.735 62.548 ;
			RECT	163.871 62.484 163.903 62.548 ;
			RECT	164.039 62.484 164.071 62.548 ;
			RECT	164.207 62.484 164.239 62.548 ;
			RECT	164.375 62.484 164.407 62.548 ;
			RECT	164.543 62.484 164.575 62.548 ;
			RECT	164.711 62.484 164.743 62.548 ;
			RECT	164.879 62.484 164.911 62.548 ;
			RECT	165.047 62.484 165.079 62.548 ;
			RECT	165.215 62.484 165.247 62.548 ;
			RECT	165.383 62.484 165.415 62.548 ;
			RECT	165.551 62.484 165.583 62.548 ;
			RECT	165.719 62.484 165.751 62.548 ;
			RECT	165.887 62.484 165.919 62.548 ;
			RECT	166.055 62.484 166.087 62.548 ;
			RECT	166.223 62.484 166.255 62.548 ;
			RECT	166.391 62.484 166.423 62.548 ;
			RECT	166.559 62.484 166.591 62.548 ;
			RECT	166.727 62.484 166.759 62.548 ;
			RECT	166.895 62.484 166.927 62.548 ;
			RECT	167.063 62.484 167.095 62.548 ;
			RECT	167.231 62.484 167.263 62.548 ;
			RECT	167.399 62.484 167.431 62.548 ;
			RECT	167.567 62.484 167.599 62.548 ;
			RECT	167.735 62.484 167.767 62.548 ;
			RECT	167.903 62.484 167.935 62.548 ;
			RECT	168.071 62.484 168.103 62.548 ;
			RECT	168.239 62.484 168.271 62.548 ;
			RECT	168.407 62.484 168.439 62.548 ;
			RECT	168.575 62.484 168.607 62.548 ;
			RECT	168.743 62.484 168.775 62.548 ;
			RECT	168.911 62.484 168.943 62.548 ;
			RECT	169.079 62.484 169.111 62.548 ;
			RECT	169.247 62.484 169.279 62.548 ;
			RECT	169.415 62.484 169.447 62.548 ;
			RECT	169.583 62.484 169.615 62.548 ;
			RECT	169.751 62.484 169.783 62.548 ;
			RECT	169.919 62.484 169.951 62.548 ;
			RECT	170.087 62.484 170.119 62.548 ;
			RECT	170.255 62.484 170.287 62.548 ;
			RECT	170.423 62.484 170.455 62.548 ;
			RECT	170.591 62.484 170.623 62.548 ;
			RECT	170.759 62.484 170.791 62.548 ;
			RECT	170.927 62.484 170.959 62.548 ;
			RECT	171.095 62.484 171.127 62.548 ;
			RECT	171.263 62.484 171.295 62.548 ;
			RECT	171.431 62.484 171.463 62.548 ;
			RECT	171.599 62.484 171.631 62.548 ;
			RECT	171.767 62.484 171.799 62.548 ;
			RECT	171.935 62.484 171.967 62.548 ;
			RECT	172.103 62.484 172.135 62.548 ;
			RECT	172.271 62.484 172.303 62.548 ;
			RECT	172.439 62.484 172.471 62.548 ;
			RECT	172.607 62.484 172.639 62.548 ;
			RECT	172.775 62.484 172.807 62.548 ;
			RECT	172.943 62.484 172.975 62.548 ;
			RECT	173.111 62.484 173.143 62.548 ;
			RECT	173.279 62.484 173.311 62.548 ;
			RECT	173.447 62.484 173.479 62.548 ;
			RECT	173.615 62.484 173.647 62.548 ;
			RECT	173.783 62.484 173.815 62.548 ;
			RECT	173.951 62.484 173.983 62.548 ;
			RECT	174.119 62.484 174.151 62.548 ;
			RECT	174.287 62.484 174.319 62.548 ;
			RECT	174.455 62.484 174.487 62.548 ;
			RECT	174.623 62.484 174.655 62.548 ;
			RECT	174.791 62.484 174.823 62.548 ;
			RECT	174.959 62.484 174.991 62.548 ;
			RECT	175.127 62.484 175.159 62.548 ;
			RECT	175.295 62.484 175.327 62.548 ;
			RECT	175.463 62.484 175.495 62.548 ;
			RECT	175.631 62.484 175.663 62.548 ;
			RECT	175.799 62.484 175.831 62.548 ;
			RECT	175.967 62.484 175.999 62.548 ;
			RECT	176.135 62.484 176.167 62.548 ;
			RECT	176.303 62.484 176.335 62.548 ;
			RECT	176.471 62.484 176.503 62.548 ;
			RECT	176.639 62.484 176.671 62.548 ;
			RECT	176.807 62.484 176.839 62.548 ;
			RECT	176.975 62.484 177.007 62.548 ;
			RECT	177.143 62.484 177.175 62.548 ;
			RECT	177.311 62.484 177.343 62.548 ;
			RECT	177.479 62.484 177.511 62.548 ;
			RECT	177.647 62.484 177.679 62.548 ;
			RECT	177.815 62.484 177.847 62.548 ;
			RECT	177.983 62.484 178.015 62.548 ;
			RECT	178.151 62.484 178.183 62.548 ;
			RECT	178.319 62.484 178.351 62.548 ;
			RECT	178.487 62.484 178.519 62.548 ;
			RECT	178.655 62.484 178.687 62.548 ;
			RECT	178.823 62.484 178.855 62.548 ;
			RECT	178.991 62.484 179.023 62.548 ;
			RECT	179.159 62.484 179.191 62.548 ;
			RECT	179.327 62.484 179.359 62.548 ;
			RECT	179.495 62.484 179.527 62.548 ;
			RECT	179.663 62.484 179.695 62.548 ;
			RECT	179.831 62.484 179.863 62.548 ;
			RECT	179.999 62.484 180.031 62.548 ;
			RECT	180.167 62.484 180.199 62.548 ;
			RECT	180.335 62.484 180.367 62.548 ;
			RECT	180.503 62.484 180.535 62.548 ;
			RECT	180.671 62.484 180.703 62.548 ;
			RECT	180.839 62.484 180.871 62.548 ;
			RECT	181.007 62.484 181.039 62.548 ;
			RECT	181.175 62.484 181.207 62.548 ;
			RECT	181.343 62.484 181.375 62.548 ;
			RECT	181.511 62.484 181.543 62.548 ;
			RECT	181.679 62.484 181.711 62.548 ;
			RECT	181.847 62.484 181.879 62.548 ;
			RECT	182.015 62.484 182.047 62.548 ;
			RECT	182.183 62.484 182.215 62.548 ;
			RECT	182.351 62.484 182.383 62.548 ;
			RECT	182.519 62.484 182.551 62.548 ;
			RECT	182.687 62.484 182.719 62.548 ;
			RECT	182.855 62.484 182.887 62.548 ;
			RECT	183.023 62.484 183.055 62.548 ;
			RECT	183.191 62.484 183.223 62.548 ;
			RECT	183.359 62.484 183.391 62.548 ;
			RECT	183.527 62.484 183.559 62.548 ;
			RECT	183.695 62.484 183.727 62.548 ;
			RECT	183.863 62.484 183.895 62.548 ;
			RECT	184.031 62.484 184.063 62.548 ;
			RECT	184.199 62.484 184.231 62.548 ;
			RECT	184.367 62.484 184.399 62.548 ;
			RECT	184.535 62.484 184.567 62.548 ;
			RECT	184.703 62.484 184.735 62.548 ;
			RECT	184.871 62.484 184.903 62.548 ;
			RECT	185.039 62.484 185.071 62.548 ;
			RECT	185.207 62.484 185.239 62.548 ;
			RECT	185.375 62.484 185.407 62.548 ;
			RECT	185.543 62.484 185.575 62.548 ;
			RECT	185.711 62.484 185.743 62.548 ;
			RECT	185.879 62.484 185.911 62.548 ;
			RECT	186.047 62.484 186.079 62.548 ;
			RECT	186.215 62.484 186.247 62.548 ;
			RECT	186.383 62.484 186.415 62.548 ;
			RECT	186.551 62.484 186.583 62.548 ;
			RECT	186.719 62.484 186.751 62.548 ;
			RECT	186.887 62.484 186.919 62.548 ;
			RECT	187.055 62.484 187.087 62.548 ;
			RECT	187.223 62.484 187.255 62.548 ;
			RECT	187.391 62.484 187.423 62.548 ;
			RECT	187.559 62.484 187.591 62.548 ;
			RECT	187.727 62.484 187.759 62.548 ;
			RECT	187.895 62.484 187.927 62.548 ;
			RECT	188.063 62.484 188.095 62.548 ;
			RECT	188.231 62.484 188.263 62.548 ;
			RECT	188.399 62.484 188.431 62.548 ;
			RECT	188.567 62.484 188.599 62.548 ;
			RECT	188.735 62.484 188.767 62.548 ;
			RECT	188.903 62.484 188.935 62.548 ;
			RECT	189.071 62.484 189.103 62.548 ;
			RECT	189.239 62.484 189.271 62.548 ;
			RECT	189.407 62.484 189.439 62.548 ;
			RECT	189.575 62.484 189.607 62.548 ;
			RECT	189.743 62.484 189.775 62.548 ;
			RECT	189.911 62.484 189.943 62.548 ;
			RECT	190.079 62.484 190.111 62.548 ;
			RECT	190.247 62.484 190.279 62.548 ;
			RECT	190.415 62.484 190.447 62.548 ;
			RECT	190.583 62.484 190.615 62.548 ;
			RECT	190.751 62.484 190.783 62.548 ;
			RECT	190.919 62.484 190.951 62.548 ;
			RECT	191.087 62.484 191.119 62.548 ;
			RECT	191.255 62.484 191.287 62.548 ;
			RECT	191.423 62.484 191.455 62.548 ;
			RECT	191.591 62.484 191.623 62.548 ;
			RECT	191.759 62.484 191.791 62.548 ;
			RECT	191.927 62.484 191.959 62.548 ;
			RECT	192.095 62.484 192.127 62.548 ;
			RECT	192.263 62.484 192.295 62.548 ;
			RECT	192.431 62.484 192.463 62.548 ;
			RECT	192.599 62.484 192.631 62.548 ;
			RECT	192.767 62.484 192.799 62.548 ;
			RECT	192.935 62.484 192.967 62.548 ;
			RECT	193.103 62.484 193.135 62.548 ;
			RECT	193.271 62.484 193.303 62.548 ;
			RECT	193.439 62.484 193.471 62.548 ;
			RECT	193.607 62.484 193.639 62.548 ;
			RECT	193.775 62.484 193.807 62.548 ;
			RECT	193.943 62.484 193.975 62.548 ;
			RECT	194.111 62.484 194.143 62.548 ;
			RECT	194.279 62.484 194.311 62.548 ;
			RECT	194.447 62.484 194.479 62.548 ;
			RECT	194.615 62.484 194.647 62.548 ;
			RECT	194.783 62.484 194.815 62.548 ;
			RECT	194.951 62.484 194.983 62.548 ;
			RECT	195.119 62.484 195.151 62.548 ;
			RECT	195.287 62.484 195.319 62.548 ;
			RECT	195.455 62.484 195.487 62.548 ;
			RECT	195.623 62.484 195.655 62.548 ;
			RECT	195.791 62.484 195.823 62.548 ;
			RECT	195.959 62.484 195.991 62.548 ;
			RECT	196.127 62.484 196.159 62.548 ;
			RECT	196.295 62.484 196.327 62.548 ;
			RECT	196.463 62.484 196.495 62.548 ;
			RECT	196.631 62.484 196.663 62.548 ;
			RECT	196.799 62.484 196.831 62.548 ;
			RECT	196.967 62.484 196.999 62.548 ;
			RECT	197.135 62.484 197.167 62.548 ;
			RECT	197.303 62.484 197.335 62.548 ;
			RECT	197.471 62.484 197.503 62.548 ;
			RECT	197.639 62.484 197.671 62.548 ;
			RECT	197.807 62.484 197.839 62.548 ;
			RECT	197.975 62.484 198.007 62.548 ;
			RECT	198.143 62.484 198.175 62.548 ;
			RECT	198.311 62.484 198.343 62.548 ;
			RECT	198.479 62.484 198.511 62.548 ;
			RECT	198.647 62.484 198.679 62.548 ;
			RECT	198.815 62.484 198.847 62.548 ;
			RECT	198.983 62.484 199.015 62.548 ;
			RECT	199.151 62.484 199.183 62.548 ;
			RECT	199.319 62.484 199.351 62.548 ;
			RECT	199.487 62.484 199.519 62.548 ;
			RECT	199.655 62.484 199.687 62.548 ;
			RECT	199.823 62.484 199.855 62.548 ;
			RECT	199.991 62.484 200.023 62.548 ;
			RECT	200.121 62.5 200.153 62.532 ;
			RECT	200.243 62.495 200.275 62.527 ;
			RECT	200.373 62.484 200.405 62.548 ;
			RECT	200.9 62.484 200.932 62.548 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 60.536 201.665 60.656 ;
			LAYER	J3 ;
			RECT	0.755 60.564 0.787 60.628 ;
			RECT	1.645 60.564 1.709 60.628 ;
			RECT	2.323 60.564 2.387 60.628 ;
			RECT	3.438 60.564 3.47 60.628 ;
			RECT	3.585 60.564 3.617 60.628 ;
			RECT	4.195 60.564 4.227 60.628 ;
			RECT	4.72 60.564 4.752 60.628 ;
			RECT	4.944 60.564 5.008 60.628 ;
			RECT	5.267 60.564 5.299 60.628 ;
			RECT	5.797 60.564 5.829 60.628 ;
			RECT	5.927 60.575 5.959 60.607 ;
			RECT	6.049 60.58 6.081 60.612 ;
			RECT	6.179 60.564 6.211 60.628 ;
			RECT	6.347 60.564 6.379 60.628 ;
			RECT	6.515 60.564 6.547 60.628 ;
			RECT	6.683 60.564 6.715 60.628 ;
			RECT	6.851 60.564 6.883 60.628 ;
			RECT	7.019 60.564 7.051 60.628 ;
			RECT	7.187 60.564 7.219 60.628 ;
			RECT	7.355 60.564 7.387 60.628 ;
			RECT	7.523 60.564 7.555 60.628 ;
			RECT	7.691 60.564 7.723 60.628 ;
			RECT	7.859 60.564 7.891 60.628 ;
			RECT	8.027 60.564 8.059 60.628 ;
			RECT	8.195 60.564 8.227 60.628 ;
			RECT	8.363 60.564 8.395 60.628 ;
			RECT	8.531 60.564 8.563 60.628 ;
			RECT	8.699 60.564 8.731 60.628 ;
			RECT	8.867 60.564 8.899 60.628 ;
			RECT	9.035 60.564 9.067 60.628 ;
			RECT	9.203 60.564 9.235 60.628 ;
			RECT	9.371 60.564 9.403 60.628 ;
			RECT	9.539 60.564 9.571 60.628 ;
			RECT	9.707 60.564 9.739 60.628 ;
			RECT	9.875 60.564 9.907 60.628 ;
			RECT	10.043 60.564 10.075 60.628 ;
			RECT	10.211 60.564 10.243 60.628 ;
			RECT	10.379 60.564 10.411 60.628 ;
			RECT	10.547 60.564 10.579 60.628 ;
			RECT	10.715 60.564 10.747 60.628 ;
			RECT	10.883 60.564 10.915 60.628 ;
			RECT	11.051 60.564 11.083 60.628 ;
			RECT	11.219 60.564 11.251 60.628 ;
			RECT	11.387 60.564 11.419 60.628 ;
			RECT	11.555 60.564 11.587 60.628 ;
			RECT	11.723 60.564 11.755 60.628 ;
			RECT	11.891 60.564 11.923 60.628 ;
			RECT	12.059 60.564 12.091 60.628 ;
			RECT	12.227 60.564 12.259 60.628 ;
			RECT	12.395 60.564 12.427 60.628 ;
			RECT	12.563 60.564 12.595 60.628 ;
			RECT	12.731 60.564 12.763 60.628 ;
			RECT	12.899 60.564 12.931 60.628 ;
			RECT	13.067 60.564 13.099 60.628 ;
			RECT	13.235 60.564 13.267 60.628 ;
			RECT	13.403 60.564 13.435 60.628 ;
			RECT	13.571 60.564 13.603 60.628 ;
			RECT	13.739 60.564 13.771 60.628 ;
			RECT	13.907 60.564 13.939 60.628 ;
			RECT	14.075 60.564 14.107 60.628 ;
			RECT	14.243 60.564 14.275 60.628 ;
			RECT	14.411 60.564 14.443 60.628 ;
			RECT	14.579 60.564 14.611 60.628 ;
			RECT	14.747 60.564 14.779 60.628 ;
			RECT	14.915 60.564 14.947 60.628 ;
			RECT	15.083 60.564 15.115 60.628 ;
			RECT	15.251 60.564 15.283 60.628 ;
			RECT	15.419 60.564 15.451 60.628 ;
			RECT	15.587 60.564 15.619 60.628 ;
			RECT	15.755 60.564 15.787 60.628 ;
			RECT	15.923 60.564 15.955 60.628 ;
			RECT	16.091 60.564 16.123 60.628 ;
			RECT	16.259 60.564 16.291 60.628 ;
			RECT	16.427 60.564 16.459 60.628 ;
			RECT	16.595 60.564 16.627 60.628 ;
			RECT	16.763 60.564 16.795 60.628 ;
			RECT	16.931 60.564 16.963 60.628 ;
			RECT	17.099 60.564 17.131 60.628 ;
			RECT	17.267 60.564 17.299 60.628 ;
			RECT	17.435 60.564 17.467 60.628 ;
			RECT	17.603 60.564 17.635 60.628 ;
			RECT	17.771 60.564 17.803 60.628 ;
			RECT	17.939 60.564 17.971 60.628 ;
			RECT	18.107 60.564 18.139 60.628 ;
			RECT	18.275 60.564 18.307 60.628 ;
			RECT	18.443 60.564 18.475 60.628 ;
			RECT	18.611 60.564 18.643 60.628 ;
			RECT	18.779 60.564 18.811 60.628 ;
			RECT	18.947 60.564 18.979 60.628 ;
			RECT	19.115 60.564 19.147 60.628 ;
			RECT	19.283 60.564 19.315 60.628 ;
			RECT	19.451 60.564 19.483 60.628 ;
			RECT	19.619 60.564 19.651 60.628 ;
			RECT	19.787 60.564 19.819 60.628 ;
			RECT	19.955 60.564 19.987 60.628 ;
			RECT	20.123 60.564 20.155 60.628 ;
			RECT	20.291 60.564 20.323 60.628 ;
			RECT	20.459 60.564 20.491 60.628 ;
			RECT	20.627 60.564 20.659 60.628 ;
			RECT	20.795 60.564 20.827 60.628 ;
			RECT	20.963 60.564 20.995 60.628 ;
			RECT	21.131 60.564 21.163 60.628 ;
			RECT	21.299 60.564 21.331 60.628 ;
			RECT	21.467 60.564 21.499 60.628 ;
			RECT	21.635 60.564 21.667 60.628 ;
			RECT	21.803 60.564 21.835 60.628 ;
			RECT	21.971 60.564 22.003 60.628 ;
			RECT	22.139 60.564 22.171 60.628 ;
			RECT	22.307 60.564 22.339 60.628 ;
			RECT	22.475 60.564 22.507 60.628 ;
			RECT	22.643 60.564 22.675 60.628 ;
			RECT	22.811 60.564 22.843 60.628 ;
			RECT	22.979 60.564 23.011 60.628 ;
			RECT	23.147 60.564 23.179 60.628 ;
			RECT	23.315 60.564 23.347 60.628 ;
			RECT	23.483 60.564 23.515 60.628 ;
			RECT	23.651 60.564 23.683 60.628 ;
			RECT	23.819 60.564 23.851 60.628 ;
			RECT	23.987 60.564 24.019 60.628 ;
			RECT	24.155 60.564 24.187 60.628 ;
			RECT	24.323 60.564 24.355 60.628 ;
			RECT	24.491 60.564 24.523 60.628 ;
			RECT	24.659 60.564 24.691 60.628 ;
			RECT	24.827 60.564 24.859 60.628 ;
			RECT	24.995 60.564 25.027 60.628 ;
			RECT	25.163 60.564 25.195 60.628 ;
			RECT	25.331 60.564 25.363 60.628 ;
			RECT	25.499 60.564 25.531 60.628 ;
			RECT	25.667 60.564 25.699 60.628 ;
			RECT	25.835 60.564 25.867 60.628 ;
			RECT	26.003 60.564 26.035 60.628 ;
			RECT	26.171 60.564 26.203 60.628 ;
			RECT	26.339 60.564 26.371 60.628 ;
			RECT	26.507 60.564 26.539 60.628 ;
			RECT	26.675 60.564 26.707 60.628 ;
			RECT	26.843 60.564 26.875 60.628 ;
			RECT	27.011 60.564 27.043 60.628 ;
			RECT	27.179 60.564 27.211 60.628 ;
			RECT	27.347 60.564 27.379 60.628 ;
			RECT	27.515 60.564 27.547 60.628 ;
			RECT	27.683 60.564 27.715 60.628 ;
			RECT	27.851 60.564 27.883 60.628 ;
			RECT	28.019 60.564 28.051 60.628 ;
			RECT	28.187 60.564 28.219 60.628 ;
			RECT	28.355 60.564 28.387 60.628 ;
			RECT	28.523 60.564 28.555 60.628 ;
			RECT	28.691 60.564 28.723 60.628 ;
			RECT	28.859 60.564 28.891 60.628 ;
			RECT	29.027 60.564 29.059 60.628 ;
			RECT	29.195 60.564 29.227 60.628 ;
			RECT	29.363 60.564 29.395 60.628 ;
			RECT	29.531 60.564 29.563 60.628 ;
			RECT	29.699 60.564 29.731 60.628 ;
			RECT	29.867 60.564 29.899 60.628 ;
			RECT	30.035 60.564 30.067 60.628 ;
			RECT	30.203 60.564 30.235 60.628 ;
			RECT	30.371 60.564 30.403 60.628 ;
			RECT	30.539 60.564 30.571 60.628 ;
			RECT	30.707 60.564 30.739 60.628 ;
			RECT	30.875 60.564 30.907 60.628 ;
			RECT	31.043 60.564 31.075 60.628 ;
			RECT	31.211 60.564 31.243 60.628 ;
			RECT	31.379 60.564 31.411 60.628 ;
			RECT	31.547 60.564 31.579 60.628 ;
			RECT	31.715 60.564 31.747 60.628 ;
			RECT	31.883 60.564 31.915 60.628 ;
			RECT	32.051 60.564 32.083 60.628 ;
			RECT	32.219 60.564 32.251 60.628 ;
			RECT	32.387 60.564 32.419 60.628 ;
			RECT	32.555 60.564 32.587 60.628 ;
			RECT	32.723 60.564 32.755 60.628 ;
			RECT	32.891 60.564 32.923 60.628 ;
			RECT	33.059 60.564 33.091 60.628 ;
			RECT	33.227 60.564 33.259 60.628 ;
			RECT	33.395 60.564 33.427 60.628 ;
			RECT	33.563 60.564 33.595 60.628 ;
			RECT	33.731 60.564 33.763 60.628 ;
			RECT	33.899 60.564 33.931 60.628 ;
			RECT	34.067 60.564 34.099 60.628 ;
			RECT	34.235 60.564 34.267 60.628 ;
			RECT	34.403 60.564 34.435 60.628 ;
			RECT	34.571 60.564 34.603 60.628 ;
			RECT	34.739 60.564 34.771 60.628 ;
			RECT	34.907 60.564 34.939 60.628 ;
			RECT	35.075 60.564 35.107 60.628 ;
			RECT	35.243 60.564 35.275 60.628 ;
			RECT	35.411 60.564 35.443 60.628 ;
			RECT	35.579 60.564 35.611 60.628 ;
			RECT	35.747 60.564 35.779 60.628 ;
			RECT	35.915 60.564 35.947 60.628 ;
			RECT	36.083 60.564 36.115 60.628 ;
			RECT	36.251 60.564 36.283 60.628 ;
			RECT	36.419 60.564 36.451 60.628 ;
			RECT	36.587 60.564 36.619 60.628 ;
			RECT	36.755 60.564 36.787 60.628 ;
			RECT	36.923 60.564 36.955 60.628 ;
			RECT	37.091 60.564 37.123 60.628 ;
			RECT	37.259 60.564 37.291 60.628 ;
			RECT	37.427 60.564 37.459 60.628 ;
			RECT	37.595 60.564 37.627 60.628 ;
			RECT	37.763 60.564 37.795 60.628 ;
			RECT	37.931 60.564 37.963 60.628 ;
			RECT	38.099 60.564 38.131 60.628 ;
			RECT	38.267 60.564 38.299 60.628 ;
			RECT	38.435 60.564 38.467 60.628 ;
			RECT	38.603 60.564 38.635 60.628 ;
			RECT	38.771 60.564 38.803 60.628 ;
			RECT	38.939 60.564 38.971 60.628 ;
			RECT	39.107 60.564 39.139 60.628 ;
			RECT	39.275 60.564 39.307 60.628 ;
			RECT	39.443 60.564 39.475 60.628 ;
			RECT	39.611 60.564 39.643 60.628 ;
			RECT	39.779 60.564 39.811 60.628 ;
			RECT	39.947 60.564 39.979 60.628 ;
			RECT	40.115 60.564 40.147 60.628 ;
			RECT	40.283 60.564 40.315 60.628 ;
			RECT	40.451 60.564 40.483 60.628 ;
			RECT	40.619 60.564 40.651 60.628 ;
			RECT	40.787 60.564 40.819 60.628 ;
			RECT	40.955 60.564 40.987 60.628 ;
			RECT	41.123 60.564 41.155 60.628 ;
			RECT	41.291 60.564 41.323 60.628 ;
			RECT	41.459 60.564 41.491 60.628 ;
			RECT	41.627 60.564 41.659 60.628 ;
			RECT	41.795 60.564 41.827 60.628 ;
			RECT	41.963 60.564 41.995 60.628 ;
			RECT	42.131 60.564 42.163 60.628 ;
			RECT	42.299 60.564 42.331 60.628 ;
			RECT	42.467 60.564 42.499 60.628 ;
			RECT	42.635 60.564 42.667 60.628 ;
			RECT	42.803 60.564 42.835 60.628 ;
			RECT	42.971 60.564 43.003 60.628 ;
			RECT	43.139 60.564 43.171 60.628 ;
			RECT	43.307 60.564 43.339 60.628 ;
			RECT	43.475 60.564 43.507 60.628 ;
			RECT	43.643 60.564 43.675 60.628 ;
			RECT	43.811 60.564 43.843 60.628 ;
			RECT	43.979 60.564 44.011 60.628 ;
			RECT	44.147 60.564 44.179 60.628 ;
			RECT	44.315 60.564 44.347 60.628 ;
			RECT	44.483 60.564 44.515 60.628 ;
			RECT	44.651 60.564 44.683 60.628 ;
			RECT	44.819 60.564 44.851 60.628 ;
			RECT	44.987 60.564 45.019 60.628 ;
			RECT	45.155 60.564 45.187 60.628 ;
			RECT	45.323 60.564 45.355 60.628 ;
			RECT	45.491 60.564 45.523 60.628 ;
			RECT	45.659 60.564 45.691 60.628 ;
			RECT	45.827 60.564 45.859 60.628 ;
			RECT	45.995 60.564 46.027 60.628 ;
			RECT	46.163 60.564 46.195 60.628 ;
			RECT	46.331 60.564 46.363 60.628 ;
			RECT	46.499 60.564 46.531 60.628 ;
			RECT	46.667 60.564 46.699 60.628 ;
			RECT	46.835 60.564 46.867 60.628 ;
			RECT	47.003 60.564 47.035 60.628 ;
			RECT	47.171 60.564 47.203 60.628 ;
			RECT	47.339 60.564 47.371 60.628 ;
			RECT	47.507 60.564 47.539 60.628 ;
			RECT	47.675 60.564 47.707 60.628 ;
			RECT	47.843 60.564 47.875 60.628 ;
			RECT	48.011 60.564 48.043 60.628 ;
			RECT	48.179 60.564 48.211 60.628 ;
			RECT	48.347 60.564 48.379 60.628 ;
			RECT	48.515 60.564 48.547 60.628 ;
			RECT	48.683 60.564 48.715 60.628 ;
			RECT	48.851 60.564 48.883 60.628 ;
			RECT	49.019 60.564 49.051 60.628 ;
			RECT	49.187 60.564 49.219 60.628 ;
			RECT	49.318 60.58 49.35 60.612 ;
			RECT	49.439 60.58 49.471 60.612 ;
			RECT	49.569 60.564 49.601 60.628 ;
			RECT	51.881 60.564 51.913 60.628 ;
			RECT	53.132 60.564 53.196 60.628 ;
			RECT	53.812 60.564 53.844 60.628 ;
			RECT	54.251 60.564 54.283 60.628 ;
			RECT	55.562 60.564 55.626 60.628 ;
			RECT	58.603 60.564 58.635 60.628 ;
			RECT	58.733 60.58 58.765 60.612 ;
			RECT	58.854 60.58 58.886 60.612 ;
			RECT	58.985 60.564 59.017 60.628 ;
			RECT	59.153 60.564 59.185 60.628 ;
			RECT	59.321 60.564 59.353 60.628 ;
			RECT	59.489 60.564 59.521 60.628 ;
			RECT	59.657 60.564 59.689 60.628 ;
			RECT	59.825 60.564 59.857 60.628 ;
			RECT	59.993 60.564 60.025 60.628 ;
			RECT	60.161 60.564 60.193 60.628 ;
			RECT	60.329 60.564 60.361 60.628 ;
			RECT	60.497 60.564 60.529 60.628 ;
			RECT	60.665 60.564 60.697 60.628 ;
			RECT	60.833 60.564 60.865 60.628 ;
			RECT	61.001 60.564 61.033 60.628 ;
			RECT	61.169 60.564 61.201 60.628 ;
			RECT	61.337 60.564 61.369 60.628 ;
			RECT	61.505 60.564 61.537 60.628 ;
			RECT	61.673 60.564 61.705 60.628 ;
			RECT	61.841 60.564 61.873 60.628 ;
			RECT	62.009 60.564 62.041 60.628 ;
			RECT	62.177 60.564 62.209 60.628 ;
			RECT	62.345 60.564 62.377 60.628 ;
			RECT	62.513 60.564 62.545 60.628 ;
			RECT	62.681 60.564 62.713 60.628 ;
			RECT	62.849 60.564 62.881 60.628 ;
			RECT	63.017 60.564 63.049 60.628 ;
			RECT	63.185 60.564 63.217 60.628 ;
			RECT	63.353 60.564 63.385 60.628 ;
			RECT	63.521 60.564 63.553 60.628 ;
			RECT	63.689 60.564 63.721 60.628 ;
			RECT	63.857 60.564 63.889 60.628 ;
			RECT	64.025 60.564 64.057 60.628 ;
			RECT	64.193 60.564 64.225 60.628 ;
			RECT	64.361 60.564 64.393 60.628 ;
			RECT	64.529 60.564 64.561 60.628 ;
			RECT	64.697 60.564 64.729 60.628 ;
			RECT	64.865 60.564 64.897 60.628 ;
			RECT	65.033 60.564 65.065 60.628 ;
			RECT	65.201 60.564 65.233 60.628 ;
			RECT	65.369 60.564 65.401 60.628 ;
			RECT	65.537 60.564 65.569 60.628 ;
			RECT	65.705 60.564 65.737 60.628 ;
			RECT	65.873 60.564 65.905 60.628 ;
			RECT	66.041 60.564 66.073 60.628 ;
			RECT	66.209 60.564 66.241 60.628 ;
			RECT	66.377 60.564 66.409 60.628 ;
			RECT	66.545 60.564 66.577 60.628 ;
			RECT	66.713 60.564 66.745 60.628 ;
			RECT	66.881 60.564 66.913 60.628 ;
			RECT	67.049 60.564 67.081 60.628 ;
			RECT	67.217 60.564 67.249 60.628 ;
			RECT	67.385 60.564 67.417 60.628 ;
			RECT	67.553 60.564 67.585 60.628 ;
			RECT	67.721 60.564 67.753 60.628 ;
			RECT	67.889 60.564 67.921 60.628 ;
			RECT	68.057 60.564 68.089 60.628 ;
			RECT	68.225 60.564 68.257 60.628 ;
			RECT	68.393 60.564 68.425 60.628 ;
			RECT	68.561 60.564 68.593 60.628 ;
			RECT	68.729 60.564 68.761 60.628 ;
			RECT	68.897 60.564 68.929 60.628 ;
			RECT	69.065 60.564 69.097 60.628 ;
			RECT	69.233 60.564 69.265 60.628 ;
			RECT	69.401 60.564 69.433 60.628 ;
			RECT	69.569 60.564 69.601 60.628 ;
			RECT	69.737 60.564 69.769 60.628 ;
			RECT	69.905 60.564 69.937 60.628 ;
			RECT	70.073 60.564 70.105 60.628 ;
			RECT	70.241 60.564 70.273 60.628 ;
			RECT	70.409 60.564 70.441 60.628 ;
			RECT	70.577 60.564 70.609 60.628 ;
			RECT	70.745 60.564 70.777 60.628 ;
			RECT	70.913 60.564 70.945 60.628 ;
			RECT	71.081 60.564 71.113 60.628 ;
			RECT	71.249 60.564 71.281 60.628 ;
			RECT	71.417 60.564 71.449 60.628 ;
			RECT	71.585 60.564 71.617 60.628 ;
			RECT	71.753 60.564 71.785 60.628 ;
			RECT	71.921 60.564 71.953 60.628 ;
			RECT	72.089 60.564 72.121 60.628 ;
			RECT	72.257 60.564 72.289 60.628 ;
			RECT	72.425 60.564 72.457 60.628 ;
			RECT	72.593 60.564 72.625 60.628 ;
			RECT	72.761 60.564 72.793 60.628 ;
			RECT	72.929 60.564 72.961 60.628 ;
			RECT	73.097 60.564 73.129 60.628 ;
			RECT	73.265 60.564 73.297 60.628 ;
			RECT	73.433 60.564 73.465 60.628 ;
			RECT	73.601 60.564 73.633 60.628 ;
			RECT	73.769 60.564 73.801 60.628 ;
			RECT	73.937 60.564 73.969 60.628 ;
			RECT	74.105 60.564 74.137 60.628 ;
			RECT	74.273 60.564 74.305 60.628 ;
			RECT	74.441 60.564 74.473 60.628 ;
			RECT	74.609 60.564 74.641 60.628 ;
			RECT	74.777 60.564 74.809 60.628 ;
			RECT	74.945 60.564 74.977 60.628 ;
			RECT	75.113 60.564 75.145 60.628 ;
			RECT	75.281 60.564 75.313 60.628 ;
			RECT	75.449 60.564 75.481 60.628 ;
			RECT	75.617 60.564 75.649 60.628 ;
			RECT	75.785 60.564 75.817 60.628 ;
			RECT	75.953 60.564 75.985 60.628 ;
			RECT	76.121 60.564 76.153 60.628 ;
			RECT	76.289 60.564 76.321 60.628 ;
			RECT	76.457 60.564 76.489 60.628 ;
			RECT	76.625 60.564 76.657 60.628 ;
			RECT	76.793 60.564 76.825 60.628 ;
			RECT	76.961 60.564 76.993 60.628 ;
			RECT	77.129 60.564 77.161 60.628 ;
			RECT	77.297 60.564 77.329 60.628 ;
			RECT	77.465 60.564 77.497 60.628 ;
			RECT	77.633 60.564 77.665 60.628 ;
			RECT	77.801 60.564 77.833 60.628 ;
			RECT	77.969 60.564 78.001 60.628 ;
			RECT	78.137 60.564 78.169 60.628 ;
			RECT	78.305 60.564 78.337 60.628 ;
			RECT	78.473 60.564 78.505 60.628 ;
			RECT	78.641 60.564 78.673 60.628 ;
			RECT	78.809 60.564 78.841 60.628 ;
			RECT	78.977 60.564 79.009 60.628 ;
			RECT	79.145 60.564 79.177 60.628 ;
			RECT	79.313 60.564 79.345 60.628 ;
			RECT	79.481 60.564 79.513 60.628 ;
			RECT	79.649 60.564 79.681 60.628 ;
			RECT	79.817 60.564 79.849 60.628 ;
			RECT	79.985 60.564 80.017 60.628 ;
			RECT	80.153 60.564 80.185 60.628 ;
			RECT	80.321 60.564 80.353 60.628 ;
			RECT	80.489 60.564 80.521 60.628 ;
			RECT	80.657 60.564 80.689 60.628 ;
			RECT	80.825 60.564 80.857 60.628 ;
			RECT	80.993 60.564 81.025 60.628 ;
			RECT	81.161 60.564 81.193 60.628 ;
			RECT	81.329 60.564 81.361 60.628 ;
			RECT	81.497 60.564 81.529 60.628 ;
			RECT	81.665 60.564 81.697 60.628 ;
			RECT	81.833 60.564 81.865 60.628 ;
			RECT	82.001 60.564 82.033 60.628 ;
			RECT	82.169 60.564 82.201 60.628 ;
			RECT	82.337 60.564 82.369 60.628 ;
			RECT	82.505 60.564 82.537 60.628 ;
			RECT	82.673 60.564 82.705 60.628 ;
			RECT	82.841 60.564 82.873 60.628 ;
			RECT	83.009 60.564 83.041 60.628 ;
			RECT	83.177 60.564 83.209 60.628 ;
			RECT	83.345 60.564 83.377 60.628 ;
			RECT	83.513 60.564 83.545 60.628 ;
			RECT	83.681 60.564 83.713 60.628 ;
			RECT	83.849 60.564 83.881 60.628 ;
			RECT	84.017 60.564 84.049 60.628 ;
			RECT	84.185 60.564 84.217 60.628 ;
			RECT	84.353 60.564 84.385 60.628 ;
			RECT	84.521 60.564 84.553 60.628 ;
			RECT	84.689 60.564 84.721 60.628 ;
			RECT	84.857 60.564 84.889 60.628 ;
			RECT	85.025 60.564 85.057 60.628 ;
			RECT	85.193 60.564 85.225 60.628 ;
			RECT	85.361 60.564 85.393 60.628 ;
			RECT	85.529 60.564 85.561 60.628 ;
			RECT	85.697 60.564 85.729 60.628 ;
			RECT	85.865 60.564 85.897 60.628 ;
			RECT	86.033 60.564 86.065 60.628 ;
			RECT	86.201 60.564 86.233 60.628 ;
			RECT	86.369 60.564 86.401 60.628 ;
			RECT	86.537 60.564 86.569 60.628 ;
			RECT	86.705 60.564 86.737 60.628 ;
			RECT	86.873 60.564 86.905 60.628 ;
			RECT	87.041 60.564 87.073 60.628 ;
			RECT	87.209 60.564 87.241 60.628 ;
			RECT	87.377 60.564 87.409 60.628 ;
			RECT	87.545 60.564 87.577 60.628 ;
			RECT	87.713 60.564 87.745 60.628 ;
			RECT	87.881 60.564 87.913 60.628 ;
			RECT	88.049 60.564 88.081 60.628 ;
			RECT	88.217 60.564 88.249 60.628 ;
			RECT	88.385 60.564 88.417 60.628 ;
			RECT	88.553 60.564 88.585 60.628 ;
			RECT	88.721 60.564 88.753 60.628 ;
			RECT	88.889 60.564 88.921 60.628 ;
			RECT	89.057 60.564 89.089 60.628 ;
			RECT	89.225 60.564 89.257 60.628 ;
			RECT	89.393 60.564 89.425 60.628 ;
			RECT	89.561 60.564 89.593 60.628 ;
			RECT	89.729 60.564 89.761 60.628 ;
			RECT	89.897 60.564 89.929 60.628 ;
			RECT	90.065 60.564 90.097 60.628 ;
			RECT	90.233 60.564 90.265 60.628 ;
			RECT	90.401 60.564 90.433 60.628 ;
			RECT	90.569 60.564 90.601 60.628 ;
			RECT	90.737 60.564 90.769 60.628 ;
			RECT	90.905 60.564 90.937 60.628 ;
			RECT	91.073 60.564 91.105 60.628 ;
			RECT	91.241 60.564 91.273 60.628 ;
			RECT	91.409 60.564 91.441 60.628 ;
			RECT	91.577 60.564 91.609 60.628 ;
			RECT	91.745 60.564 91.777 60.628 ;
			RECT	91.913 60.564 91.945 60.628 ;
			RECT	92.081 60.564 92.113 60.628 ;
			RECT	92.249 60.564 92.281 60.628 ;
			RECT	92.417 60.564 92.449 60.628 ;
			RECT	92.585 60.564 92.617 60.628 ;
			RECT	92.753 60.564 92.785 60.628 ;
			RECT	92.921 60.564 92.953 60.628 ;
			RECT	93.089 60.564 93.121 60.628 ;
			RECT	93.257 60.564 93.289 60.628 ;
			RECT	93.425 60.564 93.457 60.628 ;
			RECT	93.593 60.564 93.625 60.628 ;
			RECT	93.761 60.564 93.793 60.628 ;
			RECT	93.929 60.564 93.961 60.628 ;
			RECT	94.097 60.564 94.129 60.628 ;
			RECT	94.265 60.564 94.297 60.628 ;
			RECT	94.433 60.564 94.465 60.628 ;
			RECT	94.601 60.564 94.633 60.628 ;
			RECT	94.769 60.564 94.801 60.628 ;
			RECT	94.937 60.564 94.969 60.628 ;
			RECT	95.105 60.564 95.137 60.628 ;
			RECT	95.273 60.564 95.305 60.628 ;
			RECT	95.441 60.564 95.473 60.628 ;
			RECT	95.609 60.564 95.641 60.628 ;
			RECT	95.777 60.564 95.809 60.628 ;
			RECT	95.945 60.564 95.977 60.628 ;
			RECT	96.113 60.564 96.145 60.628 ;
			RECT	96.281 60.564 96.313 60.628 ;
			RECT	96.449 60.564 96.481 60.628 ;
			RECT	96.617 60.564 96.649 60.628 ;
			RECT	96.785 60.564 96.817 60.628 ;
			RECT	96.953 60.564 96.985 60.628 ;
			RECT	97.121 60.564 97.153 60.628 ;
			RECT	97.289 60.564 97.321 60.628 ;
			RECT	97.457 60.564 97.489 60.628 ;
			RECT	97.625 60.564 97.657 60.628 ;
			RECT	97.793 60.564 97.825 60.628 ;
			RECT	97.961 60.564 97.993 60.628 ;
			RECT	98.129 60.564 98.161 60.628 ;
			RECT	98.297 60.564 98.329 60.628 ;
			RECT	98.465 60.564 98.497 60.628 ;
			RECT	98.633 60.564 98.665 60.628 ;
			RECT	98.801 60.564 98.833 60.628 ;
			RECT	98.969 60.564 99.001 60.628 ;
			RECT	99.137 60.564 99.169 60.628 ;
			RECT	99.305 60.564 99.337 60.628 ;
			RECT	99.473 60.564 99.505 60.628 ;
			RECT	99.641 60.564 99.673 60.628 ;
			RECT	99.809 60.564 99.841 60.628 ;
			RECT	99.977 60.564 100.009 60.628 ;
			RECT	100.145 60.564 100.177 60.628 ;
			RECT	100.313 60.564 100.345 60.628 ;
			RECT	100.481 60.564 100.513 60.628 ;
			RECT	100.649 60.564 100.681 60.628 ;
			RECT	100.817 60.564 100.849 60.628 ;
			RECT	100.985 60.564 101.017 60.628 ;
			RECT	101.153 60.564 101.185 60.628 ;
			RECT	101.321 60.564 101.353 60.628 ;
			RECT	101.489 60.564 101.521 60.628 ;
			RECT	101.657 60.564 101.689 60.628 ;
			RECT	101.825 60.564 101.857 60.628 ;
			RECT	101.993 60.564 102.025 60.628 ;
			RECT	102.123 60.58 102.155 60.612 ;
			RECT	102.245 60.575 102.277 60.607 ;
			RECT	102.375 60.564 102.407 60.628 ;
			RECT	103.795 60.564 103.827 60.628 ;
			RECT	103.925 60.575 103.957 60.607 ;
			RECT	104.047 60.58 104.079 60.612 ;
			RECT	104.177 60.564 104.209 60.628 ;
			RECT	104.345 60.564 104.377 60.628 ;
			RECT	104.513 60.564 104.545 60.628 ;
			RECT	104.681 60.564 104.713 60.628 ;
			RECT	104.849 60.564 104.881 60.628 ;
			RECT	105.017 60.564 105.049 60.628 ;
			RECT	105.185 60.564 105.217 60.628 ;
			RECT	105.353 60.564 105.385 60.628 ;
			RECT	105.521 60.564 105.553 60.628 ;
			RECT	105.689 60.564 105.721 60.628 ;
			RECT	105.857 60.564 105.889 60.628 ;
			RECT	106.025 60.564 106.057 60.628 ;
			RECT	106.193 60.564 106.225 60.628 ;
			RECT	106.361 60.564 106.393 60.628 ;
			RECT	106.529 60.564 106.561 60.628 ;
			RECT	106.697 60.564 106.729 60.628 ;
			RECT	106.865 60.564 106.897 60.628 ;
			RECT	107.033 60.564 107.065 60.628 ;
			RECT	107.201 60.564 107.233 60.628 ;
			RECT	107.369 60.564 107.401 60.628 ;
			RECT	107.537 60.564 107.569 60.628 ;
			RECT	107.705 60.564 107.737 60.628 ;
			RECT	107.873 60.564 107.905 60.628 ;
			RECT	108.041 60.564 108.073 60.628 ;
			RECT	108.209 60.564 108.241 60.628 ;
			RECT	108.377 60.564 108.409 60.628 ;
			RECT	108.545 60.564 108.577 60.628 ;
			RECT	108.713 60.564 108.745 60.628 ;
			RECT	108.881 60.564 108.913 60.628 ;
			RECT	109.049 60.564 109.081 60.628 ;
			RECT	109.217 60.564 109.249 60.628 ;
			RECT	109.385 60.564 109.417 60.628 ;
			RECT	109.553 60.564 109.585 60.628 ;
			RECT	109.721 60.564 109.753 60.628 ;
			RECT	109.889 60.564 109.921 60.628 ;
			RECT	110.057 60.564 110.089 60.628 ;
			RECT	110.225 60.564 110.257 60.628 ;
			RECT	110.393 60.564 110.425 60.628 ;
			RECT	110.561 60.564 110.593 60.628 ;
			RECT	110.729 60.564 110.761 60.628 ;
			RECT	110.897 60.564 110.929 60.628 ;
			RECT	111.065 60.564 111.097 60.628 ;
			RECT	111.233 60.564 111.265 60.628 ;
			RECT	111.401 60.564 111.433 60.628 ;
			RECT	111.569 60.564 111.601 60.628 ;
			RECT	111.737 60.564 111.769 60.628 ;
			RECT	111.905 60.564 111.937 60.628 ;
			RECT	112.073 60.564 112.105 60.628 ;
			RECT	112.241 60.564 112.273 60.628 ;
			RECT	112.409 60.564 112.441 60.628 ;
			RECT	112.577 60.564 112.609 60.628 ;
			RECT	112.745 60.564 112.777 60.628 ;
			RECT	112.913 60.564 112.945 60.628 ;
			RECT	113.081 60.564 113.113 60.628 ;
			RECT	113.249 60.564 113.281 60.628 ;
			RECT	113.417 60.564 113.449 60.628 ;
			RECT	113.585 60.564 113.617 60.628 ;
			RECT	113.753 60.564 113.785 60.628 ;
			RECT	113.921 60.564 113.953 60.628 ;
			RECT	114.089 60.564 114.121 60.628 ;
			RECT	114.257 60.564 114.289 60.628 ;
			RECT	114.425 60.564 114.457 60.628 ;
			RECT	114.593 60.564 114.625 60.628 ;
			RECT	114.761 60.564 114.793 60.628 ;
			RECT	114.929 60.564 114.961 60.628 ;
			RECT	115.097 60.564 115.129 60.628 ;
			RECT	115.265 60.564 115.297 60.628 ;
			RECT	115.433 60.564 115.465 60.628 ;
			RECT	115.601 60.564 115.633 60.628 ;
			RECT	115.769 60.564 115.801 60.628 ;
			RECT	115.937 60.564 115.969 60.628 ;
			RECT	116.105 60.564 116.137 60.628 ;
			RECT	116.273 60.564 116.305 60.628 ;
			RECT	116.441 60.564 116.473 60.628 ;
			RECT	116.609 60.564 116.641 60.628 ;
			RECT	116.777 60.564 116.809 60.628 ;
			RECT	116.945 60.564 116.977 60.628 ;
			RECT	117.113 60.564 117.145 60.628 ;
			RECT	117.281 60.564 117.313 60.628 ;
			RECT	117.449 60.564 117.481 60.628 ;
			RECT	117.617 60.564 117.649 60.628 ;
			RECT	117.785 60.564 117.817 60.628 ;
			RECT	117.953 60.564 117.985 60.628 ;
			RECT	118.121 60.564 118.153 60.628 ;
			RECT	118.289 60.564 118.321 60.628 ;
			RECT	118.457 60.564 118.489 60.628 ;
			RECT	118.625 60.564 118.657 60.628 ;
			RECT	118.793 60.564 118.825 60.628 ;
			RECT	118.961 60.564 118.993 60.628 ;
			RECT	119.129 60.564 119.161 60.628 ;
			RECT	119.297 60.564 119.329 60.628 ;
			RECT	119.465 60.564 119.497 60.628 ;
			RECT	119.633 60.564 119.665 60.628 ;
			RECT	119.801 60.564 119.833 60.628 ;
			RECT	119.969 60.564 120.001 60.628 ;
			RECT	120.137 60.564 120.169 60.628 ;
			RECT	120.305 60.564 120.337 60.628 ;
			RECT	120.473 60.564 120.505 60.628 ;
			RECT	120.641 60.564 120.673 60.628 ;
			RECT	120.809 60.564 120.841 60.628 ;
			RECT	120.977 60.564 121.009 60.628 ;
			RECT	121.145 60.564 121.177 60.628 ;
			RECT	121.313 60.564 121.345 60.628 ;
			RECT	121.481 60.564 121.513 60.628 ;
			RECT	121.649 60.564 121.681 60.628 ;
			RECT	121.817 60.564 121.849 60.628 ;
			RECT	121.985 60.564 122.017 60.628 ;
			RECT	122.153 60.564 122.185 60.628 ;
			RECT	122.321 60.564 122.353 60.628 ;
			RECT	122.489 60.564 122.521 60.628 ;
			RECT	122.657 60.564 122.689 60.628 ;
			RECT	122.825 60.564 122.857 60.628 ;
			RECT	122.993 60.564 123.025 60.628 ;
			RECT	123.161 60.564 123.193 60.628 ;
			RECT	123.329 60.564 123.361 60.628 ;
			RECT	123.497 60.564 123.529 60.628 ;
			RECT	123.665 60.564 123.697 60.628 ;
			RECT	123.833 60.564 123.865 60.628 ;
			RECT	124.001 60.564 124.033 60.628 ;
			RECT	124.169 60.564 124.201 60.628 ;
			RECT	124.337 60.564 124.369 60.628 ;
			RECT	124.505 60.564 124.537 60.628 ;
			RECT	124.673 60.564 124.705 60.628 ;
			RECT	124.841 60.564 124.873 60.628 ;
			RECT	125.009 60.564 125.041 60.628 ;
			RECT	125.177 60.564 125.209 60.628 ;
			RECT	125.345 60.564 125.377 60.628 ;
			RECT	125.513 60.564 125.545 60.628 ;
			RECT	125.681 60.564 125.713 60.628 ;
			RECT	125.849 60.564 125.881 60.628 ;
			RECT	126.017 60.564 126.049 60.628 ;
			RECT	126.185 60.564 126.217 60.628 ;
			RECT	126.353 60.564 126.385 60.628 ;
			RECT	126.521 60.564 126.553 60.628 ;
			RECT	126.689 60.564 126.721 60.628 ;
			RECT	126.857 60.564 126.889 60.628 ;
			RECT	127.025 60.564 127.057 60.628 ;
			RECT	127.193 60.564 127.225 60.628 ;
			RECT	127.361 60.564 127.393 60.628 ;
			RECT	127.529 60.564 127.561 60.628 ;
			RECT	127.697 60.564 127.729 60.628 ;
			RECT	127.865 60.564 127.897 60.628 ;
			RECT	128.033 60.564 128.065 60.628 ;
			RECT	128.201 60.564 128.233 60.628 ;
			RECT	128.369 60.564 128.401 60.628 ;
			RECT	128.537 60.564 128.569 60.628 ;
			RECT	128.705 60.564 128.737 60.628 ;
			RECT	128.873 60.564 128.905 60.628 ;
			RECT	129.041 60.564 129.073 60.628 ;
			RECT	129.209 60.564 129.241 60.628 ;
			RECT	129.377 60.564 129.409 60.628 ;
			RECT	129.545 60.564 129.577 60.628 ;
			RECT	129.713 60.564 129.745 60.628 ;
			RECT	129.881 60.564 129.913 60.628 ;
			RECT	130.049 60.564 130.081 60.628 ;
			RECT	130.217 60.564 130.249 60.628 ;
			RECT	130.385 60.564 130.417 60.628 ;
			RECT	130.553 60.564 130.585 60.628 ;
			RECT	130.721 60.564 130.753 60.628 ;
			RECT	130.889 60.564 130.921 60.628 ;
			RECT	131.057 60.564 131.089 60.628 ;
			RECT	131.225 60.564 131.257 60.628 ;
			RECT	131.393 60.564 131.425 60.628 ;
			RECT	131.561 60.564 131.593 60.628 ;
			RECT	131.729 60.564 131.761 60.628 ;
			RECT	131.897 60.564 131.929 60.628 ;
			RECT	132.065 60.564 132.097 60.628 ;
			RECT	132.233 60.564 132.265 60.628 ;
			RECT	132.401 60.564 132.433 60.628 ;
			RECT	132.569 60.564 132.601 60.628 ;
			RECT	132.737 60.564 132.769 60.628 ;
			RECT	132.905 60.564 132.937 60.628 ;
			RECT	133.073 60.564 133.105 60.628 ;
			RECT	133.241 60.564 133.273 60.628 ;
			RECT	133.409 60.564 133.441 60.628 ;
			RECT	133.577 60.564 133.609 60.628 ;
			RECT	133.745 60.564 133.777 60.628 ;
			RECT	133.913 60.564 133.945 60.628 ;
			RECT	134.081 60.564 134.113 60.628 ;
			RECT	134.249 60.564 134.281 60.628 ;
			RECT	134.417 60.564 134.449 60.628 ;
			RECT	134.585 60.564 134.617 60.628 ;
			RECT	134.753 60.564 134.785 60.628 ;
			RECT	134.921 60.564 134.953 60.628 ;
			RECT	135.089 60.564 135.121 60.628 ;
			RECT	135.257 60.564 135.289 60.628 ;
			RECT	135.425 60.564 135.457 60.628 ;
			RECT	135.593 60.564 135.625 60.628 ;
			RECT	135.761 60.564 135.793 60.628 ;
			RECT	135.929 60.564 135.961 60.628 ;
			RECT	136.097 60.564 136.129 60.628 ;
			RECT	136.265 60.564 136.297 60.628 ;
			RECT	136.433 60.564 136.465 60.628 ;
			RECT	136.601 60.564 136.633 60.628 ;
			RECT	136.769 60.564 136.801 60.628 ;
			RECT	136.937 60.564 136.969 60.628 ;
			RECT	137.105 60.564 137.137 60.628 ;
			RECT	137.273 60.564 137.305 60.628 ;
			RECT	137.441 60.564 137.473 60.628 ;
			RECT	137.609 60.564 137.641 60.628 ;
			RECT	137.777 60.564 137.809 60.628 ;
			RECT	137.945 60.564 137.977 60.628 ;
			RECT	138.113 60.564 138.145 60.628 ;
			RECT	138.281 60.564 138.313 60.628 ;
			RECT	138.449 60.564 138.481 60.628 ;
			RECT	138.617 60.564 138.649 60.628 ;
			RECT	138.785 60.564 138.817 60.628 ;
			RECT	138.953 60.564 138.985 60.628 ;
			RECT	139.121 60.564 139.153 60.628 ;
			RECT	139.289 60.564 139.321 60.628 ;
			RECT	139.457 60.564 139.489 60.628 ;
			RECT	139.625 60.564 139.657 60.628 ;
			RECT	139.793 60.564 139.825 60.628 ;
			RECT	139.961 60.564 139.993 60.628 ;
			RECT	140.129 60.564 140.161 60.628 ;
			RECT	140.297 60.564 140.329 60.628 ;
			RECT	140.465 60.564 140.497 60.628 ;
			RECT	140.633 60.564 140.665 60.628 ;
			RECT	140.801 60.564 140.833 60.628 ;
			RECT	140.969 60.564 141.001 60.628 ;
			RECT	141.137 60.564 141.169 60.628 ;
			RECT	141.305 60.564 141.337 60.628 ;
			RECT	141.473 60.564 141.505 60.628 ;
			RECT	141.641 60.564 141.673 60.628 ;
			RECT	141.809 60.564 141.841 60.628 ;
			RECT	141.977 60.564 142.009 60.628 ;
			RECT	142.145 60.564 142.177 60.628 ;
			RECT	142.313 60.564 142.345 60.628 ;
			RECT	142.481 60.564 142.513 60.628 ;
			RECT	142.649 60.564 142.681 60.628 ;
			RECT	142.817 60.564 142.849 60.628 ;
			RECT	142.985 60.564 143.017 60.628 ;
			RECT	143.153 60.564 143.185 60.628 ;
			RECT	143.321 60.564 143.353 60.628 ;
			RECT	143.489 60.564 143.521 60.628 ;
			RECT	143.657 60.564 143.689 60.628 ;
			RECT	143.825 60.564 143.857 60.628 ;
			RECT	143.993 60.564 144.025 60.628 ;
			RECT	144.161 60.564 144.193 60.628 ;
			RECT	144.329 60.564 144.361 60.628 ;
			RECT	144.497 60.564 144.529 60.628 ;
			RECT	144.665 60.564 144.697 60.628 ;
			RECT	144.833 60.564 144.865 60.628 ;
			RECT	145.001 60.564 145.033 60.628 ;
			RECT	145.169 60.564 145.201 60.628 ;
			RECT	145.337 60.564 145.369 60.628 ;
			RECT	145.505 60.564 145.537 60.628 ;
			RECT	145.673 60.564 145.705 60.628 ;
			RECT	145.841 60.564 145.873 60.628 ;
			RECT	146.009 60.564 146.041 60.628 ;
			RECT	146.177 60.564 146.209 60.628 ;
			RECT	146.345 60.564 146.377 60.628 ;
			RECT	146.513 60.564 146.545 60.628 ;
			RECT	146.681 60.564 146.713 60.628 ;
			RECT	146.849 60.564 146.881 60.628 ;
			RECT	147.017 60.564 147.049 60.628 ;
			RECT	147.185 60.564 147.217 60.628 ;
			RECT	147.316 60.58 147.348 60.612 ;
			RECT	147.437 60.58 147.469 60.612 ;
			RECT	147.567 60.564 147.599 60.628 ;
			RECT	149.879 60.564 149.911 60.628 ;
			RECT	151.13 60.564 151.194 60.628 ;
			RECT	151.81 60.564 151.842 60.628 ;
			RECT	152.249 60.564 152.281 60.628 ;
			RECT	153.56 60.564 153.624 60.628 ;
			RECT	156.601 60.564 156.633 60.628 ;
			RECT	156.731 60.58 156.763 60.612 ;
			RECT	156.852 60.58 156.884 60.612 ;
			RECT	156.983 60.564 157.015 60.628 ;
			RECT	157.151 60.564 157.183 60.628 ;
			RECT	157.319 60.564 157.351 60.628 ;
			RECT	157.487 60.564 157.519 60.628 ;
			RECT	157.655 60.564 157.687 60.628 ;
			RECT	157.823 60.564 157.855 60.628 ;
			RECT	157.991 60.564 158.023 60.628 ;
			RECT	158.159 60.564 158.191 60.628 ;
			RECT	158.327 60.564 158.359 60.628 ;
			RECT	158.495 60.564 158.527 60.628 ;
			RECT	158.663 60.564 158.695 60.628 ;
			RECT	158.831 60.564 158.863 60.628 ;
			RECT	158.999 60.564 159.031 60.628 ;
			RECT	159.167 60.564 159.199 60.628 ;
			RECT	159.335 60.564 159.367 60.628 ;
			RECT	159.503 60.564 159.535 60.628 ;
			RECT	159.671 60.564 159.703 60.628 ;
			RECT	159.839 60.564 159.871 60.628 ;
			RECT	160.007 60.564 160.039 60.628 ;
			RECT	160.175 60.564 160.207 60.628 ;
			RECT	160.343 60.564 160.375 60.628 ;
			RECT	160.511 60.564 160.543 60.628 ;
			RECT	160.679 60.564 160.711 60.628 ;
			RECT	160.847 60.564 160.879 60.628 ;
			RECT	161.015 60.564 161.047 60.628 ;
			RECT	161.183 60.564 161.215 60.628 ;
			RECT	161.351 60.564 161.383 60.628 ;
			RECT	161.519 60.564 161.551 60.628 ;
			RECT	161.687 60.564 161.719 60.628 ;
			RECT	161.855 60.564 161.887 60.628 ;
			RECT	162.023 60.564 162.055 60.628 ;
			RECT	162.191 60.564 162.223 60.628 ;
			RECT	162.359 60.564 162.391 60.628 ;
			RECT	162.527 60.564 162.559 60.628 ;
			RECT	162.695 60.564 162.727 60.628 ;
			RECT	162.863 60.564 162.895 60.628 ;
			RECT	163.031 60.564 163.063 60.628 ;
			RECT	163.199 60.564 163.231 60.628 ;
			RECT	163.367 60.564 163.399 60.628 ;
			RECT	163.535 60.564 163.567 60.628 ;
			RECT	163.703 60.564 163.735 60.628 ;
			RECT	163.871 60.564 163.903 60.628 ;
			RECT	164.039 60.564 164.071 60.628 ;
			RECT	164.207 60.564 164.239 60.628 ;
			RECT	164.375 60.564 164.407 60.628 ;
			RECT	164.543 60.564 164.575 60.628 ;
			RECT	164.711 60.564 164.743 60.628 ;
			RECT	164.879 60.564 164.911 60.628 ;
			RECT	165.047 60.564 165.079 60.628 ;
			RECT	165.215 60.564 165.247 60.628 ;
			RECT	165.383 60.564 165.415 60.628 ;
			RECT	165.551 60.564 165.583 60.628 ;
			RECT	165.719 60.564 165.751 60.628 ;
			RECT	165.887 60.564 165.919 60.628 ;
			RECT	166.055 60.564 166.087 60.628 ;
			RECT	166.223 60.564 166.255 60.628 ;
			RECT	166.391 60.564 166.423 60.628 ;
			RECT	166.559 60.564 166.591 60.628 ;
			RECT	166.727 60.564 166.759 60.628 ;
			RECT	166.895 60.564 166.927 60.628 ;
			RECT	167.063 60.564 167.095 60.628 ;
			RECT	167.231 60.564 167.263 60.628 ;
			RECT	167.399 60.564 167.431 60.628 ;
			RECT	167.567 60.564 167.599 60.628 ;
			RECT	167.735 60.564 167.767 60.628 ;
			RECT	167.903 60.564 167.935 60.628 ;
			RECT	168.071 60.564 168.103 60.628 ;
			RECT	168.239 60.564 168.271 60.628 ;
			RECT	168.407 60.564 168.439 60.628 ;
			RECT	168.575 60.564 168.607 60.628 ;
			RECT	168.743 60.564 168.775 60.628 ;
			RECT	168.911 60.564 168.943 60.628 ;
			RECT	169.079 60.564 169.111 60.628 ;
			RECT	169.247 60.564 169.279 60.628 ;
			RECT	169.415 60.564 169.447 60.628 ;
			RECT	169.583 60.564 169.615 60.628 ;
			RECT	169.751 60.564 169.783 60.628 ;
			RECT	169.919 60.564 169.951 60.628 ;
			RECT	170.087 60.564 170.119 60.628 ;
			RECT	170.255 60.564 170.287 60.628 ;
			RECT	170.423 60.564 170.455 60.628 ;
			RECT	170.591 60.564 170.623 60.628 ;
			RECT	170.759 60.564 170.791 60.628 ;
			RECT	170.927 60.564 170.959 60.628 ;
			RECT	171.095 60.564 171.127 60.628 ;
			RECT	171.263 60.564 171.295 60.628 ;
			RECT	171.431 60.564 171.463 60.628 ;
			RECT	171.599 60.564 171.631 60.628 ;
			RECT	171.767 60.564 171.799 60.628 ;
			RECT	171.935 60.564 171.967 60.628 ;
			RECT	172.103 60.564 172.135 60.628 ;
			RECT	172.271 60.564 172.303 60.628 ;
			RECT	172.439 60.564 172.471 60.628 ;
			RECT	172.607 60.564 172.639 60.628 ;
			RECT	172.775 60.564 172.807 60.628 ;
			RECT	172.943 60.564 172.975 60.628 ;
			RECT	173.111 60.564 173.143 60.628 ;
			RECT	173.279 60.564 173.311 60.628 ;
			RECT	173.447 60.564 173.479 60.628 ;
			RECT	173.615 60.564 173.647 60.628 ;
			RECT	173.783 60.564 173.815 60.628 ;
			RECT	173.951 60.564 173.983 60.628 ;
			RECT	174.119 60.564 174.151 60.628 ;
			RECT	174.287 60.564 174.319 60.628 ;
			RECT	174.455 60.564 174.487 60.628 ;
			RECT	174.623 60.564 174.655 60.628 ;
			RECT	174.791 60.564 174.823 60.628 ;
			RECT	174.959 60.564 174.991 60.628 ;
			RECT	175.127 60.564 175.159 60.628 ;
			RECT	175.295 60.564 175.327 60.628 ;
			RECT	175.463 60.564 175.495 60.628 ;
			RECT	175.631 60.564 175.663 60.628 ;
			RECT	175.799 60.564 175.831 60.628 ;
			RECT	175.967 60.564 175.999 60.628 ;
			RECT	176.135 60.564 176.167 60.628 ;
			RECT	176.303 60.564 176.335 60.628 ;
			RECT	176.471 60.564 176.503 60.628 ;
			RECT	176.639 60.564 176.671 60.628 ;
			RECT	176.807 60.564 176.839 60.628 ;
			RECT	176.975 60.564 177.007 60.628 ;
			RECT	177.143 60.564 177.175 60.628 ;
			RECT	177.311 60.564 177.343 60.628 ;
			RECT	177.479 60.564 177.511 60.628 ;
			RECT	177.647 60.564 177.679 60.628 ;
			RECT	177.815 60.564 177.847 60.628 ;
			RECT	177.983 60.564 178.015 60.628 ;
			RECT	178.151 60.564 178.183 60.628 ;
			RECT	178.319 60.564 178.351 60.628 ;
			RECT	178.487 60.564 178.519 60.628 ;
			RECT	178.655 60.564 178.687 60.628 ;
			RECT	178.823 60.564 178.855 60.628 ;
			RECT	178.991 60.564 179.023 60.628 ;
			RECT	179.159 60.564 179.191 60.628 ;
			RECT	179.327 60.564 179.359 60.628 ;
			RECT	179.495 60.564 179.527 60.628 ;
			RECT	179.663 60.564 179.695 60.628 ;
			RECT	179.831 60.564 179.863 60.628 ;
			RECT	179.999 60.564 180.031 60.628 ;
			RECT	180.167 60.564 180.199 60.628 ;
			RECT	180.335 60.564 180.367 60.628 ;
			RECT	180.503 60.564 180.535 60.628 ;
			RECT	180.671 60.564 180.703 60.628 ;
			RECT	180.839 60.564 180.871 60.628 ;
			RECT	181.007 60.564 181.039 60.628 ;
			RECT	181.175 60.564 181.207 60.628 ;
			RECT	181.343 60.564 181.375 60.628 ;
			RECT	181.511 60.564 181.543 60.628 ;
			RECT	181.679 60.564 181.711 60.628 ;
			RECT	181.847 60.564 181.879 60.628 ;
			RECT	182.015 60.564 182.047 60.628 ;
			RECT	182.183 60.564 182.215 60.628 ;
			RECT	182.351 60.564 182.383 60.628 ;
			RECT	182.519 60.564 182.551 60.628 ;
			RECT	182.687 60.564 182.719 60.628 ;
			RECT	182.855 60.564 182.887 60.628 ;
			RECT	183.023 60.564 183.055 60.628 ;
			RECT	183.191 60.564 183.223 60.628 ;
			RECT	183.359 60.564 183.391 60.628 ;
			RECT	183.527 60.564 183.559 60.628 ;
			RECT	183.695 60.564 183.727 60.628 ;
			RECT	183.863 60.564 183.895 60.628 ;
			RECT	184.031 60.564 184.063 60.628 ;
			RECT	184.199 60.564 184.231 60.628 ;
			RECT	184.367 60.564 184.399 60.628 ;
			RECT	184.535 60.564 184.567 60.628 ;
			RECT	184.703 60.564 184.735 60.628 ;
			RECT	184.871 60.564 184.903 60.628 ;
			RECT	185.039 60.564 185.071 60.628 ;
			RECT	185.207 60.564 185.239 60.628 ;
			RECT	185.375 60.564 185.407 60.628 ;
			RECT	185.543 60.564 185.575 60.628 ;
			RECT	185.711 60.564 185.743 60.628 ;
			RECT	185.879 60.564 185.911 60.628 ;
			RECT	186.047 60.564 186.079 60.628 ;
			RECT	186.215 60.564 186.247 60.628 ;
			RECT	186.383 60.564 186.415 60.628 ;
			RECT	186.551 60.564 186.583 60.628 ;
			RECT	186.719 60.564 186.751 60.628 ;
			RECT	186.887 60.564 186.919 60.628 ;
			RECT	187.055 60.564 187.087 60.628 ;
			RECT	187.223 60.564 187.255 60.628 ;
			RECT	187.391 60.564 187.423 60.628 ;
			RECT	187.559 60.564 187.591 60.628 ;
			RECT	187.727 60.564 187.759 60.628 ;
			RECT	187.895 60.564 187.927 60.628 ;
			RECT	188.063 60.564 188.095 60.628 ;
			RECT	188.231 60.564 188.263 60.628 ;
			RECT	188.399 60.564 188.431 60.628 ;
			RECT	188.567 60.564 188.599 60.628 ;
			RECT	188.735 60.564 188.767 60.628 ;
			RECT	188.903 60.564 188.935 60.628 ;
			RECT	189.071 60.564 189.103 60.628 ;
			RECT	189.239 60.564 189.271 60.628 ;
			RECT	189.407 60.564 189.439 60.628 ;
			RECT	189.575 60.564 189.607 60.628 ;
			RECT	189.743 60.564 189.775 60.628 ;
			RECT	189.911 60.564 189.943 60.628 ;
			RECT	190.079 60.564 190.111 60.628 ;
			RECT	190.247 60.564 190.279 60.628 ;
			RECT	190.415 60.564 190.447 60.628 ;
			RECT	190.583 60.564 190.615 60.628 ;
			RECT	190.751 60.564 190.783 60.628 ;
			RECT	190.919 60.564 190.951 60.628 ;
			RECT	191.087 60.564 191.119 60.628 ;
			RECT	191.255 60.564 191.287 60.628 ;
			RECT	191.423 60.564 191.455 60.628 ;
			RECT	191.591 60.564 191.623 60.628 ;
			RECT	191.759 60.564 191.791 60.628 ;
			RECT	191.927 60.564 191.959 60.628 ;
			RECT	192.095 60.564 192.127 60.628 ;
			RECT	192.263 60.564 192.295 60.628 ;
			RECT	192.431 60.564 192.463 60.628 ;
			RECT	192.599 60.564 192.631 60.628 ;
			RECT	192.767 60.564 192.799 60.628 ;
			RECT	192.935 60.564 192.967 60.628 ;
			RECT	193.103 60.564 193.135 60.628 ;
			RECT	193.271 60.564 193.303 60.628 ;
			RECT	193.439 60.564 193.471 60.628 ;
			RECT	193.607 60.564 193.639 60.628 ;
			RECT	193.775 60.564 193.807 60.628 ;
			RECT	193.943 60.564 193.975 60.628 ;
			RECT	194.111 60.564 194.143 60.628 ;
			RECT	194.279 60.564 194.311 60.628 ;
			RECT	194.447 60.564 194.479 60.628 ;
			RECT	194.615 60.564 194.647 60.628 ;
			RECT	194.783 60.564 194.815 60.628 ;
			RECT	194.951 60.564 194.983 60.628 ;
			RECT	195.119 60.564 195.151 60.628 ;
			RECT	195.287 60.564 195.319 60.628 ;
			RECT	195.455 60.564 195.487 60.628 ;
			RECT	195.623 60.564 195.655 60.628 ;
			RECT	195.791 60.564 195.823 60.628 ;
			RECT	195.959 60.564 195.991 60.628 ;
			RECT	196.127 60.564 196.159 60.628 ;
			RECT	196.295 60.564 196.327 60.628 ;
			RECT	196.463 60.564 196.495 60.628 ;
			RECT	196.631 60.564 196.663 60.628 ;
			RECT	196.799 60.564 196.831 60.628 ;
			RECT	196.967 60.564 196.999 60.628 ;
			RECT	197.135 60.564 197.167 60.628 ;
			RECT	197.303 60.564 197.335 60.628 ;
			RECT	197.471 60.564 197.503 60.628 ;
			RECT	197.639 60.564 197.671 60.628 ;
			RECT	197.807 60.564 197.839 60.628 ;
			RECT	197.975 60.564 198.007 60.628 ;
			RECT	198.143 60.564 198.175 60.628 ;
			RECT	198.311 60.564 198.343 60.628 ;
			RECT	198.479 60.564 198.511 60.628 ;
			RECT	198.647 60.564 198.679 60.628 ;
			RECT	198.815 60.564 198.847 60.628 ;
			RECT	198.983 60.564 199.015 60.628 ;
			RECT	199.151 60.564 199.183 60.628 ;
			RECT	199.319 60.564 199.351 60.628 ;
			RECT	199.487 60.564 199.519 60.628 ;
			RECT	199.655 60.564 199.687 60.628 ;
			RECT	199.823 60.564 199.855 60.628 ;
			RECT	199.991 60.564 200.023 60.628 ;
			RECT	200.121 60.58 200.153 60.612 ;
			RECT	200.243 60.575 200.275 60.607 ;
			RECT	200.373 60.564 200.405 60.628 ;
			RECT	200.9 60.564 200.932 60.628 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 58.616 201.665 58.736 ;
			LAYER	J3 ;
			RECT	0.755 58.644 0.787 58.708 ;
			RECT	1.645 58.644 1.709 58.708 ;
			RECT	2.323 58.644 2.387 58.708 ;
			RECT	3.438 58.644 3.47 58.708 ;
			RECT	3.585 58.644 3.617 58.708 ;
			RECT	4.195 58.644 4.227 58.708 ;
			RECT	4.72 58.644 4.752 58.708 ;
			RECT	4.944 58.644 5.008 58.708 ;
			RECT	5.267 58.644 5.299 58.708 ;
			RECT	5.797 58.644 5.829 58.708 ;
			RECT	5.927 58.655 5.959 58.687 ;
			RECT	6.049 58.66 6.081 58.692 ;
			RECT	6.179 58.644 6.211 58.708 ;
			RECT	6.347 58.644 6.379 58.708 ;
			RECT	6.515 58.644 6.547 58.708 ;
			RECT	6.683 58.644 6.715 58.708 ;
			RECT	6.851 58.644 6.883 58.708 ;
			RECT	7.019 58.644 7.051 58.708 ;
			RECT	7.187 58.644 7.219 58.708 ;
			RECT	7.355 58.644 7.387 58.708 ;
			RECT	7.523 58.644 7.555 58.708 ;
			RECT	7.691 58.644 7.723 58.708 ;
			RECT	7.859 58.644 7.891 58.708 ;
			RECT	8.027 58.644 8.059 58.708 ;
			RECT	8.195 58.644 8.227 58.708 ;
			RECT	8.363 58.644 8.395 58.708 ;
			RECT	8.531 58.644 8.563 58.708 ;
			RECT	8.699 58.644 8.731 58.708 ;
			RECT	8.867 58.644 8.899 58.708 ;
			RECT	9.035 58.644 9.067 58.708 ;
			RECT	9.203 58.644 9.235 58.708 ;
			RECT	9.371 58.644 9.403 58.708 ;
			RECT	9.539 58.644 9.571 58.708 ;
			RECT	9.707 58.644 9.739 58.708 ;
			RECT	9.875 58.644 9.907 58.708 ;
			RECT	10.043 58.644 10.075 58.708 ;
			RECT	10.211 58.644 10.243 58.708 ;
			RECT	10.379 58.644 10.411 58.708 ;
			RECT	10.547 58.644 10.579 58.708 ;
			RECT	10.715 58.644 10.747 58.708 ;
			RECT	10.883 58.644 10.915 58.708 ;
			RECT	11.051 58.644 11.083 58.708 ;
			RECT	11.219 58.644 11.251 58.708 ;
			RECT	11.387 58.644 11.419 58.708 ;
			RECT	11.555 58.644 11.587 58.708 ;
			RECT	11.723 58.644 11.755 58.708 ;
			RECT	11.891 58.644 11.923 58.708 ;
			RECT	12.059 58.644 12.091 58.708 ;
			RECT	12.227 58.644 12.259 58.708 ;
			RECT	12.395 58.644 12.427 58.708 ;
			RECT	12.563 58.644 12.595 58.708 ;
			RECT	12.731 58.644 12.763 58.708 ;
			RECT	12.899 58.644 12.931 58.708 ;
			RECT	13.067 58.644 13.099 58.708 ;
			RECT	13.235 58.644 13.267 58.708 ;
			RECT	13.403 58.644 13.435 58.708 ;
			RECT	13.571 58.644 13.603 58.708 ;
			RECT	13.739 58.644 13.771 58.708 ;
			RECT	13.907 58.644 13.939 58.708 ;
			RECT	14.075 58.644 14.107 58.708 ;
			RECT	14.243 58.644 14.275 58.708 ;
			RECT	14.411 58.644 14.443 58.708 ;
			RECT	14.579 58.644 14.611 58.708 ;
			RECT	14.747 58.644 14.779 58.708 ;
			RECT	14.915 58.644 14.947 58.708 ;
			RECT	15.083 58.644 15.115 58.708 ;
			RECT	15.251 58.644 15.283 58.708 ;
			RECT	15.419 58.644 15.451 58.708 ;
			RECT	15.587 58.644 15.619 58.708 ;
			RECT	15.755 58.644 15.787 58.708 ;
			RECT	15.923 58.644 15.955 58.708 ;
			RECT	16.091 58.644 16.123 58.708 ;
			RECT	16.259 58.644 16.291 58.708 ;
			RECT	16.427 58.644 16.459 58.708 ;
			RECT	16.595 58.644 16.627 58.708 ;
			RECT	16.763 58.644 16.795 58.708 ;
			RECT	16.931 58.644 16.963 58.708 ;
			RECT	17.099 58.644 17.131 58.708 ;
			RECT	17.267 58.644 17.299 58.708 ;
			RECT	17.435 58.644 17.467 58.708 ;
			RECT	17.603 58.644 17.635 58.708 ;
			RECT	17.771 58.644 17.803 58.708 ;
			RECT	17.939 58.644 17.971 58.708 ;
			RECT	18.107 58.644 18.139 58.708 ;
			RECT	18.275 58.644 18.307 58.708 ;
			RECT	18.443 58.644 18.475 58.708 ;
			RECT	18.611 58.644 18.643 58.708 ;
			RECT	18.779 58.644 18.811 58.708 ;
			RECT	18.947 58.644 18.979 58.708 ;
			RECT	19.115 58.644 19.147 58.708 ;
			RECT	19.283 58.644 19.315 58.708 ;
			RECT	19.451 58.644 19.483 58.708 ;
			RECT	19.619 58.644 19.651 58.708 ;
			RECT	19.787 58.644 19.819 58.708 ;
			RECT	19.955 58.644 19.987 58.708 ;
			RECT	20.123 58.644 20.155 58.708 ;
			RECT	20.291 58.644 20.323 58.708 ;
			RECT	20.459 58.644 20.491 58.708 ;
			RECT	20.627 58.644 20.659 58.708 ;
			RECT	20.795 58.644 20.827 58.708 ;
			RECT	20.963 58.644 20.995 58.708 ;
			RECT	21.131 58.644 21.163 58.708 ;
			RECT	21.299 58.644 21.331 58.708 ;
			RECT	21.467 58.644 21.499 58.708 ;
			RECT	21.635 58.644 21.667 58.708 ;
			RECT	21.803 58.644 21.835 58.708 ;
			RECT	21.971 58.644 22.003 58.708 ;
			RECT	22.139 58.644 22.171 58.708 ;
			RECT	22.307 58.644 22.339 58.708 ;
			RECT	22.475 58.644 22.507 58.708 ;
			RECT	22.643 58.644 22.675 58.708 ;
			RECT	22.811 58.644 22.843 58.708 ;
			RECT	22.979 58.644 23.011 58.708 ;
			RECT	23.147 58.644 23.179 58.708 ;
			RECT	23.315 58.644 23.347 58.708 ;
			RECT	23.483 58.644 23.515 58.708 ;
			RECT	23.651 58.644 23.683 58.708 ;
			RECT	23.819 58.644 23.851 58.708 ;
			RECT	23.987 58.644 24.019 58.708 ;
			RECT	24.155 58.644 24.187 58.708 ;
			RECT	24.323 58.644 24.355 58.708 ;
			RECT	24.491 58.644 24.523 58.708 ;
			RECT	24.659 58.644 24.691 58.708 ;
			RECT	24.827 58.644 24.859 58.708 ;
			RECT	24.995 58.644 25.027 58.708 ;
			RECT	25.163 58.644 25.195 58.708 ;
			RECT	25.331 58.644 25.363 58.708 ;
			RECT	25.499 58.644 25.531 58.708 ;
			RECT	25.667 58.644 25.699 58.708 ;
			RECT	25.835 58.644 25.867 58.708 ;
			RECT	26.003 58.644 26.035 58.708 ;
			RECT	26.171 58.644 26.203 58.708 ;
			RECT	26.339 58.644 26.371 58.708 ;
			RECT	26.507 58.644 26.539 58.708 ;
			RECT	26.675 58.644 26.707 58.708 ;
			RECT	26.843 58.644 26.875 58.708 ;
			RECT	27.011 58.644 27.043 58.708 ;
			RECT	27.179 58.644 27.211 58.708 ;
			RECT	27.347 58.644 27.379 58.708 ;
			RECT	27.515 58.644 27.547 58.708 ;
			RECT	27.683 58.644 27.715 58.708 ;
			RECT	27.851 58.644 27.883 58.708 ;
			RECT	28.019 58.644 28.051 58.708 ;
			RECT	28.187 58.644 28.219 58.708 ;
			RECT	28.355 58.644 28.387 58.708 ;
			RECT	28.523 58.644 28.555 58.708 ;
			RECT	28.691 58.644 28.723 58.708 ;
			RECT	28.859 58.644 28.891 58.708 ;
			RECT	29.027 58.644 29.059 58.708 ;
			RECT	29.195 58.644 29.227 58.708 ;
			RECT	29.363 58.644 29.395 58.708 ;
			RECT	29.531 58.644 29.563 58.708 ;
			RECT	29.699 58.644 29.731 58.708 ;
			RECT	29.867 58.644 29.899 58.708 ;
			RECT	30.035 58.644 30.067 58.708 ;
			RECT	30.203 58.644 30.235 58.708 ;
			RECT	30.371 58.644 30.403 58.708 ;
			RECT	30.539 58.644 30.571 58.708 ;
			RECT	30.707 58.644 30.739 58.708 ;
			RECT	30.875 58.644 30.907 58.708 ;
			RECT	31.043 58.644 31.075 58.708 ;
			RECT	31.211 58.644 31.243 58.708 ;
			RECT	31.379 58.644 31.411 58.708 ;
			RECT	31.547 58.644 31.579 58.708 ;
			RECT	31.715 58.644 31.747 58.708 ;
			RECT	31.883 58.644 31.915 58.708 ;
			RECT	32.051 58.644 32.083 58.708 ;
			RECT	32.219 58.644 32.251 58.708 ;
			RECT	32.387 58.644 32.419 58.708 ;
			RECT	32.555 58.644 32.587 58.708 ;
			RECT	32.723 58.644 32.755 58.708 ;
			RECT	32.891 58.644 32.923 58.708 ;
			RECT	33.059 58.644 33.091 58.708 ;
			RECT	33.227 58.644 33.259 58.708 ;
			RECT	33.395 58.644 33.427 58.708 ;
			RECT	33.563 58.644 33.595 58.708 ;
			RECT	33.731 58.644 33.763 58.708 ;
			RECT	33.899 58.644 33.931 58.708 ;
			RECT	34.067 58.644 34.099 58.708 ;
			RECT	34.235 58.644 34.267 58.708 ;
			RECT	34.403 58.644 34.435 58.708 ;
			RECT	34.571 58.644 34.603 58.708 ;
			RECT	34.739 58.644 34.771 58.708 ;
			RECT	34.907 58.644 34.939 58.708 ;
			RECT	35.075 58.644 35.107 58.708 ;
			RECT	35.243 58.644 35.275 58.708 ;
			RECT	35.411 58.644 35.443 58.708 ;
			RECT	35.579 58.644 35.611 58.708 ;
			RECT	35.747 58.644 35.779 58.708 ;
			RECT	35.915 58.644 35.947 58.708 ;
			RECT	36.083 58.644 36.115 58.708 ;
			RECT	36.251 58.644 36.283 58.708 ;
			RECT	36.419 58.644 36.451 58.708 ;
			RECT	36.587 58.644 36.619 58.708 ;
			RECT	36.755 58.644 36.787 58.708 ;
			RECT	36.923 58.644 36.955 58.708 ;
			RECT	37.091 58.644 37.123 58.708 ;
			RECT	37.259 58.644 37.291 58.708 ;
			RECT	37.427 58.644 37.459 58.708 ;
			RECT	37.595 58.644 37.627 58.708 ;
			RECT	37.763 58.644 37.795 58.708 ;
			RECT	37.931 58.644 37.963 58.708 ;
			RECT	38.099 58.644 38.131 58.708 ;
			RECT	38.267 58.644 38.299 58.708 ;
			RECT	38.435 58.644 38.467 58.708 ;
			RECT	38.603 58.644 38.635 58.708 ;
			RECT	38.771 58.644 38.803 58.708 ;
			RECT	38.939 58.644 38.971 58.708 ;
			RECT	39.107 58.644 39.139 58.708 ;
			RECT	39.275 58.644 39.307 58.708 ;
			RECT	39.443 58.644 39.475 58.708 ;
			RECT	39.611 58.644 39.643 58.708 ;
			RECT	39.779 58.644 39.811 58.708 ;
			RECT	39.947 58.644 39.979 58.708 ;
			RECT	40.115 58.644 40.147 58.708 ;
			RECT	40.283 58.644 40.315 58.708 ;
			RECT	40.451 58.644 40.483 58.708 ;
			RECT	40.619 58.644 40.651 58.708 ;
			RECT	40.787 58.644 40.819 58.708 ;
			RECT	40.955 58.644 40.987 58.708 ;
			RECT	41.123 58.644 41.155 58.708 ;
			RECT	41.291 58.644 41.323 58.708 ;
			RECT	41.459 58.644 41.491 58.708 ;
			RECT	41.627 58.644 41.659 58.708 ;
			RECT	41.795 58.644 41.827 58.708 ;
			RECT	41.963 58.644 41.995 58.708 ;
			RECT	42.131 58.644 42.163 58.708 ;
			RECT	42.299 58.644 42.331 58.708 ;
			RECT	42.467 58.644 42.499 58.708 ;
			RECT	42.635 58.644 42.667 58.708 ;
			RECT	42.803 58.644 42.835 58.708 ;
			RECT	42.971 58.644 43.003 58.708 ;
			RECT	43.139 58.644 43.171 58.708 ;
			RECT	43.307 58.644 43.339 58.708 ;
			RECT	43.475 58.644 43.507 58.708 ;
			RECT	43.643 58.644 43.675 58.708 ;
			RECT	43.811 58.644 43.843 58.708 ;
			RECT	43.979 58.644 44.011 58.708 ;
			RECT	44.147 58.644 44.179 58.708 ;
			RECT	44.315 58.644 44.347 58.708 ;
			RECT	44.483 58.644 44.515 58.708 ;
			RECT	44.651 58.644 44.683 58.708 ;
			RECT	44.819 58.644 44.851 58.708 ;
			RECT	44.987 58.644 45.019 58.708 ;
			RECT	45.155 58.644 45.187 58.708 ;
			RECT	45.323 58.644 45.355 58.708 ;
			RECT	45.491 58.644 45.523 58.708 ;
			RECT	45.659 58.644 45.691 58.708 ;
			RECT	45.827 58.644 45.859 58.708 ;
			RECT	45.995 58.644 46.027 58.708 ;
			RECT	46.163 58.644 46.195 58.708 ;
			RECT	46.331 58.644 46.363 58.708 ;
			RECT	46.499 58.644 46.531 58.708 ;
			RECT	46.667 58.644 46.699 58.708 ;
			RECT	46.835 58.644 46.867 58.708 ;
			RECT	47.003 58.644 47.035 58.708 ;
			RECT	47.171 58.644 47.203 58.708 ;
			RECT	47.339 58.644 47.371 58.708 ;
			RECT	47.507 58.644 47.539 58.708 ;
			RECT	47.675 58.644 47.707 58.708 ;
			RECT	47.843 58.644 47.875 58.708 ;
			RECT	48.011 58.644 48.043 58.708 ;
			RECT	48.179 58.644 48.211 58.708 ;
			RECT	48.347 58.644 48.379 58.708 ;
			RECT	48.515 58.644 48.547 58.708 ;
			RECT	48.683 58.644 48.715 58.708 ;
			RECT	48.851 58.644 48.883 58.708 ;
			RECT	49.019 58.644 49.051 58.708 ;
			RECT	49.187 58.644 49.219 58.708 ;
			RECT	49.318 58.66 49.35 58.692 ;
			RECT	49.439 58.66 49.471 58.692 ;
			RECT	49.569 58.644 49.601 58.708 ;
			RECT	51.881 58.644 51.913 58.708 ;
			RECT	53.132 58.644 53.196 58.708 ;
			RECT	53.812 58.644 53.844 58.708 ;
			RECT	54.251 58.644 54.283 58.708 ;
			RECT	55.562 58.644 55.626 58.708 ;
			RECT	58.603 58.644 58.635 58.708 ;
			RECT	58.733 58.66 58.765 58.692 ;
			RECT	58.854 58.66 58.886 58.692 ;
			RECT	58.985 58.644 59.017 58.708 ;
			RECT	59.153 58.644 59.185 58.708 ;
			RECT	59.321 58.644 59.353 58.708 ;
			RECT	59.489 58.644 59.521 58.708 ;
			RECT	59.657 58.644 59.689 58.708 ;
			RECT	59.825 58.644 59.857 58.708 ;
			RECT	59.993 58.644 60.025 58.708 ;
			RECT	60.161 58.644 60.193 58.708 ;
			RECT	60.329 58.644 60.361 58.708 ;
			RECT	60.497 58.644 60.529 58.708 ;
			RECT	60.665 58.644 60.697 58.708 ;
			RECT	60.833 58.644 60.865 58.708 ;
			RECT	61.001 58.644 61.033 58.708 ;
			RECT	61.169 58.644 61.201 58.708 ;
			RECT	61.337 58.644 61.369 58.708 ;
			RECT	61.505 58.644 61.537 58.708 ;
			RECT	61.673 58.644 61.705 58.708 ;
			RECT	61.841 58.644 61.873 58.708 ;
			RECT	62.009 58.644 62.041 58.708 ;
			RECT	62.177 58.644 62.209 58.708 ;
			RECT	62.345 58.644 62.377 58.708 ;
			RECT	62.513 58.644 62.545 58.708 ;
			RECT	62.681 58.644 62.713 58.708 ;
			RECT	62.849 58.644 62.881 58.708 ;
			RECT	63.017 58.644 63.049 58.708 ;
			RECT	63.185 58.644 63.217 58.708 ;
			RECT	63.353 58.644 63.385 58.708 ;
			RECT	63.521 58.644 63.553 58.708 ;
			RECT	63.689 58.644 63.721 58.708 ;
			RECT	63.857 58.644 63.889 58.708 ;
			RECT	64.025 58.644 64.057 58.708 ;
			RECT	64.193 58.644 64.225 58.708 ;
			RECT	64.361 58.644 64.393 58.708 ;
			RECT	64.529 58.644 64.561 58.708 ;
			RECT	64.697 58.644 64.729 58.708 ;
			RECT	64.865 58.644 64.897 58.708 ;
			RECT	65.033 58.644 65.065 58.708 ;
			RECT	65.201 58.644 65.233 58.708 ;
			RECT	65.369 58.644 65.401 58.708 ;
			RECT	65.537 58.644 65.569 58.708 ;
			RECT	65.705 58.644 65.737 58.708 ;
			RECT	65.873 58.644 65.905 58.708 ;
			RECT	66.041 58.644 66.073 58.708 ;
			RECT	66.209 58.644 66.241 58.708 ;
			RECT	66.377 58.644 66.409 58.708 ;
			RECT	66.545 58.644 66.577 58.708 ;
			RECT	66.713 58.644 66.745 58.708 ;
			RECT	66.881 58.644 66.913 58.708 ;
			RECT	67.049 58.644 67.081 58.708 ;
			RECT	67.217 58.644 67.249 58.708 ;
			RECT	67.385 58.644 67.417 58.708 ;
			RECT	67.553 58.644 67.585 58.708 ;
			RECT	67.721 58.644 67.753 58.708 ;
			RECT	67.889 58.644 67.921 58.708 ;
			RECT	68.057 58.644 68.089 58.708 ;
			RECT	68.225 58.644 68.257 58.708 ;
			RECT	68.393 58.644 68.425 58.708 ;
			RECT	68.561 58.644 68.593 58.708 ;
			RECT	68.729 58.644 68.761 58.708 ;
			RECT	68.897 58.644 68.929 58.708 ;
			RECT	69.065 58.644 69.097 58.708 ;
			RECT	69.233 58.644 69.265 58.708 ;
			RECT	69.401 58.644 69.433 58.708 ;
			RECT	69.569 58.644 69.601 58.708 ;
			RECT	69.737 58.644 69.769 58.708 ;
			RECT	69.905 58.644 69.937 58.708 ;
			RECT	70.073 58.644 70.105 58.708 ;
			RECT	70.241 58.644 70.273 58.708 ;
			RECT	70.409 58.644 70.441 58.708 ;
			RECT	70.577 58.644 70.609 58.708 ;
			RECT	70.745 58.644 70.777 58.708 ;
			RECT	70.913 58.644 70.945 58.708 ;
			RECT	71.081 58.644 71.113 58.708 ;
			RECT	71.249 58.644 71.281 58.708 ;
			RECT	71.417 58.644 71.449 58.708 ;
			RECT	71.585 58.644 71.617 58.708 ;
			RECT	71.753 58.644 71.785 58.708 ;
			RECT	71.921 58.644 71.953 58.708 ;
			RECT	72.089 58.644 72.121 58.708 ;
			RECT	72.257 58.644 72.289 58.708 ;
			RECT	72.425 58.644 72.457 58.708 ;
			RECT	72.593 58.644 72.625 58.708 ;
			RECT	72.761 58.644 72.793 58.708 ;
			RECT	72.929 58.644 72.961 58.708 ;
			RECT	73.097 58.644 73.129 58.708 ;
			RECT	73.265 58.644 73.297 58.708 ;
			RECT	73.433 58.644 73.465 58.708 ;
			RECT	73.601 58.644 73.633 58.708 ;
			RECT	73.769 58.644 73.801 58.708 ;
			RECT	73.937 58.644 73.969 58.708 ;
			RECT	74.105 58.644 74.137 58.708 ;
			RECT	74.273 58.644 74.305 58.708 ;
			RECT	74.441 58.644 74.473 58.708 ;
			RECT	74.609 58.644 74.641 58.708 ;
			RECT	74.777 58.644 74.809 58.708 ;
			RECT	74.945 58.644 74.977 58.708 ;
			RECT	75.113 58.644 75.145 58.708 ;
			RECT	75.281 58.644 75.313 58.708 ;
			RECT	75.449 58.644 75.481 58.708 ;
			RECT	75.617 58.644 75.649 58.708 ;
			RECT	75.785 58.644 75.817 58.708 ;
			RECT	75.953 58.644 75.985 58.708 ;
			RECT	76.121 58.644 76.153 58.708 ;
			RECT	76.289 58.644 76.321 58.708 ;
			RECT	76.457 58.644 76.489 58.708 ;
			RECT	76.625 58.644 76.657 58.708 ;
			RECT	76.793 58.644 76.825 58.708 ;
			RECT	76.961 58.644 76.993 58.708 ;
			RECT	77.129 58.644 77.161 58.708 ;
			RECT	77.297 58.644 77.329 58.708 ;
			RECT	77.465 58.644 77.497 58.708 ;
			RECT	77.633 58.644 77.665 58.708 ;
			RECT	77.801 58.644 77.833 58.708 ;
			RECT	77.969 58.644 78.001 58.708 ;
			RECT	78.137 58.644 78.169 58.708 ;
			RECT	78.305 58.644 78.337 58.708 ;
			RECT	78.473 58.644 78.505 58.708 ;
			RECT	78.641 58.644 78.673 58.708 ;
			RECT	78.809 58.644 78.841 58.708 ;
			RECT	78.977 58.644 79.009 58.708 ;
			RECT	79.145 58.644 79.177 58.708 ;
			RECT	79.313 58.644 79.345 58.708 ;
			RECT	79.481 58.644 79.513 58.708 ;
			RECT	79.649 58.644 79.681 58.708 ;
			RECT	79.817 58.644 79.849 58.708 ;
			RECT	79.985 58.644 80.017 58.708 ;
			RECT	80.153 58.644 80.185 58.708 ;
			RECT	80.321 58.644 80.353 58.708 ;
			RECT	80.489 58.644 80.521 58.708 ;
			RECT	80.657 58.644 80.689 58.708 ;
			RECT	80.825 58.644 80.857 58.708 ;
			RECT	80.993 58.644 81.025 58.708 ;
			RECT	81.161 58.644 81.193 58.708 ;
			RECT	81.329 58.644 81.361 58.708 ;
			RECT	81.497 58.644 81.529 58.708 ;
			RECT	81.665 58.644 81.697 58.708 ;
			RECT	81.833 58.644 81.865 58.708 ;
			RECT	82.001 58.644 82.033 58.708 ;
			RECT	82.169 58.644 82.201 58.708 ;
			RECT	82.337 58.644 82.369 58.708 ;
			RECT	82.505 58.644 82.537 58.708 ;
			RECT	82.673 58.644 82.705 58.708 ;
			RECT	82.841 58.644 82.873 58.708 ;
			RECT	83.009 58.644 83.041 58.708 ;
			RECT	83.177 58.644 83.209 58.708 ;
			RECT	83.345 58.644 83.377 58.708 ;
			RECT	83.513 58.644 83.545 58.708 ;
			RECT	83.681 58.644 83.713 58.708 ;
			RECT	83.849 58.644 83.881 58.708 ;
			RECT	84.017 58.644 84.049 58.708 ;
			RECT	84.185 58.644 84.217 58.708 ;
			RECT	84.353 58.644 84.385 58.708 ;
			RECT	84.521 58.644 84.553 58.708 ;
			RECT	84.689 58.644 84.721 58.708 ;
			RECT	84.857 58.644 84.889 58.708 ;
			RECT	85.025 58.644 85.057 58.708 ;
			RECT	85.193 58.644 85.225 58.708 ;
			RECT	85.361 58.644 85.393 58.708 ;
			RECT	85.529 58.644 85.561 58.708 ;
			RECT	85.697 58.644 85.729 58.708 ;
			RECT	85.865 58.644 85.897 58.708 ;
			RECT	86.033 58.644 86.065 58.708 ;
			RECT	86.201 58.644 86.233 58.708 ;
			RECT	86.369 58.644 86.401 58.708 ;
			RECT	86.537 58.644 86.569 58.708 ;
			RECT	86.705 58.644 86.737 58.708 ;
			RECT	86.873 58.644 86.905 58.708 ;
			RECT	87.041 58.644 87.073 58.708 ;
			RECT	87.209 58.644 87.241 58.708 ;
			RECT	87.377 58.644 87.409 58.708 ;
			RECT	87.545 58.644 87.577 58.708 ;
			RECT	87.713 58.644 87.745 58.708 ;
			RECT	87.881 58.644 87.913 58.708 ;
			RECT	88.049 58.644 88.081 58.708 ;
			RECT	88.217 58.644 88.249 58.708 ;
			RECT	88.385 58.644 88.417 58.708 ;
			RECT	88.553 58.644 88.585 58.708 ;
			RECT	88.721 58.644 88.753 58.708 ;
			RECT	88.889 58.644 88.921 58.708 ;
			RECT	89.057 58.644 89.089 58.708 ;
			RECT	89.225 58.644 89.257 58.708 ;
			RECT	89.393 58.644 89.425 58.708 ;
			RECT	89.561 58.644 89.593 58.708 ;
			RECT	89.729 58.644 89.761 58.708 ;
			RECT	89.897 58.644 89.929 58.708 ;
			RECT	90.065 58.644 90.097 58.708 ;
			RECT	90.233 58.644 90.265 58.708 ;
			RECT	90.401 58.644 90.433 58.708 ;
			RECT	90.569 58.644 90.601 58.708 ;
			RECT	90.737 58.644 90.769 58.708 ;
			RECT	90.905 58.644 90.937 58.708 ;
			RECT	91.073 58.644 91.105 58.708 ;
			RECT	91.241 58.644 91.273 58.708 ;
			RECT	91.409 58.644 91.441 58.708 ;
			RECT	91.577 58.644 91.609 58.708 ;
			RECT	91.745 58.644 91.777 58.708 ;
			RECT	91.913 58.644 91.945 58.708 ;
			RECT	92.081 58.644 92.113 58.708 ;
			RECT	92.249 58.644 92.281 58.708 ;
			RECT	92.417 58.644 92.449 58.708 ;
			RECT	92.585 58.644 92.617 58.708 ;
			RECT	92.753 58.644 92.785 58.708 ;
			RECT	92.921 58.644 92.953 58.708 ;
			RECT	93.089 58.644 93.121 58.708 ;
			RECT	93.257 58.644 93.289 58.708 ;
			RECT	93.425 58.644 93.457 58.708 ;
			RECT	93.593 58.644 93.625 58.708 ;
			RECT	93.761 58.644 93.793 58.708 ;
			RECT	93.929 58.644 93.961 58.708 ;
			RECT	94.097 58.644 94.129 58.708 ;
			RECT	94.265 58.644 94.297 58.708 ;
			RECT	94.433 58.644 94.465 58.708 ;
			RECT	94.601 58.644 94.633 58.708 ;
			RECT	94.769 58.644 94.801 58.708 ;
			RECT	94.937 58.644 94.969 58.708 ;
			RECT	95.105 58.644 95.137 58.708 ;
			RECT	95.273 58.644 95.305 58.708 ;
			RECT	95.441 58.644 95.473 58.708 ;
			RECT	95.609 58.644 95.641 58.708 ;
			RECT	95.777 58.644 95.809 58.708 ;
			RECT	95.945 58.644 95.977 58.708 ;
			RECT	96.113 58.644 96.145 58.708 ;
			RECT	96.281 58.644 96.313 58.708 ;
			RECT	96.449 58.644 96.481 58.708 ;
			RECT	96.617 58.644 96.649 58.708 ;
			RECT	96.785 58.644 96.817 58.708 ;
			RECT	96.953 58.644 96.985 58.708 ;
			RECT	97.121 58.644 97.153 58.708 ;
			RECT	97.289 58.644 97.321 58.708 ;
			RECT	97.457 58.644 97.489 58.708 ;
			RECT	97.625 58.644 97.657 58.708 ;
			RECT	97.793 58.644 97.825 58.708 ;
			RECT	97.961 58.644 97.993 58.708 ;
			RECT	98.129 58.644 98.161 58.708 ;
			RECT	98.297 58.644 98.329 58.708 ;
			RECT	98.465 58.644 98.497 58.708 ;
			RECT	98.633 58.644 98.665 58.708 ;
			RECT	98.801 58.644 98.833 58.708 ;
			RECT	98.969 58.644 99.001 58.708 ;
			RECT	99.137 58.644 99.169 58.708 ;
			RECT	99.305 58.644 99.337 58.708 ;
			RECT	99.473 58.644 99.505 58.708 ;
			RECT	99.641 58.644 99.673 58.708 ;
			RECT	99.809 58.644 99.841 58.708 ;
			RECT	99.977 58.644 100.009 58.708 ;
			RECT	100.145 58.644 100.177 58.708 ;
			RECT	100.313 58.644 100.345 58.708 ;
			RECT	100.481 58.644 100.513 58.708 ;
			RECT	100.649 58.644 100.681 58.708 ;
			RECT	100.817 58.644 100.849 58.708 ;
			RECT	100.985 58.644 101.017 58.708 ;
			RECT	101.153 58.644 101.185 58.708 ;
			RECT	101.321 58.644 101.353 58.708 ;
			RECT	101.489 58.644 101.521 58.708 ;
			RECT	101.657 58.644 101.689 58.708 ;
			RECT	101.825 58.644 101.857 58.708 ;
			RECT	101.993 58.644 102.025 58.708 ;
			RECT	102.123 58.66 102.155 58.692 ;
			RECT	102.245 58.655 102.277 58.687 ;
			RECT	102.375 58.644 102.407 58.708 ;
			RECT	103.795 58.644 103.827 58.708 ;
			RECT	103.925 58.655 103.957 58.687 ;
			RECT	104.047 58.66 104.079 58.692 ;
			RECT	104.177 58.644 104.209 58.708 ;
			RECT	104.345 58.644 104.377 58.708 ;
			RECT	104.513 58.644 104.545 58.708 ;
			RECT	104.681 58.644 104.713 58.708 ;
			RECT	104.849 58.644 104.881 58.708 ;
			RECT	105.017 58.644 105.049 58.708 ;
			RECT	105.185 58.644 105.217 58.708 ;
			RECT	105.353 58.644 105.385 58.708 ;
			RECT	105.521 58.644 105.553 58.708 ;
			RECT	105.689 58.644 105.721 58.708 ;
			RECT	105.857 58.644 105.889 58.708 ;
			RECT	106.025 58.644 106.057 58.708 ;
			RECT	106.193 58.644 106.225 58.708 ;
			RECT	106.361 58.644 106.393 58.708 ;
			RECT	106.529 58.644 106.561 58.708 ;
			RECT	106.697 58.644 106.729 58.708 ;
			RECT	106.865 58.644 106.897 58.708 ;
			RECT	107.033 58.644 107.065 58.708 ;
			RECT	107.201 58.644 107.233 58.708 ;
			RECT	107.369 58.644 107.401 58.708 ;
			RECT	107.537 58.644 107.569 58.708 ;
			RECT	107.705 58.644 107.737 58.708 ;
			RECT	107.873 58.644 107.905 58.708 ;
			RECT	108.041 58.644 108.073 58.708 ;
			RECT	108.209 58.644 108.241 58.708 ;
			RECT	108.377 58.644 108.409 58.708 ;
			RECT	108.545 58.644 108.577 58.708 ;
			RECT	108.713 58.644 108.745 58.708 ;
			RECT	108.881 58.644 108.913 58.708 ;
			RECT	109.049 58.644 109.081 58.708 ;
			RECT	109.217 58.644 109.249 58.708 ;
			RECT	109.385 58.644 109.417 58.708 ;
			RECT	109.553 58.644 109.585 58.708 ;
			RECT	109.721 58.644 109.753 58.708 ;
			RECT	109.889 58.644 109.921 58.708 ;
			RECT	110.057 58.644 110.089 58.708 ;
			RECT	110.225 58.644 110.257 58.708 ;
			RECT	110.393 58.644 110.425 58.708 ;
			RECT	110.561 58.644 110.593 58.708 ;
			RECT	110.729 58.644 110.761 58.708 ;
			RECT	110.897 58.644 110.929 58.708 ;
			RECT	111.065 58.644 111.097 58.708 ;
			RECT	111.233 58.644 111.265 58.708 ;
			RECT	111.401 58.644 111.433 58.708 ;
			RECT	111.569 58.644 111.601 58.708 ;
			RECT	111.737 58.644 111.769 58.708 ;
			RECT	111.905 58.644 111.937 58.708 ;
			RECT	112.073 58.644 112.105 58.708 ;
			RECT	112.241 58.644 112.273 58.708 ;
			RECT	112.409 58.644 112.441 58.708 ;
			RECT	112.577 58.644 112.609 58.708 ;
			RECT	112.745 58.644 112.777 58.708 ;
			RECT	112.913 58.644 112.945 58.708 ;
			RECT	113.081 58.644 113.113 58.708 ;
			RECT	113.249 58.644 113.281 58.708 ;
			RECT	113.417 58.644 113.449 58.708 ;
			RECT	113.585 58.644 113.617 58.708 ;
			RECT	113.753 58.644 113.785 58.708 ;
			RECT	113.921 58.644 113.953 58.708 ;
			RECT	114.089 58.644 114.121 58.708 ;
			RECT	114.257 58.644 114.289 58.708 ;
			RECT	114.425 58.644 114.457 58.708 ;
			RECT	114.593 58.644 114.625 58.708 ;
			RECT	114.761 58.644 114.793 58.708 ;
			RECT	114.929 58.644 114.961 58.708 ;
			RECT	115.097 58.644 115.129 58.708 ;
			RECT	115.265 58.644 115.297 58.708 ;
			RECT	115.433 58.644 115.465 58.708 ;
			RECT	115.601 58.644 115.633 58.708 ;
			RECT	115.769 58.644 115.801 58.708 ;
			RECT	115.937 58.644 115.969 58.708 ;
			RECT	116.105 58.644 116.137 58.708 ;
			RECT	116.273 58.644 116.305 58.708 ;
			RECT	116.441 58.644 116.473 58.708 ;
			RECT	116.609 58.644 116.641 58.708 ;
			RECT	116.777 58.644 116.809 58.708 ;
			RECT	116.945 58.644 116.977 58.708 ;
			RECT	117.113 58.644 117.145 58.708 ;
			RECT	117.281 58.644 117.313 58.708 ;
			RECT	117.449 58.644 117.481 58.708 ;
			RECT	117.617 58.644 117.649 58.708 ;
			RECT	117.785 58.644 117.817 58.708 ;
			RECT	117.953 58.644 117.985 58.708 ;
			RECT	118.121 58.644 118.153 58.708 ;
			RECT	118.289 58.644 118.321 58.708 ;
			RECT	118.457 58.644 118.489 58.708 ;
			RECT	118.625 58.644 118.657 58.708 ;
			RECT	118.793 58.644 118.825 58.708 ;
			RECT	118.961 58.644 118.993 58.708 ;
			RECT	119.129 58.644 119.161 58.708 ;
			RECT	119.297 58.644 119.329 58.708 ;
			RECT	119.465 58.644 119.497 58.708 ;
			RECT	119.633 58.644 119.665 58.708 ;
			RECT	119.801 58.644 119.833 58.708 ;
			RECT	119.969 58.644 120.001 58.708 ;
			RECT	120.137 58.644 120.169 58.708 ;
			RECT	120.305 58.644 120.337 58.708 ;
			RECT	120.473 58.644 120.505 58.708 ;
			RECT	120.641 58.644 120.673 58.708 ;
			RECT	120.809 58.644 120.841 58.708 ;
			RECT	120.977 58.644 121.009 58.708 ;
			RECT	121.145 58.644 121.177 58.708 ;
			RECT	121.313 58.644 121.345 58.708 ;
			RECT	121.481 58.644 121.513 58.708 ;
			RECT	121.649 58.644 121.681 58.708 ;
			RECT	121.817 58.644 121.849 58.708 ;
			RECT	121.985 58.644 122.017 58.708 ;
			RECT	122.153 58.644 122.185 58.708 ;
			RECT	122.321 58.644 122.353 58.708 ;
			RECT	122.489 58.644 122.521 58.708 ;
			RECT	122.657 58.644 122.689 58.708 ;
			RECT	122.825 58.644 122.857 58.708 ;
			RECT	122.993 58.644 123.025 58.708 ;
			RECT	123.161 58.644 123.193 58.708 ;
			RECT	123.329 58.644 123.361 58.708 ;
			RECT	123.497 58.644 123.529 58.708 ;
			RECT	123.665 58.644 123.697 58.708 ;
			RECT	123.833 58.644 123.865 58.708 ;
			RECT	124.001 58.644 124.033 58.708 ;
			RECT	124.169 58.644 124.201 58.708 ;
			RECT	124.337 58.644 124.369 58.708 ;
			RECT	124.505 58.644 124.537 58.708 ;
			RECT	124.673 58.644 124.705 58.708 ;
			RECT	124.841 58.644 124.873 58.708 ;
			RECT	125.009 58.644 125.041 58.708 ;
			RECT	125.177 58.644 125.209 58.708 ;
			RECT	125.345 58.644 125.377 58.708 ;
			RECT	125.513 58.644 125.545 58.708 ;
			RECT	125.681 58.644 125.713 58.708 ;
			RECT	125.849 58.644 125.881 58.708 ;
			RECT	126.017 58.644 126.049 58.708 ;
			RECT	126.185 58.644 126.217 58.708 ;
			RECT	126.353 58.644 126.385 58.708 ;
			RECT	126.521 58.644 126.553 58.708 ;
			RECT	126.689 58.644 126.721 58.708 ;
			RECT	126.857 58.644 126.889 58.708 ;
			RECT	127.025 58.644 127.057 58.708 ;
			RECT	127.193 58.644 127.225 58.708 ;
			RECT	127.361 58.644 127.393 58.708 ;
			RECT	127.529 58.644 127.561 58.708 ;
			RECT	127.697 58.644 127.729 58.708 ;
			RECT	127.865 58.644 127.897 58.708 ;
			RECT	128.033 58.644 128.065 58.708 ;
			RECT	128.201 58.644 128.233 58.708 ;
			RECT	128.369 58.644 128.401 58.708 ;
			RECT	128.537 58.644 128.569 58.708 ;
			RECT	128.705 58.644 128.737 58.708 ;
			RECT	128.873 58.644 128.905 58.708 ;
			RECT	129.041 58.644 129.073 58.708 ;
			RECT	129.209 58.644 129.241 58.708 ;
			RECT	129.377 58.644 129.409 58.708 ;
			RECT	129.545 58.644 129.577 58.708 ;
			RECT	129.713 58.644 129.745 58.708 ;
			RECT	129.881 58.644 129.913 58.708 ;
			RECT	130.049 58.644 130.081 58.708 ;
			RECT	130.217 58.644 130.249 58.708 ;
			RECT	130.385 58.644 130.417 58.708 ;
			RECT	130.553 58.644 130.585 58.708 ;
			RECT	130.721 58.644 130.753 58.708 ;
			RECT	130.889 58.644 130.921 58.708 ;
			RECT	131.057 58.644 131.089 58.708 ;
			RECT	131.225 58.644 131.257 58.708 ;
			RECT	131.393 58.644 131.425 58.708 ;
			RECT	131.561 58.644 131.593 58.708 ;
			RECT	131.729 58.644 131.761 58.708 ;
			RECT	131.897 58.644 131.929 58.708 ;
			RECT	132.065 58.644 132.097 58.708 ;
			RECT	132.233 58.644 132.265 58.708 ;
			RECT	132.401 58.644 132.433 58.708 ;
			RECT	132.569 58.644 132.601 58.708 ;
			RECT	132.737 58.644 132.769 58.708 ;
			RECT	132.905 58.644 132.937 58.708 ;
			RECT	133.073 58.644 133.105 58.708 ;
			RECT	133.241 58.644 133.273 58.708 ;
			RECT	133.409 58.644 133.441 58.708 ;
			RECT	133.577 58.644 133.609 58.708 ;
			RECT	133.745 58.644 133.777 58.708 ;
			RECT	133.913 58.644 133.945 58.708 ;
			RECT	134.081 58.644 134.113 58.708 ;
			RECT	134.249 58.644 134.281 58.708 ;
			RECT	134.417 58.644 134.449 58.708 ;
			RECT	134.585 58.644 134.617 58.708 ;
			RECT	134.753 58.644 134.785 58.708 ;
			RECT	134.921 58.644 134.953 58.708 ;
			RECT	135.089 58.644 135.121 58.708 ;
			RECT	135.257 58.644 135.289 58.708 ;
			RECT	135.425 58.644 135.457 58.708 ;
			RECT	135.593 58.644 135.625 58.708 ;
			RECT	135.761 58.644 135.793 58.708 ;
			RECT	135.929 58.644 135.961 58.708 ;
			RECT	136.097 58.644 136.129 58.708 ;
			RECT	136.265 58.644 136.297 58.708 ;
			RECT	136.433 58.644 136.465 58.708 ;
			RECT	136.601 58.644 136.633 58.708 ;
			RECT	136.769 58.644 136.801 58.708 ;
			RECT	136.937 58.644 136.969 58.708 ;
			RECT	137.105 58.644 137.137 58.708 ;
			RECT	137.273 58.644 137.305 58.708 ;
			RECT	137.441 58.644 137.473 58.708 ;
			RECT	137.609 58.644 137.641 58.708 ;
			RECT	137.777 58.644 137.809 58.708 ;
			RECT	137.945 58.644 137.977 58.708 ;
			RECT	138.113 58.644 138.145 58.708 ;
			RECT	138.281 58.644 138.313 58.708 ;
			RECT	138.449 58.644 138.481 58.708 ;
			RECT	138.617 58.644 138.649 58.708 ;
			RECT	138.785 58.644 138.817 58.708 ;
			RECT	138.953 58.644 138.985 58.708 ;
			RECT	139.121 58.644 139.153 58.708 ;
			RECT	139.289 58.644 139.321 58.708 ;
			RECT	139.457 58.644 139.489 58.708 ;
			RECT	139.625 58.644 139.657 58.708 ;
			RECT	139.793 58.644 139.825 58.708 ;
			RECT	139.961 58.644 139.993 58.708 ;
			RECT	140.129 58.644 140.161 58.708 ;
			RECT	140.297 58.644 140.329 58.708 ;
			RECT	140.465 58.644 140.497 58.708 ;
			RECT	140.633 58.644 140.665 58.708 ;
			RECT	140.801 58.644 140.833 58.708 ;
			RECT	140.969 58.644 141.001 58.708 ;
			RECT	141.137 58.644 141.169 58.708 ;
			RECT	141.305 58.644 141.337 58.708 ;
			RECT	141.473 58.644 141.505 58.708 ;
			RECT	141.641 58.644 141.673 58.708 ;
			RECT	141.809 58.644 141.841 58.708 ;
			RECT	141.977 58.644 142.009 58.708 ;
			RECT	142.145 58.644 142.177 58.708 ;
			RECT	142.313 58.644 142.345 58.708 ;
			RECT	142.481 58.644 142.513 58.708 ;
			RECT	142.649 58.644 142.681 58.708 ;
			RECT	142.817 58.644 142.849 58.708 ;
			RECT	142.985 58.644 143.017 58.708 ;
			RECT	143.153 58.644 143.185 58.708 ;
			RECT	143.321 58.644 143.353 58.708 ;
			RECT	143.489 58.644 143.521 58.708 ;
			RECT	143.657 58.644 143.689 58.708 ;
			RECT	143.825 58.644 143.857 58.708 ;
			RECT	143.993 58.644 144.025 58.708 ;
			RECT	144.161 58.644 144.193 58.708 ;
			RECT	144.329 58.644 144.361 58.708 ;
			RECT	144.497 58.644 144.529 58.708 ;
			RECT	144.665 58.644 144.697 58.708 ;
			RECT	144.833 58.644 144.865 58.708 ;
			RECT	145.001 58.644 145.033 58.708 ;
			RECT	145.169 58.644 145.201 58.708 ;
			RECT	145.337 58.644 145.369 58.708 ;
			RECT	145.505 58.644 145.537 58.708 ;
			RECT	145.673 58.644 145.705 58.708 ;
			RECT	145.841 58.644 145.873 58.708 ;
			RECT	146.009 58.644 146.041 58.708 ;
			RECT	146.177 58.644 146.209 58.708 ;
			RECT	146.345 58.644 146.377 58.708 ;
			RECT	146.513 58.644 146.545 58.708 ;
			RECT	146.681 58.644 146.713 58.708 ;
			RECT	146.849 58.644 146.881 58.708 ;
			RECT	147.017 58.644 147.049 58.708 ;
			RECT	147.185 58.644 147.217 58.708 ;
			RECT	147.316 58.66 147.348 58.692 ;
			RECT	147.437 58.66 147.469 58.692 ;
			RECT	147.567 58.644 147.599 58.708 ;
			RECT	149.879 58.644 149.911 58.708 ;
			RECT	151.13 58.644 151.194 58.708 ;
			RECT	151.81 58.644 151.842 58.708 ;
			RECT	152.249 58.644 152.281 58.708 ;
			RECT	153.56 58.644 153.624 58.708 ;
			RECT	156.601 58.644 156.633 58.708 ;
			RECT	156.731 58.66 156.763 58.692 ;
			RECT	156.852 58.66 156.884 58.692 ;
			RECT	156.983 58.644 157.015 58.708 ;
			RECT	157.151 58.644 157.183 58.708 ;
			RECT	157.319 58.644 157.351 58.708 ;
			RECT	157.487 58.644 157.519 58.708 ;
			RECT	157.655 58.644 157.687 58.708 ;
			RECT	157.823 58.644 157.855 58.708 ;
			RECT	157.991 58.644 158.023 58.708 ;
			RECT	158.159 58.644 158.191 58.708 ;
			RECT	158.327 58.644 158.359 58.708 ;
			RECT	158.495 58.644 158.527 58.708 ;
			RECT	158.663 58.644 158.695 58.708 ;
			RECT	158.831 58.644 158.863 58.708 ;
			RECT	158.999 58.644 159.031 58.708 ;
			RECT	159.167 58.644 159.199 58.708 ;
			RECT	159.335 58.644 159.367 58.708 ;
			RECT	159.503 58.644 159.535 58.708 ;
			RECT	159.671 58.644 159.703 58.708 ;
			RECT	159.839 58.644 159.871 58.708 ;
			RECT	160.007 58.644 160.039 58.708 ;
			RECT	160.175 58.644 160.207 58.708 ;
			RECT	160.343 58.644 160.375 58.708 ;
			RECT	160.511 58.644 160.543 58.708 ;
			RECT	160.679 58.644 160.711 58.708 ;
			RECT	160.847 58.644 160.879 58.708 ;
			RECT	161.015 58.644 161.047 58.708 ;
			RECT	161.183 58.644 161.215 58.708 ;
			RECT	161.351 58.644 161.383 58.708 ;
			RECT	161.519 58.644 161.551 58.708 ;
			RECT	161.687 58.644 161.719 58.708 ;
			RECT	161.855 58.644 161.887 58.708 ;
			RECT	162.023 58.644 162.055 58.708 ;
			RECT	162.191 58.644 162.223 58.708 ;
			RECT	162.359 58.644 162.391 58.708 ;
			RECT	162.527 58.644 162.559 58.708 ;
			RECT	162.695 58.644 162.727 58.708 ;
			RECT	162.863 58.644 162.895 58.708 ;
			RECT	163.031 58.644 163.063 58.708 ;
			RECT	163.199 58.644 163.231 58.708 ;
			RECT	163.367 58.644 163.399 58.708 ;
			RECT	163.535 58.644 163.567 58.708 ;
			RECT	163.703 58.644 163.735 58.708 ;
			RECT	163.871 58.644 163.903 58.708 ;
			RECT	164.039 58.644 164.071 58.708 ;
			RECT	164.207 58.644 164.239 58.708 ;
			RECT	164.375 58.644 164.407 58.708 ;
			RECT	164.543 58.644 164.575 58.708 ;
			RECT	164.711 58.644 164.743 58.708 ;
			RECT	164.879 58.644 164.911 58.708 ;
			RECT	165.047 58.644 165.079 58.708 ;
			RECT	165.215 58.644 165.247 58.708 ;
			RECT	165.383 58.644 165.415 58.708 ;
			RECT	165.551 58.644 165.583 58.708 ;
			RECT	165.719 58.644 165.751 58.708 ;
			RECT	165.887 58.644 165.919 58.708 ;
			RECT	166.055 58.644 166.087 58.708 ;
			RECT	166.223 58.644 166.255 58.708 ;
			RECT	166.391 58.644 166.423 58.708 ;
			RECT	166.559 58.644 166.591 58.708 ;
			RECT	166.727 58.644 166.759 58.708 ;
			RECT	166.895 58.644 166.927 58.708 ;
			RECT	167.063 58.644 167.095 58.708 ;
			RECT	167.231 58.644 167.263 58.708 ;
			RECT	167.399 58.644 167.431 58.708 ;
			RECT	167.567 58.644 167.599 58.708 ;
			RECT	167.735 58.644 167.767 58.708 ;
			RECT	167.903 58.644 167.935 58.708 ;
			RECT	168.071 58.644 168.103 58.708 ;
			RECT	168.239 58.644 168.271 58.708 ;
			RECT	168.407 58.644 168.439 58.708 ;
			RECT	168.575 58.644 168.607 58.708 ;
			RECT	168.743 58.644 168.775 58.708 ;
			RECT	168.911 58.644 168.943 58.708 ;
			RECT	169.079 58.644 169.111 58.708 ;
			RECT	169.247 58.644 169.279 58.708 ;
			RECT	169.415 58.644 169.447 58.708 ;
			RECT	169.583 58.644 169.615 58.708 ;
			RECT	169.751 58.644 169.783 58.708 ;
			RECT	169.919 58.644 169.951 58.708 ;
			RECT	170.087 58.644 170.119 58.708 ;
			RECT	170.255 58.644 170.287 58.708 ;
			RECT	170.423 58.644 170.455 58.708 ;
			RECT	170.591 58.644 170.623 58.708 ;
			RECT	170.759 58.644 170.791 58.708 ;
			RECT	170.927 58.644 170.959 58.708 ;
			RECT	171.095 58.644 171.127 58.708 ;
			RECT	171.263 58.644 171.295 58.708 ;
			RECT	171.431 58.644 171.463 58.708 ;
			RECT	171.599 58.644 171.631 58.708 ;
			RECT	171.767 58.644 171.799 58.708 ;
			RECT	171.935 58.644 171.967 58.708 ;
			RECT	172.103 58.644 172.135 58.708 ;
			RECT	172.271 58.644 172.303 58.708 ;
			RECT	172.439 58.644 172.471 58.708 ;
			RECT	172.607 58.644 172.639 58.708 ;
			RECT	172.775 58.644 172.807 58.708 ;
			RECT	172.943 58.644 172.975 58.708 ;
			RECT	173.111 58.644 173.143 58.708 ;
			RECT	173.279 58.644 173.311 58.708 ;
			RECT	173.447 58.644 173.479 58.708 ;
			RECT	173.615 58.644 173.647 58.708 ;
			RECT	173.783 58.644 173.815 58.708 ;
			RECT	173.951 58.644 173.983 58.708 ;
			RECT	174.119 58.644 174.151 58.708 ;
			RECT	174.287 58.644 174.319 58.708 ;
			RECT	174.455 58.644 174.487 58.708 ;
			RECT	174.623 58.644 174.655 58.708 ;
			RECT	174.791 58.644 174.823 58.708 ;
			RECT	174.959 58.644 174.991 58.708 ;
			RECT	175.127 58.644 175.159 58.708 ;
			RECT	175.295 58.644 175.327 58.708 ;
			RECT	175.463 58.644 175.495 58.708 ;
			RECT	175.631 58.644 175.663 58.708 ;
			RECT	175.799 58.644 175.831 58.708 ;
			RECT	175.967 58.644 175.999 58.708 ;
			RECT	176.135 58.644 176.167 58.708 ;
			RECT	176.303 58.644 176.335 58.708 ;
			RECT	176.471 58.644 176.503 58.708 ;
			RECT	176.639 58.644 176.671 58.708 ;
			RECT	176.807 58.644 176.839 58.708 ;
			RECT	176.975 58.644 177.007 58.708 ;
			RECT	177.143 58.644 177.175 58.708 ;
			RECT	177.311 58.644 177.343 58.708 ;
			RECT	177.479 58.644 177.511 58.708 ;
			RECT	177.647 58.644 177.679 58.708 ;
			RECT	177.815 58.644 177.847 58.708 ;
			RECT	177.983 58.644 178.015 58.708 ;
			RECT	178.151 58.644 178.183 58.708 ;
			RECT	178.319 58.644 178.351 58.708 ;
			RECT	178.487 58.644 178.519 58.708 ;
			RECT	178.655 58.644 178.687 58.708 ;
			RECT	178.823 58.644 178.855 58.708 ;
			RECT	178.991 58.644 179.023 58.708 ;
			RECT	179.159 58.644 179.191 58.708 ;
			RECT	179.327 58.644 179.359 58.708 ;
			RECT	179.495 58.644 179.527 58.708 ;
			RECT	179.663 58.644 179.695 58.708 ;
			RECT	179.831 58.644 179.863 58.708 ;
			RECT	179.999 58.644 180.031 58.708 ;
			RECT	180.167 58.644 180.199 58.708 ;
			RECT	180.335 58.644 180.367 58.708 ;
			RECT	180.503 58.644 180.535 58.708 ;
			RECT	180.671 58.644 180.703 58.708 ;
			RECT	180.839 58.644 180.871 58.708 ;
			RECT	181.007 58.644 181.039 58.708 ;
			RECT	181.175 58.644 181.207 58.708 ;
			RECT	181.343 58.644 181.375 58.708 ;
			RECT	181.511 58.644 181.543 58.708 ;
			RECT	181.679 58.644 181.711 58.708 ;
			RECT	181.847 58.644 181.879 58.708 ;
			RECT	182.015 58.644 182.047 58.708 ;
			RECT	182.183 58.644 182.215 58.708 ;
			RECT	182.351 58.644 182.383 58.708 ;
			RECT	182.519 58.644 182.551 58.708 ;
			RECT	182.687 58.644 182.719 58.708 ;
			RECT	182.855 58.644 182.887 58.708 ;
			RECT	183.023 58.644 183.055 58.708 ;
			RECT	183.191 58.644 183.223 58.708 ;
			RECT	183.359 58.644 183.391 58.708 ;
			RECT	183.527 58.644 183.559 58.708 ;
			RECT	183.695 58.644 183.727 58.708 ;
			RECT	183.863 58.644 183.895 58.708 ;
			RECT	184.031 58.644 184.063 58.708 ;
			RECT	184.199 58.644 184.231 58.708 ;
			RECT	184.367 58.644 184.399 58.708 ;
			RECT	184.535 58.644 184.567 58.708 ;
			RECT	184.703 58.644 184.735 58.708 ;
			RECT	184.871 58.644 184.903 58.708 ;
			RECT	185.039 58.644 185.071 58.708 ;
			RECT	185.207 58.644 185.239 58.708 ;
			RECT	185.375 58.644 185.407 58.708 ;
			RECT	185.543 58.644 185.575 58.708 ;
			RECT	185.711 58.644 185.743 58.708 ;
			RECT	185.879 58.644 185.911 58.708 ;
			RECT	186.047 58.644 186.079 58.708 ;
			RECT	186.215 58.644 186.247 58.708 ;
			RECT	186.383 58.644 186.415 58.708 ;
			RECT	186.551 58.644 186.583 58.708 ;
			RECT	186.719 58.644 186.751 58.708 ;
			RECT	186.887 58.644 186.919 58.708 ;
			RECT	187.055 58.644 187.087 58.708 ;
			RECT	187.223 58.644 187.255 58.708 ;
			RECT	187.391 58.644 187.423 58.708 ;
			RECT	187.559 58.644 187.591 58.708 ;
			RECT	187.727 58.644 187.759 58.708 ;
			RECT	187.895 58.644 187.927 58.708 ;
			RECT	188.063 58.644 188.095 58.708 ;
			RECT	188.231 58.644 188.263 58.708 ;
			RECT	188.399 58.644 188.431 58.708 ;
			RECT	188.567 58.644 188.599 58.708 ;
			RECT	188.735 58.644 188.767 58.708 ;
			RECT	188.903 58.644 188.935 58.708 ;
			RECT	189.071 58.644 189.103 58.708 ;
			RECT	189.239 58.644 189.271 58.708 ;
			RECT	189.407 58.644 189.439 58.708 ;
			RECT	189.575 58.644 189.607 58.708 ;
			RECT	189.743 58.644 189.775 58.708 ;
			RECT	189.911 58.644 189.943 58.708 ;
			RECT	190.079 58.644 190.111 58.708 ;
			RECT	190.247 58.644 190.279 58.708 ;
			RECT	190.415 58.644 190.447 58.708 ;
			RECT	190.583 58.644 190.615 58.708 ;
			RECT	190.751 58.644 190.783 58.708 ;
			RECT	190.919 58.644 190.951 58.708 ;
			RECT	191.087 58.644 191.119 58.708 ;
			RECT	191.255 58.644 191.287 58.708 ;
			RECT	191.423 58.644 191.455 58.708 ;
			RECT	191.591 58.644 191.623 58.708 ;
			RECT	191.759 58.644 191.791 58.708 ;
			RECT	191.927 58.644 191.959 58.708 ;
			RECT	192.095 58.644 192.127 58.708 ;
			RECT	192.263 58.644 192.295 58.708 ;
			RECT	192.431 58.644 192.463 58.708 ;
			RECT	192.599 58.644 192.631 58.708 ;
			RECT	192.767 58.644 192.799 58.708 ;
			RECT	192.935 58.644 192.967 58.708 ;
			RECT	193.103 58.644 193.135 58.708 ;
			RECT	193.271 58.644 193.303 58.708 ;
			RECT	193.439 58.644 193.471 58.708 ;
			RECT	193.607 58.644 193.639 58.708 ;
			RECT	193.775 58.644 193.807 58.708 ;
			RECT	193.943 58.644 193.975 58.708 ;
			RECT	194.111 58.644 194.143 58.708 ;
			RECT	194.279 58.644 194.311 58.708 ;
			RECT	194.447 58.644 194.479 58.708 ;
			RECT	194.615 58.644 194.647 58.708 ;
			RECT	194.783 58.644 194.815 58.708 ;
			RECT	194.951 58.644 194.983 58.708 ;
			RECT	195.119 58.644 195.151 58.708 ;
			RECT	195.287 58.644 195.319 58.708 ;
			RECT	195.455 58.644 195.487 58.708 ;
			RECT	195.623 58.644 195.655 58.708 ;
			RECT	195.791 58.644 195.823 58.708 ;
			RECT	195.959 58.644 195.991 58.708 ;
			RECT	196.127 58.644 196.159 58.708 ;
			RECT	196.295 58.644 196.327 58.708 ;
			RECT	196.463 58.644 196.495 58.708 ;
			RECT	196.631 58.644 196.663 58.708 ;
			RECT	196.799 58.644 196.831 58.708 ;
			RECT	196.967 58.644 196.999 58.708 ;
			RECT	197.135 58.644 197.167 58.708 ;
			RECT	197.303 58.644 197.335 58.708 ;
			RECT	197.471 58.644 197.503 58.708 ;
			RECT	197.639 58.644 197.671 58.708 ;
			RECT	197.807 58.644 197.839 58.708 ;
			RECT	197.975 58.644 198.007 58.708 ;
			RECT	198.143 58.644 198.175 58.708 ;
			RECT	198.311 58.644 198.343 58.708 ;
			RECT	198.479 58.644 198.511 58.708 ;
			RECT	198.647 58.644 198.679 58.708 ;
			RECT	198.815 58.644 198.847 58.708 ;
			RECT	198.983 58.644 199.015 58.708 ;
			RECT	199.151 58.644 199.183 58.708 ;
			RECT	199.319 58.644 199.351 58.708 ;
			RECT	199.487 58.644 199.519 58.708 ;
			RECT	199.655 58.644 199.687 58.708 ;
			RECT	199.823 58.644 199.855 58.708 ;
			RECT	199.991 58.644 200.023 58.708 ;
			RECT	200.121 58.66 200.153 58.692 ;
			RECT	200.243 58.655 200.275 58.687 ;
			RECT	200.373 58.644 200.405 58.708 ;
			RECT	200.9 58.644 200.932 58.708 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 56.696 201.665 56.816 ;
			LAYER	J3 ;
			RECT	0.755 56.724 0.787 56.788 ;
			RECT	1.645 56.724 1.709 56.788 ;
			RECT	2.323 56.724 2.387 56.788 ;
			RECT	3.438 56.724 3.47 56.788 ;
			RECT	3.585 56.724 3.617 56.788 ;
			RECT	4.195 56.724 4.227 56.788 ;
			RECT	4.72 56.724 4.752 56.788 ;
			RECT	4.944 56.724 5.008 56.788 ;
			RECT	5.267 56.724 5.299 56.788 ;
			RECT	5.797 56.724 5.829 56.788 ;
			RECT	5.927 56.735 5.959 56.767 ;
			RECT	6.049 56.74 6.081 56.772 ;
			RECT	6.179 56.724 6.211 56.788 ;
			RECT	6.347 56.724 6.379 56.788 ;
			RECT	6.515 56.724 6.547 56.788 ;
			RECT	6.683 56.724 6.715 56.788 ;
			RECT	6.851 56.724 6.883 56.788 ;
			RECT	7.019 56.724 7.051 56.788 ;
			RECT	7.187 56.724 7.219 56.788 ;
			RECT	7.355 56.724 7.387 56.788 ;
			RECT	7.523 56.724 7.555 56.788 ;
			RECT	7.691 56.724 7.723 56.788 ;
			RECT	7.859 56.724 7.891 56.788 ;
			RECT	8.027 56.724 8.059 56.788 ;
			RECT	8.195 56.724 8.227 56.788 ;
			RECT	8.363 56.724 8.395 56.788 ;
			RECT	8.531 56.724 8.563 56.788 ;
			RECT	8.699 56.724 8.731 56.788 ;
			RECT	8.867 56.724 8.899 56.788 ;
			RECT	9.035 56.724 9.067 56.788 ;
			RECT	9.203 56.724 9.235 56.788 ;
			RECT	9.371 56.724 9.403 56.788 ;
			RECT	9.539 56.724 9.571 56.788 ;
			RECT	9.707 56.724 9.739 56.788 ;
			RECT	9.875 56.724 9.907 56.788 ;
			RECT	10.043 56.724 10.075 56.788 ;
			RECT	10.211 56.724 10.243 56.788 ;
			RECT	10.379 56.724 10.411 56.788 ;
			RECT	10.547 56.724 10.579 56.788 ;
			RECT	10.715 56.724 10.747 56.788 ;
			RECT	10.883 56.724 10.915 56.788 ;
			RECT	11.051 56.724 11.083 56.788 ;
			RECT	11.219 56.724 11.251 56.788 ;
			RECT	11.387 56.724 11.419 56.788 ;
			RECT	11.555 56.724 11.587 56.788 ;
			RECT	11.723 56.724 11.755 56.788 ;
			RECT	11.891 56.724 11.923 56.788 ;
			RECT	12.059 56.724 12.091 56.788 ;
			RECT	12.227 56.724 12.259 56.788 ;
			RECT	12.395 56.724 12.427 56.788 ;
			RECT	12.563 56.724 12.595 56.788 ;
			RECT	12.731 56.724 12.763 56.788 ;
			RECT	12.899 56.724 12.931 56.788 ;
			RECT	13.067 56.724 13.099 56.788 ;
			RECT	13.235 56.724 13.267 56.788 ;
			RECT	13.403 56.724 13.435 56.788 ;
			RECT	13.571 56.724 13.603 56.788 ;
			RECT	13.739 56.724 13.771 56.788 ;
			RECT	13.907 56.724 13.939 56.788 ;
			RECT	14.075 56.724 14.107 56.788 ;
			RECT	14.243 56.724 14.275 56.788 ;
			RECT	14.411 56.724 14.443 56.788 ;
			RECT	14.579 56.724 14.611 56.788 ;
			RECT	14.747 56.724 14.779 56.788 ;
			RECT	14.915 56.724 14.947 56.788 ;
			RECT	15.083 56.724 15.115 56.788 ;
			RECT	15.251 56.724 15.283 56.788 ;
			RECT	15.419 56.724 15.451 56.788 ;
			RECT	15.587 56.724 15.619 56.788 ;
			RECT	15.755 56.724 15.787 56.788 ;
			RECT	15.923 56.724 15.955 56.788 ;
			RECT	16.091 56.724 16.123 56.788 ;
			RECT	16.259 56.724 16.291 56.788 ;
			RECT	16.427 56.724 16.459 56.788 ;
			RECT	16.595 56.724 16.627 56.788 ;
			RECT	16.763 56.724 16.795 56.788 ;
			RECT	16.931 56.724 16.963 56.788 ;
			RECT	17.099 56.724 17.131 56.788 ;
			RECT	17.267 56.724 17.299 56.788 ;
			RECT	17.435 56.724 17.467 56.788 ;
			RECT	17.603 56.724 17.635 56.788 ;
			RECT	17.771 56.724 17.803 56.788 ;
			RECT	17.939 56.724 17.971 56.788 ;
			RECT	18.107 56.724 18.139 56.788 ;
			RECT	18.275 56.724 18.307 56.788 ;
			RECT	18.443 56.724 18.475 56.788 ;
			RECT	18.611 56.724 18.643 56.788 ;
			RECT	18.779 56.724 18.811 56.788 ;
			RECT	18.947 56.724 18.979 56.788 ;
			RECT	19.115 56.724 19.147 56.788 ;
			RECT	19.283 56.724 19.315 56.788 ;
			RECT	19.451 56.724 19.483 56.788 ;
			RECT	19.619 56.724 19.651 56.788 ;
			RECT	19.787 56.724 19.819 56.788 ;
			RECT	19.955 56.724 19.987 56.788 ;
			RECT	20.123 56.724 20.155 56.788 ;
			RECT	20.291 56.724 20.323 56.788 ;
			RECT	20.459 56.724 20.491 56.788 ;
			RECT	20.627 56.724 20.659 56.788 ;
			RECT	20.795 56.724 20.827 56.788 ;
			RECT	20.963 56.724 20.995 56.788 ;
			RECT	21.131 56.724 21.163 56.788 ;
			RECT	21.299 56.724 21.331 56.788 ;
			RECT	21.467 56.724 21.499 56.788 ;
			RECT	21.635 56.724 21.667 56.788 ;
			RECT	21.803 56.724 21.835 56.788 ;
			RECT	21.971 56.724 22.003 56.788 ;
			RECT	22.139 56.724 22.171 56.788 ;
			RECT	22.307 56.724 22.339 56.788 ;
			RECT	22.475 56.724 22.507 56.788 ;
			RECT	22.643 56.724 22.675 56.788 ;
			RECT	22.811 56.724 22.843 56.788 ;
			RECT	22.979 56.724 23.011 56.788 ;
			RECT	23.147 56.724 23.179 56.788 ;
			RECT	23.315 56.724 23.347 56.788 ;
			RECT	23.483 56.724 23.515 56.788 ;
			RECT	23.651 56.724 23.683 56.788 ;
			RECT	23.819 56.724 23.851 56.788 ;
			RECT	23.987 56.724 24.019 56.788 ;
			RECT	24.155 56.724 24.187 56.788 ;
			RECT	24.323 56.724 24.355 56.788 ;
			RECT	24.491 56.724 24.523 56.788 ;
			RECT	24.659 56.724 24.691 56.788 ;
			RECT	24.827 56.724 24.859 56.788 ;
			RECT	24.995 56.724 25.027 56.788 ;
			RECT	25.163 56.724 25.195 56.788 ;
			RECT	25.331 56.724 25.363 56.788 ;
			RECT	25.499 56.724 25.531 56.788 ;
			RECT	25.667 56.724 25.699 56.788 ;
			RECT	25.835 56.724 25.867 56.788 ;
			RECT	26.003 56.724 26.035 56.788 ;
			RECT	26.171 56.724 26.203 56.788 ;
			RECT	26.339 56.724 26.371 56.788 ;
			RECT	26.507 56.724 26.539 56.788 ;
			RECT	26.675 56.724 26.707 56.788 ;
			RECT	26.843 56.724 26.875 56.788 ;
			RECT	27.011 56.724 27.043 56.788 ;
			RECT	27.179 56.724 27.211 56.788 ;
			RECT	27.347 56.724 27.379 56.788 ;
			RECT	27.515 56.724 27.547 56.788 ;
			RECT	27.683 56.724 27.715 56.788 ;
			RECT	27.851 56.724 27.883 56.788 ;
			RECT	28.019 56.724 28.051 56.788 ;
			RECT	28.187 56.724 28.219 56.788 ;
			RECT	28.355 56.724 28.387 56.788 ;
			RECT	28.523 56.724 28.555 56.788 ;
			RECT	28.691 56.724 28.723 56.788 ;
			RECT	28.859 56.724 28.891 56.788 ;
			RECT	29.027 56.724 29.059 56.788 ;
			RECT	29.195 56.724 29.227 56.788 ;
			RECT	29.363 56.724 29.395 56.788 ;
			RECT	29.531 56.724 29.563 56.788 ;
			RECT	29.699 56.724 29.731 56.788 ;
			RECT	29.867 56.724 29.899 56.788 ;
			RECT	30.035 56.724 30.067 56.788 ;
			RECT	30.203 56.724 30.235 56.788 ;
			RECT	30.371 56.724 30.403 56.788 ;
			RECT	30.539 56.724 30.571 56.788 ;
			RECT	30.707 56.724 30.739 56.788 ;
			RECT	30.875 56.724 30.907 56.788 ;
			RECT	31.043 56.724 31.075 56.788 ;
			RECT	31.211 56.724 31.243 56.788 ;
			RECT	31.379 56.724 31.411 56.788 ;
			RECT	31.547 56.724 31.579 56.788 ;
			RECT	31.715 56.724 31.747 56.788 ;
			RECT	31.883 56.724 31.915 56.788 ;
			RECT	32.051 56.724 32.083 56.788 ;
			RECT	32.219 56.724 32.251 56.788 ;
			RECT	32.387 56.724 32.419 56.788 ;
			RECT	32.555 56.724 32.587 56.788 ;
			RECT	32.723 56.724 32.755 56.788 ;
			RECT	32.891 56.724 32.923 56.788 ;
			RECT	33.059 56.724 33.091 56.788 ;
			RECT	33.227 56.724 33.259 56.788 ;
			RECT	33.395 56.724 33.427 56.788 ;
			RECT	33.563 56.724 33.595 56.788 ;
			RECT	33.731 56.724 33.763 56.788 ;
			RECT	33.899 56.724 33.931 56.788 ;
			RECT	34.067 56.724 34.099 56.788 ;
			RECT	34.235 56.724 34.267 56.788 ;
			RECT	34.403 56.724 34.435 56.788 ;
			RECT	34.571 56.724 34.603 56.788 ;
			RECT	34.739 56.724 34.771 56.788 ;
			RECT	34.907 56.724 34.939 56.788 ;
			RECT	35.075 56.724 35.107 56.788 ;
			RECT	35.243 56.724 35.275 56.788 ;
			RECT	35.411 56.724 35.443 56.788 ;
			RECT	35.579 56.724 35.611 56.788 ;
			RECT	35.747 56.724 35.779 56.788 ;
			RECT	35.915 56.724 35.947 56.788 ;
			RECT	36.083 56.724 36.115 56.788 ;
			RECT	36.251 56.724 36.283 56.788 ;
			RECT	36.419 56.724 36.451 56.788 ;
			RECT	36.587 56.724 36.619 56.788 ;
			RECT	36.755 56.724 36.787 56.788 ;
			RECT	36.923 56.724 36.955 56.788 ;
			RECT	37.091 56.724 37.123 56.788 ;
			RECT	37.259 56.724 37.291 56.788 ;
			RECT	37.427 56.724 37.459 56.788 ;
			RECT	37.595 56.724 37.627 56.788 ;
			RECT	37.763 56.724 37.795 56.788 ;
			RECT	37.931 56.724 37.963 56.788 ;
			RECT	38.099 56.724 38.131 56.788 ;
			RECT	38.267 56.724 38.299 56.788 ;
			RECT	38.435 56.724 38.467 56.788 ;
			RECT	38.603 56.724 38.635 56.788 ;
			RECT	38.771 56.724 38.803 56.788 ;
			RECT	38.939 56.724 38.971 56.788 ;
			RECT	39.107 56.724 39.139 56.788 ;
			RECT	39.275 56.724 39.307 56.788 ;
			RECT	39.443 56.724 39.475 56.788 ;
			RECT	39.611 56.724 39.643 56.788 ;
			RECT	39.779 56.724 39.811 56.788 ;
			RECT	39.947 56.724 39.979 56.788 ;
			RECT	40.115 56.724 40.147 56.788 ;
			RECT	40.283 56.724 40.315 56.788 ;
			RECT	40.451 56.724 40.483 56.788 ;
			RECT	40.619 56.724 40.651 56.788 ;
			RECT	40.787 56.724 40.819 56.788 ;
			RECT	40.955 56.724 40.987 56.788 ;
			RECT	41.123 56.724 41.155 56.788 ;
			RECT	41.291 56.724 41.323 56.788 ;
			RECT	41.459 56.724 41.491 56.788 ;
			RECT	41.627 56.724 41.659 56.788 ;
			RECT	41.795 56.724 41.827 56.788 ;
			RECT	41.963 56.724 41.995 56.788 ;
			RECT	42.131 56.724 42.163 56.788 ;
			RECT	42.299 56.724 42.331 56.788 ;
			RECT	42.467 56.724 42.499 56.788 ;
			RECT	42.635 56.724 42.667 56.788 ;
			RECT	42.803 56.724 42.835 56.788 ;
			RECT	42.971 56.724 43.003 56.788 ;
			RECT	43.139 56.724 43.171 56.788 ;
			RECT	43.307 56.724 43.339 56.788 ;
			RECT	43.475 56.724 43.507 56.788 ;
			RECT	43.643 56.724 43.675 56.788 ;
			RECT	43.811 56.724 43.843 56.788 ;
			RECT	43.979 56.724 44.011 56.788 ;
			RECT	44.147 56.724 44.179 56.788 ;
			RECT	44.315 56.724 44.347 56.788 ;
			RECT	44.483 56.724 44.515 56.788 ;
			RECT	44.651 56.724 44.683 56.788 ;
			RECT	44.819 56.724 44.851 56.788 ;
			RECT	44.987 56.724 45.019 56.788 ;
			RECT	45.155 56.724 45.187 56.788 ;
			RECT	45.323 56.724 45.355 56.788 ;
			RECT	45.491 56.724 45.523 56.788 ;
			RECT	45.659 56.724 45.691 56.788 ;
			RECT	45.827 56.724 45.859 56.788 ;
			RECT	45.995 56.724 46.027 56.788 ;
			RECT	46.163 56.724 46.195 56.788 ;
			RECT	46.331 56.724 46.363 56.788 ;
			RECT	46.499 56.724 46.531 56.788 ;
			RECT	46.667 56.724 46.699 56.788 ;
			RECT	46.835 56.724 46.867 56.788 ;
			RECT	47.003 56.724 47.035 56.788 ;
			RECT	47.171 56.724 47.203 56.788 ;
			RECT	47.339 56.724 47.371 56.788 ;
			RECT	47.507 56.724 47.539 56.788 ;
			RECT	47.675 56.724 47.707 56.788 ;
			RECT	47.843 56.724 47.875 56.788 ;
			RECT	48.011 56.724 48.043 56.788 ;
			RECT	48.179 56.724 48.211 56.788 ;
			RECT	48.347 56.724 48.379 56.788 ;
			RECT	48.515 56.724 48.547 56.788 ;
			RECT	48.683 56.724 48.715 56.788 ;
			RECT	48.851 56.724 48.883 56.788 ;
			RECT	49.019 56.724 49.051 56.788 ;
			RECT	49.187 56.724 49.219 56.788 ;
			RECT	49.318 56.74 49.35 56.772 ;
			RECT	49.439 56.74 49.471 56.772 ;
			RECT	49.569 56.724 49.601 56.788 ;
			RECT	51.881 56.724 51.913 56.788 ;
			RECT	53.132 56.724 53.196 56.788 ;
			RECT	53.812 56.724 53.844 56.788 ;
			RECT	54.251 56.724 54.283 56.788 ;
			RECT	55.562 56.724 55.626 56.788 ;
			RECT	58.603 56.724 58.635 56.788 ;
			RECT	58.733 56.74 58.765 56.772 ;
			RECT	58.854 56.74 58.886 56.772 ;
			RECT	58.985 56.724 59.017 56.788 ;
			RECT	59.153 56.724 59.185 56.788 ;
			RECT	59.321 56.724 59.353 56.788 ;
			RECT	59.489 56.724 59.521 56.788 ;
			RECT	59.657 56.724 59.689 56.788 ;
			RECT	59.825 56.724 59.857 56.788 ;
			RECT	59.993 56.724 60.025 56.788 ;
			RECT	60.161 56.724 60.193 56.788 ;
			RECT	60.329 56.724 60.361 56.788 ;
			RECT	60.497 56.724 60.529 56.788 ;
			RECT	60.665 56.724 60.697 56.788 ;
			RECT	60.833 56.724 60.865 56.788 ;
			RECT	61.001 56.724 61.033 56.788 ;
			RECT	61.169 56.724 61.201 56.788 ;
			RECT	61.337 56.724 61.369 56.788 ;
			RECT	61.505 56.724 61.537 56.788 ;
			RECT	61.673 56.724 61.705 56.788 ;
			RECT	61.841 56.724 61.873 56.788 ;
			RECT	62.009 56.724 62.041 56.788 ;
			RECT	62.177 56.724 62.209 56.788 ;
			RECT	62.345 56.724 62.377 56.788 ;
			RECT	62.513 56.724 62.545 56.788 ;
			RECT	62.681 56.724 62.713 56.788 ;
			RECT	62.849 56.724 62.881 56.788 ;
			RECT	63.017 56.724 63.049 56.788 ;
			RECT	63.185 56.724 63.217 56.788 ;
			RECT	63.353 56.724 63.385 56.788 ;
			RECT	63.521 56.724 63.553 56.788 ;
			RECT	63.689 56.724 63.721 56.788 ;
			RECT	63.857 56.724 63.889 56.788 ;
			RECT	64.025 56.724 64.057 56.788 ;
			RECT	64.193 56.724 64.225 56.788 ;
			RECT	64.361 56.724 64.393 56.788 ;
			RECT	64.529 56.724 64.561 56.788 ;
			RECT	64.697 56.724 64.729 56.788 ;
			RECT	64.865 56.724 64.897 56.788 ;
			RECT	65.033 56.724 65.065 56.788 ;
			RECT	65.201 56.724 65.233 56.788 ;
			RECT	65.369 56.724 65.401 56.788 ;
			RECT	65.537 56.724 65.569 56.788 ;
			RECT	65.705 56.724 65.737 56.788 ;
			RECT	65.873 56.724 65.905 56.788 ;
			RECT	66.041 56.724 66.073 56.788 ;
			RECT	66.209 56.724 66.241 56.788 ;
			RECT	66.377 56.724 66.409 56.788 ;
			RECT	66.545 56.724 66.577 56.788 ;
			RECT	66.713 56.724 66.745 56.788 ;
			RECT	66.881 56.724 66.913 56.788 ;
			RECT	67.049 56.724 67.081 56.788 ;
			RECT	67.217 56.724 67.249 56.788 ;
			RECT	67.385 56.724 67.417 56.788 ;
			RECT	67.553 56.724 67.585 56.788 ;
			RECT	67.721 56.724 67.753 56.788 ;
			RECT	67.889 56.724 67.921 56.788 ;
			RECT	68.057 56.724 68.089 56.788 ;
			RECT	68.225 56.724 68.257 56.788 ;
			RECT	68.393 56.724 68.425 56.788 ;
			RECT	68.561 56.724 68.593 56.788 ;
			RECT	68.729 56.724 68.761 56.788 ;
			RECT	68.897 56.724 68.929 56.788 ;
			RECT	69.065 56.724 69.097 56.788 ;
			RECT	69.233 56.724 69.265 56.788 ;
			RECT	69.401 56.724 69.433 56.788 ;
			RECT	69.569 56.724 69.601 56.788 ;
			RECT	69.737 56.724 69.769 56.788 ;
			RECT	69.905 56.724 69.937 56.788 ;
			RECT	70.073 56.724 70.105 56.788 ;
			RECT	70.241 56.724 70.273 56.788 ;
			RECT	70.409 56.724 70.441 56.788 ;
			RECT	70.577 56.724 70.609 56.788 ;
			RECT	70.745 56.724 70.777 56.788 ;
			RECT	70.913 56.724 70.945 56.788 ;
			RECT	71.081 56.724 71.113 56.788 ;
			RECT	71.249 56.724 71.281 56.788 ;
			RECT	71.417 56.724 71.449 56.788 ;
			RECT	71.585 56.724 71.617 56.788 ;
			RECT	71.753 56.724 71.785 56.788 ;
			RECT	71.921 56.724 71.953 56.788 ;
			RECT	72.089 56.724 72.121 56.788 ;
			RECT	72.257 56.724 72.289 56.788 ;
			RECT	72.425 56.724 72.457 56.788 ;
			RECT	72.593 56.724 72.625 56.788 ;
			RECT	72.761 56.724 72.793 56.788 ;
			RECT	72.929 56.724 72.961 56.788 ;
			RECT	73.097 56.724 73.129 56.788 ;
			RECT	73.265 56.724 73.297 56.788 ;
			RECT	73.433 56.724 73.465 56.788 ;
			RECT	73.601 56.724 73.633 56.788 ;
			RECT	73.769 56.724 73.801 56.788 ;
			RECT	73.937 56.724 73.969 56.788 ;
			RECT	74.105 56.724 74.137 56.788 ;
			RECT	74.273 56.724 74.305 56.788 ;
			RECT	74.441 56.724 74.473 56.788 ;
			RECT	74.609 56.724 74.641 56.788 ;
			RECT	74.777 56.724 74.809 56.788 ;
			RECT	74.945 56.724 74.977 56.788 ;
			RECT	75.113 56.724 75.145 56.788 ;
			RECT	75.281 56.724 75.313 56.788 ;
			RECT	75.449 56.724 75.481 56.788 ;
			RECT	75.617 56.724 75.649 56.788 ;
			RECT	75.785 56.724 75.817 56.788 ;
			RECT	75.953 56.724 75.985 56.788 ;
			RECT	76.121 56.724 76.153 56.788 ;
			RECT	76.289 56.724 76.321 56.788 ;
			RECT	76.457 56.724 76.489 56.788 ;
			RECT	76.625 56.724 76.657 56.788 ;
			RECT	76.793 56.724 76.825 56.788 ;
			RECT	76.961 56.724 76.993 56.788 ;
			RECT	77.129 56.724 77.161 56.788 ;
			RECT	77.297 56.724 77.329 56.788 ;
			RECT	77.465 56.724 77.497 56.788 ;
			RECT	77.633 56.724 77.665 56.788 ;
			RECT	77.801 56.724 77.833 56.788 ;
			RECT	77.969 56.724 78.001 56.788 ;
			RECT	78.137 56.724 78.169 56.788 ;
			RECT	78.305 56.724 78.337 56.788 ;
			RECT	78.473 56.724 78.505 56.788 ;
			RECT	78.641 56.724 78.673 56.788 ;
			RECT	78.809 56.724 78.841 56.788 ;
			RECT	78.977 56.724 79.009 56.788 ;
			RECT	79.145 56.724 79.177 56.788 ;
			RECT	79.313 56.724 79.345 56.788 ;
			RECT	79.481 56.724 79.513 56.788 ;
			RECT	79.649 56.724 79.681 56.788 ;
			RECT	79.817 56.724 79.849 56.788 ;
			RECT	79.985 56.724 80.017 56.788 ;
			RECT	80.153 56.724 80.185 56.788 ;
			RECT	80.321 56.724 80.353 56.788 ;
			RECT	80.489 56.724 80.521 56.788 ;
			RECT	80.657 56.724 80.689 56.788 ;
			RECT	80.825 56.724 80.857 56.788 ;
			RECT	80.993 56.724 81.025 56.788 ;
			RECT	81.161 56.724 81.193 56.788 ;
			RECT	81.329 56.724 81.361 56.788 ;
			RECT	81.497 56.724 81.529 56.788 ;
			RECT	81.665 56.724 81.697 56.788 ;
			RECT	81.833 56.724 81.865 56.788 ;
			RECT	82.001 56.724 82.033 56.788 ;
			RECT	82.169 56.724 82.201 56.788 ;
			RECT	82.337 56.724 82.369 56.788 ;
			RECT	82.505 56.724 82.537 56.788 ;
			RECT	82.673 56.724 82.705 56.788 ;
			RECT	82.841 56.724 82.873 56.788 ;
			RECT	83.009 56.724 83.041 56.788 ;
			RECT	83.177 56.724 83.209 56.788 ;
			RECT	83.345 56.724 83.377 56.788 ;
			RECT	83.513 56.724 83.545 56.788 ;
			RECT	83.681 56.724 83.713 56.788 ;
			RECT	83.849 56.724 83.881 56.788 ;
			RECT	84.017 56.724 84.049 56.788 ;
			RECT	84.185 56.724 84.217 56.788 ;
			RECT	84.353 56.724 84.385 56.788 ;
			RECT	84.521 56.724 84.553 56.788 ;
			RECT	84.689 56.724 84.721 56.788 ;
			RECT	84.857 56.724 84.889 56.788 ;
			RECT	85.025 56.724 85.057 56.788 ;
			RECT	85.193 56.724 85.225 56.788 ;
			RECT	85.361 56.724 85.393 56.788 ;
			RECT	85.529 56.724 85.561 56.788 ;
			RECT	85.697 56.724 85.729 56.788 ;
			RECT	85.865 56.724 85.897 56.788 ;
			RECT	86.033 56.724 86.065 56.788 ;
			RECT	86.201 56.724 86.233 56.788 ;
			RECT	86.369 56.724 86.401 56.788 ;
			RECT	86.537 56.724 86.569 56.788 ;
			RECT	86.705 56.724 86.737 56.788 ;
			RECT	86.873 56.724 86.905 56.788 ;
			RECT	87.041 56.724 87.073 56.788 ;
			RECT	87.209 56.724 87.241 56.788 ;
			RECT	87.377 56.724 87.409 56.788 ;
			RECT	87.545 56.724 87.577 56.788 ;
			RECT	87.713 56.724 87.745 56.788 ;
			RECT	87.881 56.724 87.913 56.788 ;
			RECT	88.049 56.724 88.081 56.788 ;
			RECT	88.217 56.724 88.249 56.788 ;
			RECT	88.385 56.724 88.417 56.788 ;
			RECT	88.553 56.724 88.585 56.788 ;
			RECT	88.721 56.724 88.753 56.788 ;
			RECT	88.889 56.724 88.921 56.788 ;
			RECT	89.057 56.724 89.089 56.788 ;
			RECT	89.225 56.724 89.257 56.788 ;
			RECT	89.393 56.724 89.425 56.788 ;
			RECT	89.561 56.724 89.593 56.788 ;
			RECT	89.729 56.724 89.761 56.788 ;
			RECT	89.897 56.724 89.929 56.788 ;
			RECT	90.065 56.724 90.097 56.788 ;
			RECT	90.233 56.724 90.265 56.788 ;
			RECT	90.401 56.724 90.433 56.788 ;
			RECT	90.569 56.724 90.601 56.788 ;
			RECT	90.737 56.724 90.769 56.788 ;
			RECT	90.905 56.724 90.937 56.788 ;
			RECT	91.073 56.724 91.105 56.788 ;
			RECT	91.241 56.724 91.273 56.788 ;
			RECT	91.409 56.724 91.441 56.788 ;
			RECT	91.577 56.724 91.609 56.788 ;
			RECT	91.745 56.724 91.777 56.788 ;
			RECT	91.913 56.724 91.945 56.788 ;
			RECT	92.081 56.724 92.113 56.788 ;
			RECT	92.249 56.724 92.281 56.788 ;
			RECT	92.417 56.724 92.449 56.788 ;
			RECT	92.585 56.724 92.617 56.788 ;
			RECT	92.753 56.724 92.785 56.788 ;
			RECT	92.921 56.724 92.953 56.788 ;
			RECT	93.089 56.724 93.121 56.788 ;
			RECT	93.257 56.724 93.289 56.788 ;
			RECT	93.425 56.724 93.457 56.788 ;
			RECT	93.593 56.724 93.625 56.788 ;
			RECT	93.761 56.724 93.793 56.788 ;
			RECT	93.929 56.724 93.961 56.788 ;
			RECT	94.097 56.724 94.129 56.788 ;
			RECT	94.265 56.724 94.297 56.788 ;
			RECT	94.433 56.724 94.465 56.788 ;
			RECT	94.601 56.724 94.633 56.788 ;
			RECT	94.769 56.724 94.801 56.788 ;
			RECT	94.937 56.724 94.969 56.788 ;
			RECT	95.105 56.724 95.137 56.788 ;
			RECT	95.273 56.724 95.305 56.788 ;
			RECT	95.441 56.724 95.473 56.788 ;
			RECT	95.609 56.724 95.641 56.788 ;
			RECT	95.777 56.724 95.809 56.788 ;
			RECT	95.945 56.724 95.977 56.788 ;
			RECT	96.113 56.724 96.145 56.788 ;
			RECT	96.281 56.724 96.313 56.788 ;
			RECT	96.449 56.724 96.481 56.788 ;
			RECT	96.617 56.724 96.649 56.788 ;
			RECT	96.785 56.724 96.817 56.788 ;
			RECT	96.953 56.724 96.985 56.788 ;
			RECT	97.121 56.724 97.153 56.788 ;
			RECT	97.289 56.724 97.321 56.788 ;
			RECT	97.457 56.724 97.489 56.788 ;
			RECT	97.625 56.724 97.657 56.788 ;
			RECT	97.793 56.724 97.825 56.788 ;
			RECT	97.961 56.724 97.993 56.788 ;
			RECT	98.129 56.724 98.161 56.788 ;
			RECT	98.297 56.724 98.329 56.788 ;
			RECT	98.465 56.724 98.497 56.788 ;
			RECT	98.633 56.724 98.665 56.788 ;
			RECT	98.801 56.724 98.833 56.788 ;
			RECT	98.969 56.724 99.001 56.788 ;
			RECT	99.137 56.724 99.169 56.788 ;
			RECT	99.305 56.724 99.337 56.788 ;
			RECT	99.473 56.724 99.505 56.788 ;
			RECT	99.641 56.724 99.673 56.788 ;
			RECT	99.809 56.724 99.841 56.788 ;
			RECT	99.977 56.724 100.009 56.788 ;
			RECT	100.145 56.724 100.177 56.788 ;
			RECT	100.313 56.724 100.345 56.788 ;
			RECT	100.481 56.724 100.513 56.788 ;
			RECT	100.649 56.724 100.681 56.788 ;
			RECT	100.817 56.724 100.849 56.788 ;
			RECT	100.985 56.724 101.017 56.788 ;
			RECT	101.153 56.724 101.185 56.788 ;
			RECT	101.321 56.724 101.353 56.788 ;
			RECT	101.489 56.724 101.521 56.788 ;
			RECT	101.657 56.724 101.689 56.788 ;
			RECT	101.825 56.724 101.857 56.788 ;
			RECT	101.993 56.724 102.025 56.788 ;
			RECT	102.123 56.74 102.155 56.772 ;
			RECT	102.245 56.735 102.277 56.767 ;
			RECT	102.375 56.724 102.407 56.788 ;
			RECT	103.795 56.724 103.827 56.788 ;
			RECT	103.925 56.735 103.957 56.767 ;
			RECT	104.047 56.74 104.079 56.772 ;
			RECT	104.177 56.724 104.209 56.788 ;
			RECT	104.345 56.724 104.377 56.788 ;
			RECT	104.513 56.724 104.545 56.788 ;
			RECT	104.681 56.724 104.713 56.788 ;
			RECT	104.849 56.724 104.881 56.788 ;
			RECT	105.017 56.724 105.049 56.788 ;
			RECT	105.185 56.724 105.217 56.788 ;
			RECT	105.353 56.724 105.385 56.788 ;
			RECT	105.521 56.724 105.553 56.788 ;
			RECT	105.689 56.724 105.721 56.788 ;
			RECT	105.857 56.724 105.889 56.788 ;
			RECT	106.025 56.724 106.057 56.788 ;
			RECT	106.193 56.724 106.225 56.788 ;
			RECT	106.361 56.724 106.393 56.788 ;
			RECT	106.529 56.724 106.561 56.788 ;
			RECT	106.697 56.724 106.729 56.788 ;
			RECT	106.865 56.724 106.897 56.788 ;
			RECT	107.033 56.724 107.065 56.788 ;
			RECT	107.201 56.724 107.233 56.788 ;
			RECT	107.369 56.724 107.401 56.788 ;
			RECT	107.537 56.724 107.569 56.788 ;
			RECT	107.705 56.724 107.737 56.788 ;
			RECT	107.873 56.724 107.905 56.788 ;
			RECT	108.041 56.724 108.073 56.788 ;
			RECT	108.209 56.724 108.241 56.788 ;
			RECT	108.377 56.724 108.409 56.788 ;
			RECT	108.545 56.724 108.577 56.788 ;
			RECT	108.713 56.724 108.745 56.788 ;
			RECT	108.881 56.724 108.913 56.788 ;
			RECT	109.049 56.724 109.081 56.788 ;
			RECT	109.217 56.724 109.249 56.788 ;
			RECT	109.385 56.724 109.417 56.788 ;
			RECT	109.553 56.724 109.585 56.788 ;
			RECT	109.721 56.724 109.753 56.788 ;
			RECT	109.889 56.724 109.921 56.788 ;
			RECT	110.057 56.724 110.089 56.788 ;
			RECT	110.225 56.724 110.257 56.788 ;
			RECT	110.393 56.724 110.425 56.788 ;
			RECT	110.561 56.724 110.593 56.788 ;
			RECT	110.729 56.724 110.761 56.788 ;
			RECT	110.897 56.724 110.929 56.788 ;
			RECT	111.065 56.724 111.097 56.788 ;
			RECT	111.233 56.724 111.265 56.788 ;
			RECT	111.401 56.724 111.433 56.788 ;
			RECT	111.569 56.724 111.601 56.788 ;
			RECT	111.737 56.724 111.769 56.788 ;
			RECT	111.905 56.724 111.937 56.788 ;
			RECT	112.073 56.724 112.105 56.788 ;
			RECT	112.241 56.724 112.273 56.788 ;
			RECT	112.409 56.724 112.441 56.788 ;
			RECT	112.577 56.724 112.609 56.788 ;
			RECT	112.745 56.724 112.777 56.788 ;
			RECT	112.913 56.724 112.945 56.788 ;
			RECT	113.081 56.724 113.113 56.788 ;
			RECT	113.249 56.724 113.281 56.788 ;
			RECT	113.417 56.724 113.449 56.788 ;
			RECT	113.585 56.724 113.617 56.788 ;
			RECT	113.753 56.724 113.785 56.788 ;
			RECT	113.921 56.724 113.953 56.788 ;
			RECT	114.089 56.724 114.121 56.788 ;
			RECT	114.257 56.724 114.289 56.788 ;
			RECT	114.425 56.724 114.457 56.788 ;
			RECT	114.593 56.724 114.625 56.788 ;
			RECT	114.761 56.724 114.793 56.788 ;
			RECT	114.929 56.724 114.961 56.788 ;
			RECT	115.097 56.724 115.129 56.788 ;
			RECT	115.265 56.724 115.297 56.788 ;
			RECT	115.433 56.724 115.465 56.788 ;
			RECT	115.601 56.724 115.633 56.788 ;
			RECT	115.769 56.724 115.801 56.788 ;
			RECT	115.937 56.724 115.969 56.788 ;
			RECT	116.105 56.724 116.137 56.788 ;
			RECT	116.273 56.724 116.305 56.788 ;
			RECT	116.441 56.724 116.473 56.788 ;
			RECT	116.609 56.724 116.641 56.788 ;
			RECT	116.777 56.724 116.809 56.788 ;
			RECT	116.945 56.724 116.977 56.788 ;
			RECT	117.113 56.724 117.145 56.788 ;
			RECT	117.281 56.724 117.313 56.788 ;
			RECT	117.449 56.724 117.481 56.788 ;
			RECT	117.617 56.724 117.649 56.788 ;
			RECT	117.785 56.724 117.817 56.788 ;
			RECT	117.953 56.724 117.985 56.788 ;
			RECT	118.121 56.724 118.153 56.788 ;
			RECT	118.289 56.724 118.321 56.788 ;
			RECT	118.457 56.724 118.489 56.788 ;
			RECT	118.625 56.724 118.657 56.788 ;
			RECT	118.793 56.724 118.825 56.788 ;
			RECT	118.961 56.724 118.993 56.788 ;
			RECT	119.129 56.724 119.161 56.788 ;
			RECT	119.297 56.724 119.329 56.788 ;
			RECT	119.465 56.724 119.497 56.788 ;
			RECT	119.633 56.724 119.665 56.788 ;
			RECT	119.801 56.724 119.833 56.788 ;
			RECT	119.969 56.724 120.001 56.788 ;
			RECT	120.137 56.724 120.169 56.788 ;
			RECT	120.305 56.724 120.337 56.788 ;
			RECT	120.473 56.724 120.505 56.788 ;
			RECT	120.641 56.724 120.673 56.788 ;
			RECT	120.809 56.724 120.841 56.788 ;
			RECT	120.977 56.724 121.009 56.788 ;
			RECT	121.145 56.724 121.177 56.788 ;
			RECT	121.313 56.724 121.345 56.788 ;
			RECT	121.481 56.724 121.513 56.788 ;
			RECT	121.649 56.724 121.681 56.788 ;
			RECT	121.817 56.724 121.849 56.788 ;
			RECT	121.985 56.724 122.017 56.788 ;
			RECT	122.153 56.724 122.185 56.788 ;
			RECT	122.321 56.724 122.353 56.788 ;
			RECT	122.489 56.724 122.521 56.788 ;
			RECT	122.657 56.724 122.689 56.788 ;
			RECT	122.825 56.724 122.857 56.788 ;
			RECT	122.993 56.724 123.025 56.788 ;
			RECT	123.161 56.724 123.193 56.788 ;
			RECT	123.329 56.724 123.361 56.788 ;
			RECT	123.497 56.724 123.529 56.788 ;
			RECT	123.665 56.724 123.697 56.788 ;
			RECT	123.833 56.724 123.865 56.788 ;
			RECT	124.001 56.724 124.033 56.788 ;
			RECT	124.169 56.724 124.201 56.788 ;
			RECT	124.337 56.724 124.369 56.788 ;
			RECT	124.505 56.724 124.537 56.788 ;
			RECT	124.673 56.724 124.705 56.788 ;
			RECT	124.841 56.724 124.873 56.788 ;
			RECT	125.009 56.724 125.041 56.788 ;
			RECT	125.177 56.724 125.209 56.788 ;
			RECT	125.345 56.724 125.377 56.788 ;
			RECT	125.513 56.724 125.545 56.788 ;
			RECT	125.681 56.724 125.713 56.788 ;
			RECT	125.849 56.724 125.881 56.788 ;
			RECT	126.017 56.724 126.049 56.788 ;
			RECT	126.185 56.724 126.217 56.788 ;
			RECT	126.353 56.724 126.385 56.788 ;
			RECT	126.521 56.724 126.553 56.788 ;
			RECT	126.689 56.724 126.721 56.788 ;
			RECT	126.857 56.724 126.889 56.788 ;
			RECT	127.025 56.724 127.057 56.788 ;
			RECT	127.193 56.724 127.225 56.788 ;
			RECT	127.361 56.724 127.393 56.788 ;
			RECT	127.529 56.724 127.561 56.788 ;
			RECT	127.697 56.724 127.729 56.788 ;
			RECT	127.865 56.724 127.897 56.788 ;
			RECT	128.033 56.724 128.065 56.788 ;
			RECT	128.201 56.724 128.233 56.788 ;
			RECT	128.369 56.724 128.401 56.788 ;
			RECT	128.537 56.724 128.569 56.788 ;
			RECT	128.705 56.724 128.737 56.788 ;
			RECT	128.873 56.724 128.905 56.788 ;
			RECT	129.041 56.724 129.073 56.788 ;
			RECT	129.209 56.724 129.241 56.788 ;
			RECT	129.377 56.724 129.409 56.788 ;
			RECT	129.545 56.724 129.577 56.788 ;
			RECT	129.713 56.724 129.745 56.788 ;
			RECT	129.881 56.724 129.913 56.788 ;
			RECT	130.049 56.724 130.081 56.788 ;
			RECT	130.217 56.724 130.249 56.788 ;
			RECT	130.385 56.724 130.417 56.788 ;
			RECT	130.553 56.724 130.585 56.788 ;
			RECT	130.721 56.724 130.753 56.788 ;
			RECT	130.889 56.724 130.921 56.788 ;
			RECT	131.057 56.724 131.089 56.788 ;
			RECT	131.225 56.724 131.257 56.788 ;
			RECT	131.393 56.724 131.425 56.788 ;
			RECT	131.561 56.724 131.593 56.788 ;
			RECT	131.729 56.724 131.761 56.788 ;
			RECT	131.897 56.724 131.929 56.788 ;
			RECT	132.065 56.724 132.097 56.788 ;
			RECT	132.233 56.724 132.265 56.788 ;
			RECT	132.401 56.724 132.433 56.788 ;
			RECT	132.569 56.724 132.601 56.788 ;
			RECT	132.737 56.724 132.769 56.788 ;
			RECT	132.905 56.724 132.937 56.788 ;
			RECT	133.073 56.724 133.105 56.788 ;
			RECT	133.241 56.724 133.273 56.788 ;
			RECT	133.409 56.724 133.441 56.788 ;
			RECT	133.577 56.724 133.609 56.788 ;
			RECT	133.745 56.724 133.777 56.788 ;
			RECT	133.913 56.724 133.945 56.788 ;
			RECT	134.081 56.724 134.113 56.788 ;
			RECT	134.249 56.724 134.281 56.788 ;
			RECT	134.417 56.724 134.449 56.788 ;
			RECT	134.585 56.724 134.617 56.788 ;
			RECT	134.753 56.724 134.785 56.788 ;
			RECT	134.921 56.724 134.953 56.788 ;
			RECT	135.089 56.724 135.121 56.788 ;
			RECT	135.257 56.724 135.289 56.788 ;
			RECT	135.425 56.724 135.457 56.788 ;
			RECT	135.593 56.724 135.625 56.788 ;
			RECT	135.761 56.724 135.793 56.788 ;
			RECT	135.929 56.724 135.961 56.788 ;
			RECT	136.097 56.724 136.129 56.788 ;
			RECT	136.265 56.724 136.297 56.788 ;
			RECT	136.433 56.724 136.465 56.788 ;
			RECT	136.601 56.724 136.633 56.788 ;
			RECT	136.769 56.724 136.801 56.788 ;
			RECT	136.937 56.724 136.969 56.788 ;
			RECT	137.105 56.724 137.137 56.788 ;
			RECT	137.273 56.724 137.305 56.788 ;
			RECT	137.441 56.724 137.473 56.788 ;
			RECT	137.609 56.724 137.641 56.788 ;
			RECT	137.777 56.724 137.809 56.788 ;
			RECT	137.945 56.724 137.977 56.788 ;
			RECT	138.113 56.724 138.145 56.788 ;
			RECT	138.281 56.724 138.313 56.788 ;
			RECT	138.449 56.724 138.481 56.788 ;
			RECT	138.617 56.724 138.649 56.788 ;
			RECT	138.785 56.724 138.817 56.788 ;
			RECT	138.953 56.724 138.985 56.788 ;
			RECT	139.121 56.724 139.153 56.788 ;
			RECT	139.289 56.724 139.321 56.788 ;
			RECT	139.457 56.724 139.489 56.788 ;
			RECT	139.625 56.724 139.657 56.788 ;
			RECT	139.793 56.724 139.825 56.788 ;
			RECT	139.961 56.724 139.993 56.788 ;
			RECT	140.129 56.724 140.161 56.788 ;
			RECT	140.297 56.724 140.329 56.788 ;
			RECT	140.465 56.724 140.497 56.788 ;
			RECT	140.633 56.724 140.665 56.788 ;
			RECT	140.801 56.724 140.833 56.788 ;
			RECT	140.969 56.724 141.001 56.788 ;
			RECT	141.137 56.724 141.169 56.788 ;
			RECT	141.305 56.724 141.337 56.788 ;
			RECT	141.473 56.724 141.505 56.788 ;
			RECT	141.641 56.724 141.673 56.788 ;
			RECT	141.809 56.724 141.841 56.788 ;
			RECT	141.977 56.724 142.009 56.788 ;
			RECT	142.145 56.724 142.177 56.788 ;
			RECT	142.313 56.724 142.345 56.788 ;
			RECT	142.481 56.724 142.513 56.788 ;
			RECT	142.649 56.724 142.681 56.788 ;
			RECT	142.817 56.724 142.849 56.788 ;
			RECT	142.985 56.724 143.017 56.788 ;
			RECT	143.153 56.724 143.185 56.788 ;
			RECT	143.321 56.724 143.353 56.788 ;
			RECT	143.489 56.724 143.521 56.788 ;
			RECT	143.657 56.724 143.689 56.788 ;
			RECT	143.825 56.724 143.857 56.788 ;
			RECT	143.993 56.724 144.025 56.788 ;
			RECT	144.161 56.724 144.193 56.788 ;
			RECT	144.329 56.724 144.361 56.788 ;
			RECT	144.497 56.724 144.529 56.788 ;
			RECT	144.665 56.724 144.697 56.788 ;
			RECT	144.833 56.724 144.865 56.788 ;
			RECT	145.001 56.724 145.033 56.788 ;
			RECT	145.169 56.724 145.201 56.788 ;
			RECT	145.337 56.724 145.369 56.788 ;
			RECT	145.505 56.724 145.537 56.788 ;
			RECT	145.673 56.724 145.705 56.788 ;
			RECT	145.841 56.724 145.873 56.788 ;
			RECT	146.009 56.724 146.041 56.788 ;
			RECT	146.177 56.724 146.209 56.788 ;
			RECT	146.345 56.724 146.377 56.788 ;
			RECT	146.513 56.724 146.545 56.788 ;
			RECT	146.681 56.724 146.713 56.788 ;
			RECT	146.849 56.724 146.881 56.788 ;
			RECT	147.017 56.724 147.049 56.788 ;
			RECT	147.185 56.724 147.217 56.788 ;
			RECT	147.316 56.74 147.348 56.772 ;
			RECT	147.437 56.74 147.469 56.772 ;
			RECT	147.567 56.724 147.599 56.788 ;
			RECT	149.879 56.724 149.911 56.788 ;
			RECT	151.13 56.724 151.194 56.788 ;
			RECT	151.81 56.724 151.842 56.788 ;
			RECT	152.249 56.724 152.281 56.788 ;
			RECT	153.56 56.724 153.624 56.788 ;
			RECT	156.601 56.724 156.633 56.788 ;
			RECT	156.731 56.74 156.763 56.772 ;
			RECT	156.852 56.74 156.884 56.772 ;
			RECT	156.983 56.724 157.015 56.788 ;
			RECT	157.151 56.724 157.183 56.788 ;
			RECT	157.319 56.724 157.351 56.788 ;
			RECT	157.487 56.724 157.519 56.788 ;
			RECT	157.655 56.724 157.687 56.788 ;
			RECT	157.823 56.724 157.855 56.788 ;
			RECT	157.991 56.724 158.023 56.788 ;
			RECT	158.159 56.724 158.191 56.788 ;
			RECT	158.327 56.724 158.359 56.788 ;
			RECT	158.495 56.724 158.527 56.788 ;
			RECT	158.663 56.724 158.695 56.788 ;
			RECT	158.831 56.724 158.863 56.788 ;
			RECT	158.999 56.724 159.031 56.788 ;
			RECT	159.167 56.724 159.199 56.788 ;
			RECT	159.335 56.724 159.367 56.788 ;
			RECT	159.503 56.724 159.535 56.788 ;
			RECT	159.671 56.724 159.703 56.788 ;
			RECT	159.839 56.724 159.871 56.788 ;
			RECT	160.007 56.724 160.039 56.788 ;
			RECT	160.175 56.724 160.207 56.788 ;
			RECT	160.343 56.724 160.375 56.788 ;
			RECT	160.511 56.724 160.543 56.788 ;
			RECT	160.679 56.724 160.711 56.788 ;
			RECT	160.847 56.724 160.879 56.788 ;
			RECT	161.015 56.724 161.047 56.788 ;
			RECT	161.183 56.724 161.215 56.788 ;
			RECT	161.351 56.724 161.383 56.788 ;
			RECT	161.519 56.724 161.551 56.788 ;
			RECT	161.687 56.724 161.719 56.788 ;
			RECT	161.855 56.724 161.887 56.788 ;
			RECT	162.023 56.724 162.055 56.788 ;
			RECT	162.191 56.724 162.223 56.788 ;
			RECT	162.359 56.724 162.391 56.788 ;
			RECT	162.527 56.724 162.559 56.788 ;
			RECT	162.695 56.724 162.727 56.788 ;
			RECT	162.863 56.724 162.895 56.788 ;
			RECT	163.031 56.724 163.063 56.788 ;
			RECT	163.199 56.724 163.231 56.788 ;
			RECT	163.367 56.724 163.399 56.788 ;
			RECT	163.535 56.724 163.567 56.788 ;
			RECT	163.703 56.724 163.735 56.788 ;
			RECT	163.871 56.724 163.903 56.788 ;
			RECT	164.039 56.724 164.071 56.788 ;
			RECT	164.207 56.724 164.239 56.788 ;
			RECT	164.375 56.724 164.407 56.788 ;
			RECT	164.543 56.724 164.575 56.788 ;
			RECT	164.711 56.724 164.743 56.788 ;
			RECT	164.879 56.724 164.911 56.788 ;
			RECT	165.047 56.724 165.079 56.788 ;
			RECT	165.215 56.724 165.247 56.788 ;
			RECT	165.383 56.724 165.415 56.788 ;
			RECT	165.551 56.724 165.583 56.788 ;
			RECT	165.719 56.724 165.751 56.788 ;
			RECT	165.887 56.724 165.919 56.788 ;
			RECT	166.055 56.724 166.087 56.788 ;
			RECT	166.223 56.724 166.255 56.788 ;
			RECT	166.391 56.724 166.423 56.788 ;
			RECT	166.559 56.724 166.591 56.788 ;
			RECT	166.727 56.724 166.759 56.788 ;
			RECT	166.895 56.724 166.927 56.788 ;
			RECT	167.063 56.724 167.095 56.788 ;
			RECT	167.231 56.724 167.263 56.788 ;
			RECT	167.399 56.724 167.431 56.788 ;
			RECT	167.567 56.724 167.599 56.788 ;
			RECT	167.735 56.724 167.767 56.788 ;
			RECT	167.903 56.724 167.935 56.788 ;
			RECT	168.071 56.724 168.103 56.788 ;
			RECT	168.239 56.724 168.271 56.788 ;
			RECT	168.407 56.724 168.439 56.788 ;
			RECT	168.575 56.724 168.607 56.788 ;
			RECT	168.743 56.724 168.775 56.788 ;
			RECT	168.911 56.724 168.943 56.788 ;
			RECT	169.079 56.724 169.111 56.788 ;
			RECT	169.247 56.724 169.279 56.788 ;
			RECT	169.415 56.724 169.447 56.788 ;
			RECT	169.583 56.724 169.615 56.788 ;
			RECT	169.751 56.724 169.783 56.788 ;
			RECT	169.919 56.724 169.951 56.788 ;
			RECT	170.087 56.724 170.119 56.788 ;
			RECT	170.255 56.724 170.287 56.788 ;
			RECT	170.423 56.724 170.455 56.788 ;
			RECT	170.591 56.724 170.623 56.788 ;
			RECT	170.759 56.724 170.791 56.788 ;
			RECT	170.927 56.724 170.959 56.788 ;
			RECT	171.095 56.724 171.127 56.788 ;
			RECT	171.263 56.724 171.295 56.788 ;
			RECT	171.431 56.724 171.463 56.788 ;
			RECT	171.599 56.724 171.631 56.788 ;
			RECT	171.767 56.724 171.799 56.788 ;
			RECT	171.935 56.724 171.967 56.788 ;
			RECT	172.103 56.724 172.135 56.788 ;
			RECT	172.271 56.724 172.303 56.788 ;
			RECT	172.439 56.724 172.471 56.788 ;
			RECT	172.607 56.724 172.639 56.788 ;
			RECT	172.775 56.724 172.807 56.788 ;
			RECT	172.943 56.724 172.975 56.788 ;
			RECT	173.111 56.724 173.143 56.788 ;
			RECT	173.279 56.724 173.311 56.788 ;
			RECT	173.447 56.724 173.479 56.788 ;
			RECT	173.615 56.724 173.647 56.788 ;
			RECT	173.783 56.724 173.815 56.788 ;
			RECT	173.951 56.724 173.983 56.788 ;
			RECT	174.119 56.724 174.151 56.788 ;
			RECT	174.287 56.724 174.319 56.788 ;
			RECT	174.455 56.724 174.487 56.788 ;
			RECT	174.623 56.724 174.655 56.788 ;
			RECT	174.791 56.724 174.823 56.788 ;
			RECT	174.959 56.724 174.991 56.788 ;
			RECT	175.127 56.724 175.159 56.788 ;
			RECT	175.295 56.724 175.327 56.788 ;
			RECT	175.463 56.724 175.495 56.788 ;
			RECT	175.631 56.724 175.663 56.788 ;
			RECT	175.799 56.724 175.831 56.788 ;
			RECT	175.967 56.724 175.999 56.788 ;
			RECT	176.135 56.724 176.167 56.788 ;
			RECT	176.303 56.724 176.335 56.788 ;
			RECT	176.471 56.724 176.503 56.788 ;
			RECT	176.639 56.724 176.671 56.788 ;
			RECT	176.807 56.724 176.839 56.788 ;
			RECT	176.975 56.724 177.007 56.788 ;
			RECT	177.143 56.724 177.175 56.788 ;
			RECT	177.311 56.724 177.343 56.788 ;
			RECT	177.479 56.724 177.511 56.788 ;
			RECT	177.647 56.724 177.679 56.788 ;
			RECT	177.815 56.724 177.847 56.788 ;
			RECT	177.983 56.724 178.015 56.788 ;
			RECT	178.151 56.724 178.183 56.788 ;
			RECT	178.319 56.724 178.351 56.788 ;
			RECT	178.487 56.724 178.519 56.788 ;
			RECT	178.655 56.724 178.687 56.788 ;
			RECT	178.823 56.724 178.855 56.788 ;
			RECT	178.991 56.724 179.023 56.788 ;
			RECT	179.159 56.724 179.191 56.788 ;
			RECT	179.327 56.724 179.359 56.788 ;
			RECT	179.495 56.724 179.527 56.788 ;
			RECT	179.663 56.724 179.695 56.788 ;
			RECT	179.831 56.724 179.863 56.788 ;
			RECT	179.999 56.724 180.031 56.788 ;
			RECT	180.167 56.724 180.199 56.788 ;
			RECT	180.335 56.724 180.367 56.788 ;
			RECT	180.503 56.724 180.535 56.788 ;
			RECT	180.671 56.724 180.703 56.788 ;
			RECT	180.839 56.724 180.871 56.788 ;
			RECT	181.007 56.724 181.039 56.788 ;
			RECT	181.175 56.724 181.207 56.788 ;
			RECT	181.343 56.724 181.375 56.788 ;
			RECT	181.511 56.724 181.543 56.788 ;
			RECT	181.679 56.724 181.711 56.788 ;
			RECT	181.847 56.724 181.879 56.788 ;
			RECT	182.015 56.724 182.047 56.788 ;
			RECT	182.183 56.724 182.215 56.788 ;
			RECT	182.351 56.724 182.383 56.788 ;
			RECT	182.519 56.724 182.551 56.788 ;
			RECT	182.687 56.724 182.719 56.788 ;
			RECT	182.855 56.724 182.887 56.788 ;
			RECT	183.023 56.724 183.055 56.788 ;
			RECT	183.191 56.724 183.223 56.788 ;
			RECT	183.359 56.724 183.391 56.788 ;
			RECT	183.527 56.724 183.559 56.788 ;
			RECT	183.695 56.724 183.727 56.788 ;
			RECT	183.863 56.724 183.895 56.788 ;
			RECT	184.031 56.724 184.063 56.788 ;
			RECT	184.199 56.724 184.231 56.788 ;
			RECT	184.367 56.724 184.399 56.788 ;
			RECT	184.535 56.724 184.567 56.788 ;
			RECT	184.703 56.724 184.735 56.788 ;
			RECT	184.871 56.724 184.903 56.788 ;
			RECT	185.039 56.724 185.071 56.788 ;
			RECT	185.207 56.724 185.239 56.788 ;
			RECT	185.375 56.724 185.407 56.788 ;
			RECT	185.543 56.724 185.575 56.788 ;
			RECT	185.711 56.724 185.743 56.788 ;
			RECT	185.879 56.724 185.911 56.788 ;
			RECT	186.047 56.724 186.079 56.788 ;
			RECT	186.215 56.724 186.247 56.788 ;
			RECT	186.383 56.724 186.415 56.788 ;
			RECT	186.551 56.724 186.583 56.788 ;
			RECT	186.719 56.724 186.751 56.788 ;
			RECT	186.887 56.724 186.919 56.788 ;
			RECT	187.055 56.724 187.087 56.788 ;
			RECT	187.223 56.724 187.255 56.788 ;
			RECT	187.391 56.724 187.423 56.788 ;
			RECT	187.559 56.724 187.591 56.788 ;
			RECT	187.727 56.724 187.759 56.788 ;
			RECT	187.895 56.724 187.927 56.788 ;
			RECT	188.063 56.724 188.095 56.788 ;
			RECT	188.231 56.724 188.263 56.788 ;
			RECT	188.399 56.724 188.431 56.788 ;
			RECT	188.567 56.724 188.599 56.788 ;
			RECT	188.735 56.724 188.767 56.788 ;
			RECT	188.903 56.724 188.935 56.788 ;
			RECT	189.071 56.724 189.103 56.788 ;
			RECT	189.239 56.724 189.271 56.788 ;
			RECT	189.407 56.724 189.439 56.788 ;
			RECT	189.575 56.724 189.607 56.788 ;
			RECT	189.743 56.724 189.775 56.788 ;
			RECT	189.911 56.724 189.943 56.788 ;
			RECT	190.079 56.724 190.111 56.788 ;
			RECT	190.247 56.724 190.279 56.788 ;
			RECT	190.415 56.724 190.447 56.788 ;
			RECT	190.583 56.724 190.615 56.788 ;
			RECT	190.751 56.724 190.783 56.788 ;
			RECT	190.919 56.724 190.951 56.788 ;
			RECT	191.087 56.724 191.119 56.788 ;
			RECT	191.255 56.724 191.287 56.788 ;
			RECT	191.423 56.724 191.455 56.788 ;
			RECT	191.591 56.724 191.623 56.788 ;
			RECT	191.759 56.724 191.791 56.788 ;
			RECT	191.927 56.724 191.959 56.788 ;
			RECT	192.095 56.724 192.127 56.788 ;
			RECT	192.263 56.724 192.295 56.788 ;
			RECT	192.431 56.724 192.463 56.788 ;
			RECT	192.599 56.724 192.631 56.788 ;
			RECT	192.767 56.724 192.799 56.788 ;
			RECT	192.935 56.724 192.967 56.788 ;
			RECT	193.103 56.724 193.135 56.788 ;
			RECT	193.271 56.724 193.303 56.788 ;
			RECT	193.439 56.724 193.471 56.788 ;
			RECT	193.607 56.724 193.639 56.788 ;
			RECT	193.775 56.724 193.807 56.788 ;
			RECT	193.943 56.724 193.975 56.788 ;
			RECT	194.111 56.724 194.143 56.788 ;
			RECT	194.279 56.724 194.311 56.788 ;
			RECT	194.447 56.724 194.479 56.788 ;
			RECT	194.615 56.724 194.647 56.788 ;
			RECT	194.783 56.724 194.815 56.788 ;
			RECT	194.951 56.724 194.983 56.788 ;
			RECT	195.119 56.724 195.151 56.788 ;
			RECT	195.287 56.724 195.319 56.788 ;
			RECT	195.455 56.724 195.487 56.788 ;
			RECT	195.623 56.724 195.655 56.788 ;
			RECT	195.791 56.724 195.823 56.788 ;
			RECT	195.959 56.724 195.991 56.788 ;
			RECT	196.127 56.724 196.159 56.788 ;
			RECT	196.295 56.724 196.327 56.788 ;
			RECT	196.463 56.724 196.495 56.788 ;
			RECT	196.631 56.724 196.663 56.788 ;
			RECT	196.799 56.724 196.831 56.788 ;
			RECT	196.967 56.724 196.999 56.788 ;
			RECT	197.135 56.724 197.167 56.788 ;
			RECT	197.303 56.724 197.335 56.788 ;
			RECT	197.471 56.724 197.503 56.788 ;
			RECT	197.639 56.724 197.671 56.788 ;
			RECT	197.807 56.724 197.839 56.788 ;
			RECT	197.975 56.724 198.007 56.788 ;
			RECT	198.143 56.724 198.175 56.788 ;
			RECT	198.311 56.724 198.343 56.788 ;
			RECT	198.479 56.724 198.511 56.788 ;
			RECT	198.647 56.724 198.679 56.788 ;
			RECT	198.815 56.724 198.847 56.788 ;
			RECT	198.983 56.724 199.015 56.788 ;
			RECT	199.151 56.724 199.183 56.788 ;
			RECT	199.319 56.724 199.351 56.788 ;
			RECT	199.487 56.724 199.519 56.788 ;
			RECT	199.655 56.724 199.687 56.788 ;
			RECT	199.823 56.724 199.855 56.788 ;
			RECT	199.991 56.724 200.023 56.788 ;
			RECT	200.121 56.74 200.153 56.772 ;
			RECT	200.243 56.735 200.275 56.767 ;
			RECT	200.373 56.724 200.405 56.788 ;
			RECT	200.9 56.724 200.932 56.788 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 54.776 201.665 54.896 ;
			LAYER	J3 ;
			RECT	0.755 54.804 0.787 54.868 ;
			RECT	1.645 54.804 1.709 54.868 ;
			RECT	2.323 54.804 2.387 54.868 ;
			RECT	3.438 54.804 3.47 54.868 ;
			RECT	3.585 54.804 3.617 54.868 ;
			RECT	4.195 54.804 4.227 54.868 ;
			RECT	4.72 54.804 4.752 54.868 ;
			RECT	4.944 54.804 5.008 54.868 ;
			RECT	5.267 54.804 5.299 54.868 ;
			RECT	5.797 54.804 5.829 54.868 ;
			RECT	5.927 54.815 5.959 54.847 ;
			RECT	6.049 54.82 6.081 54.852 ;
			RECT	6.179 54.804 6.211 54.868 ;
			RECT	6.347 54.804 6.379 54.868 ;
			RECT	6.515 54.804 6.547 54.868 ;
			RECT	6.683 54.804 6.715 54.868 ;
			RECT	6.851 54.804 6.883 54.868 ;
			RECT	7.019 54.804 7.051 54.868 ;
			RECT	7.187 54.804 7.219 54.868 ;
			RECT	7.355 54.804 7.387 54.868 ;
			RECT	7.523 54.804 7.555 54.868 ;
			RECT	7.691 54.804 7.723 54.868 ;
			RECT	7.859 54.804 7.891 54.868 ;
			RECT	8.027 54.804 8.059 54.868 ;
			RECT	8.195 54.804 8.227 54.868 ;
			RECT	8.363 54.804 8.395 54.868 ;
			RECT	8.531 54.804 8.563 54.868 ;
			RECT	8.699 54.804 8.731 54.868 ;
			RECT	8.867 54.804 8.899 54.868 ;
			RECT	9.035 54.804 9.067 54.868 ;
			RECT	9.203 54.804 9.235 54.868 ;
			RECT	9.371 54.804 9.403 54.868 ;
			RECT	9.539 54.804 9.571 54.868 ;
			RECT	9.707 54.804 9.739 54.868 ;
			RECT	9.875 54.804 9.907 54.868 ;
			RECT	10.043 54.804 10.075 54.868 ;
			RECT	10.211 54.804 10.243 54.868 ;
			RECT	10.379 54.804 10.411 54.868 ;
			RECT	10.547 54.804 10.579 54.868 ;
			RECT	10.715 54.804 10.747 54.868 ;
			RECT	10.883 54.804 10.915 54.868 ;
			RECT	11.051 54.804 11.083 54.868 ;
			RECT	11.219 54.804 11.251 54.868 ;
			RECT	11.387 54.804 11.419 54.868 ;
			RECT	11.555 54.804 11.587 54.868 ;
			RECT	11.723 54.804 11.755 54.868 ;
			RECT	11.891 54.804 11.923 54.868 ;
			RECT	12.059 54.804 12.091 54.868 ;
			RECT	12.227 54.804 12.259 54.868 ;
			RECT	12.395 54.804 12.427 54.868 ;
			RECT	12.563 54.804 12.595 54.868 ;
			RECT	12.731 54.804 12.763 54.868 ;
			RECT	12.899 54.804 12.931 54.868 ;
			RECT	13.067 54.804 13.099 54.868 ;
			RECT	13.235 54.804 13.267 54.868 ;
			RECT	13.403 54.804 13.435 54.868 ;
			RECT	13.571 54.804 13.603 54.868 ;
			RECT	13.739 54.804 13.771 54.868 ;
			RECT	13.907 54.804 13.939 54.868 ;
			RECT	14.075 54.804 14.107 54.868 ;
			RECT	14.243 54.804 14.275 54.868 ;
			RECT	14.411 54.804 14.443 54.868 ;
			RECT	14.579 54.804 14.611 54.868 ;
			RECT	14.747 54.804 14.779 54.868 ;
			RECT	14.915 54.804 14.947 54.868 ;
			RECT	15.083 54.804 15.115 54.868 ;
			RECT	15.251 54.804 15.283 54.868 ;
			RECT	15.419 54.804 15.451 54.868 ;
			RECT	15.587 54.804 15.619 54.868 ;
			RECT	15.755 54.804 15.787 54.868 ;
			RECT	15.923 54.804 15.955 54.868 ;
			RECT	16.091 54.804 16.123 54.868 ;
			RECT	16.259 54.804 16.291 54.868 ;
			RECT	16.427 54.804 16.459 54.868 ;
			RECT	16.595 54.804 16.627 54.868 ;
			RECT	16.763 54.804 16.795 54.868 ;
			RECT	16.931 54.804 16.963 54.868 ;
			RECT	17.099 54.804 17.131 54.868 ;
			RECT	17.267 54.804 17.299 54.868 ;
			RECT	17.435 54.804 17.467 54.868 ;
			RECT	17.603 54.804 17.635 54.868 ;
			RECT	17.771 54.804 17.803 54.868 ;
			RECT	17.939 54.804 17.971 54.868 ;
			RECT	18.107 54.804 18.139 54.868 ;
			RECT	18.275 54.804 18.307 54.868 ;
			RECT	18.443 54.804 18.475 54.868 ;
			RECT	18.611 54.804 18.643 54.868 ;
			RECT	18.779 54.804 18.811 54.868 ;
			RECT	18.947 54.804 18.979 54.868 ;
			RECT	19.115 54.804 19.147 54.868 ;
			RECT	19.283 54.804 19.315 54.868 ;
			RECT	19.451 54.804 19.483 54.868 ;
			RECT	19.619 54.804 19.651 54.868 ;
			RECT	19.787 54.804 19.819 54.868 ;
			RECT	19.955 54.804 19.987 54.868 ;
			RECT	20.123 54.804 20.155 54.868 ;
			RECT	20.291 54.804 20.323 54.868 ;
			RECT	20.459 54.804 20.491 54.868 ;
			RECT	20.627 54.804 20.659 54.868 ;
			RECT	20.795 54.804 20.827 54.868 ;
			RECT	20.963 54.804 20.995 54.868 ;
			RECT	21.131 54.804 21.163 54.868 ;
			RECT	21.299 54.804 21.331 54.868 ;
			RECT	21.467 54.804 21.499 54.868 ;
			RECT	21.635 54.804 21.667 54.868 ;
			RECT	21.803 54.804 21.835 54.868 ;
			RECT	21.971 54.804 22.003 54.868 ;
			RECT	22.139 54.804 22.171 54.868 ;
			RECT	22.307 54.804 22.339 54.868 ;
			RECT	22.475 54.804 22.507 54.868 ;
			RECT	22.643 54.804 22.675 54.868 ;
			RECT	22.811 54.804 22.843 54.868 ;
			RECT	22.979 54.804 23.011 54.868 ;
			RECT	23.147 54.804 23.179 54.868 ;
			RECT	23.315 54.804 23.347 54.868 ;
			RECT	23.483 54.804 23.515 54.868 ;
			RECT	23.651 54.804 23.683 54.868 ;
			RECT	23.819 54.804 23.851 54.868 ;
			RECT	23.987 54.804 24.019 54.868 ;
			RECT	24.155 54.804 24.187 54.868 ;
			RECT	24.323 54.804 24.355 54.868 ;
			RECT	24.491 54.804 24.523 54.868 ;
			RECT	24.659 54.804 24.691 54.868 ;
			RECT	24.827 54.804 24.859 54.868 ;
			RECT	24.995 54.804 25.027 54.868 ;
			RECT	25.163 54.804 25.195 54.868 ;
			RECT	25.331 54.804 25.363 54.868 ;
			RECT	25.499 54.804 25.531 54.868 ;
			RECT	25.667 54.804 25.699 54.868 ;
			RECT	25.835 54.804 25.867 54.868 ;
			RECT	26.003 54.804 26.035 54.868 ;
			RECT	26.171 54.804 26.203 54.868 ;
			RECT	26.339 54.804 26.371 54.868 ;
			RECT	26.507 54.804 26.539 54.868 ;
			RECT	26.675 54.804 26.707 54.868 ;
			RECT	26.843 54.804 26.875 54.868 ;
			RECT	27.011 54.804 27.043 54.868 ;
			RECT	27.179 54.804 27.211 54.868 ;
			RECT	27.347 54.804 27.379 54.868 ;
			RECT	27.515 54.804 27.547 54.868 ;
			RECT	27.683 54.804 27.715 54.868 ;
			RECT	27.851 54.804 27.883 54.868 ;
			RECT	28.019 54.804 28.051 54.868 ;
			RECT	28.187 54.804 28.219 54.868 ;
			RECT	28.355 54.804 28.387 54.868 ;
			RECT	28.523 54.804 28.555 54.868 ;
			RECT	28.691 54.804 28.723 54.868 ;
			RECT	28.859 54.804 28.891 54.868 ;
			RECT	29.027 54.804 29.059 54.868 ;
			RECT	29.195 54.804 29.227 54.868 ;
			RECT	29.363 54.804 29.395 54.868 ;
			RECT	29.531 54.804 29.563 54.868 ;
			RECT	29.699 54.804 29.731 54.868 ;
			RECT	29.867 54.804 29.899 54.868 ;
			RECT	30.035 54.804 30.067 54.868 ;
			RECT	30.203 54.804 30.235 54.868 ;
			RECT	30.371 54.804 30.403 54.868 ;
			RECT	30.539 54.804 30.571 54.868 ;
			RECT	30.707 54.804 30.739 54.868 ;
			RECT	30.875 54.804 30.907 54.868 ;
			RECT	31.043 54.804 31.075 54.868 ;
			RECT	31.211 54.804 31.243 54.868 ;
			RECT	31.379 54.804 31.411 54.868 ;
			RECT	31.547 54.804 31.579 54.868 ;
			RECT	31.715 54.804 31.747 54.868 ;
			RECT	31.883 54.804 31.915 54.868 ;
			RECT	32.051 54.804 32.083 54.868 ;
			RECT	32.219 54.804 32.251 54.868 ;
			RECT	32.387 54.804 32.419 54.868 ;
			RECT	32.555 54.804 32.587 54.868 ;
			RECT	32.723 54.804 32.755 54.868 ;
			RECT	32.891 54.804 32.923 54.868 ;
			RECT	33.059 54.804 33.091 54.868 ;
			RECT	33.227 54.804 33.259 54.868 ;
			RECT	33.395 54.804 33.427 54.868 ;
			RECT	33.563 54.804 33.595 54.868 ;
			RECT	33.731 54.804 33.763 54.868 ;
			RECT	33.899 54.804 33.931 54.868 ;
			RECT	34.067 54.804 34.099 54.868 ;
			RECT	34.235 54.804 34.267 54.868 ;
			RECT	34.403 54.804 34.435 54.868 ;
			RECT	34.571 54.804 34.603 54.868 ;
			RECT	34.739 54.804 34.771 54.868 ;
			RECT	34.907 54.804 34.939 54.868 ;
			RECT	35.075 54.804 35.107 54.868 ;
			RECT	35.243 54.804 35.275 54.868 ;
			RECT	35.411 54.804 35.443 54.868 ;
			RECT	35.579 54.804 35.611 54.868 ;
			RECT	35.747 54.804 35.779 54.868 ;
			RECT	35.915 54.804 35.947 54.868 ;
			RECT	36.083 54.804 36.115 54.868 ;
			RECT	36.251 54.804 36.283 54.868 ;
			RECT	36.419 54.804 36.451 54.868 ;
			RECT	36.587 54.804 36.619 54.868 ;
			RECT	36.755 54.804 36.787 54.868 ;
			RECT	36.923 54.804 36.955 54.868 ;
			RECT	37.091 54.804 37.123 54.868 ;
			RECT	37.259 54.804 37.291 54.868 ;
			RECT	37.427 54.804 37.459 54.868 ;
			RECT	37.595 54.804 37.627 54.868 ;
			RECT	37.763 54.804 37.795 54.868 ;
			RECT	37.931 54.804 37.963 54.868 ;
			RECT	38.099 54.804 38.131 54.868 ;
			RECT	38.267 54.804 38.299 54.868 ;
			RECT	38.435 54.804 38.467 54.868 ;
			RECT	38.603 54.804 38.635 54.868 ;
			RECT	38.771 54.804 38.803 54.868 ;
			RECT	38.939 54.804 38.971 54.868 ;
			RECT	39.107 54.804 39.139 54.868 ;
			RECT	39.275 54.804 39.307 54.868 ;
			RECT	39.443 54.804 39.475 54.868 ;
			RECT	39.611 54.804 39.643 54.868 ;
			RECT	39.779 54.804 39.811 54.868 ;
			RECT	39.947 54.804 39.979 54.868 ;
			RECT	40.115 54.804 40.147 54.868 ;
			RECT	40.283 54.804 40.315 54.868 ;
			RECT	40.451 54.804 40.483 54.868 ;
			RECT	40.619 54.804 40.651 54.868 ;
			RECT	40.787 54.804 40.819 54.868 ;
			RECT	40.955 54.804 40.987 54.868 ;
			RECT	41.123 54.804 41.155 54.868 ;
			RECT	41.291 54.804 41.323 54.868 ;
			RECT	41.459 54.804 41.491 54.868 ;
			RECT	41.627 54.804 41.659 54.868 ;
			RECT	41.795 54.804 41.827 54.868 ;
			RECT	41.963 54.804 41.995 54.868 ;
			RECT	42.131 54.804 42.163 54.868 ;
			RECT	42.299 54.804 42.331 54.868 ;
			RECT	42.467 54.804 42.499 54.868 ;
			RECT	42.635 54.804 42.667 54.868 ;
			RECT	42.803 54.804 42.835 54.868 ;
			RECT	42.971 54.804 43.003 54.868 ;
			RECT	43.139 54.804 43.171 54.868 ;
			RECT	43.307 54.804 43.339 54.868 ;
			RECT	43.475 54.804 43.507 54.868 ;
			RECT	43.643 54.804 43.675 54.868 ;
			RECT	43.811 54.804 43.843 54.868 ;
			RECT	43.979 54.804 44.011 54.868 ;
			RECT	44.147 54.804 44.179 54.868 ;
			RECT	44.315 54.804 44.347 54.868 ;
			RECT	44.483 54.804 44.515 54.868 ;
			RECT	44.651 54.804 44.683 54.868 ;
			RECT	44.819 54.804 44.851 54.868 ;
			RECT	44.987 54.804 45.019 54.868 ;
			RECT	45.155 54.804 45.187 54.868 ;
			RECT	45.323 54.804 45.355 54.868 ;
			RECT	45.491 54.804 45.523 54.868 ;
			RECT	45.659 54.804 45.691 54.868 ;
			RECT	45.827 54.804 45.859 54.868 ;
			RECT	45.995 54.804 46.027 54.868 ;
			RECT	46.163 54.804 46.195 54.868 ;
			RECT	46.331 54.804 46.363 54.868 ;
			RECT	46.499 54.804 46.531 54.868 ;
			RECT	46.667 54.804 46.699 54.868 ;
			RECT	46.835 54.804 46.867 54.868 ;
			RECT	47.003 54.804 47.035 54.868 ;
			RECT	47.171 54.804 47.203 54.868 ;
			RECT	47.339 54.804 47.371 54.868 ;
			RECT	47.507 54.804 47.539 54.868 ;
			RECT	47.675 54.804 47.707 54.868 ;
			RECT	47.843 54.804 47.875 54.868 ;
			RECT	48.011 54.804 48.043 54.868 ;
			RECT	48.179 54.804 48.211 54.868 ;
			RECT	48.347 54.804 48.379 54.868 ;
			RECT	48.515 54.804 48.547 54.868 ;
			RECT	48.683 54.804 48.715 54.868 ;
			RECT	48.851 54.804 48.883 54.868 ;
			RECT	49.019 54.804 49.051 54.868 ;
			RECT	49.187 54.804 49.219 54.868 ;
			RECT	49.318 54.82 49.35 54.852 ;
			RECT	49.439 54.82 49.471 54.852 ;
			RECT	49.569 54.804 49.601 54.868 ;
			RECT	51.881 54.804 51.913 54.868 ;
			RECT	53.132 54.804 53.196 54.868 ;
			RECT	53.812 54.804 53.844 54.868 ;
			RECT	54.251 54.804 54.283 54.868 ;
			RECT	55.562 54.804 55.626 54.868 ;
			RECT	58.603 54.804 58.635 54.868 ;
			RECT	58.733 54.82 58.765 54.852 ;
			RECT	58.854 54.82 58.886 54.852 ;
			RECT	58.985 54.804 59.017 54.868 ;
			RECT	59.153 54.804 59.185 54.868 ;
			RECT	59.321 54.804 59.353 54.868 ;
			RECT	59.489 54.804 59.521 54.868 ;
			RECT	59.657 54.804 59.689 54.868 ;
			RECT	59.825 54.804 59.857 54.868 ;
			RECT	59.993 54.804 60.025 54.868 ;
			RECT	60.161 54.804 60.193 54.868 ;
			RECT	60.329 54.804 60.361 54.868 ;
			RECT	60.497 54.804 60.529 54.868 ;
			RECT	60.665 54.804 60.697 54.868 ;
			RECT	60.833 54.804 60.865 54.868 ;
			RECT	61.001 54.804 61.033 54.868 ;
			RECT	61.169 54.804 61.201 54.868 ;
			RECT	61.337 54.804 61.369 54.868 ;
			RECT	61.505 54.804 61.537 54.868 ;
			RECT	61.673 54.804 61.705 54.868 ;
			RECT	61.841 54.804 61.873 54.868 ;
			RECT	62.009 54.804 62.041 54.868 ;
			RECT	62.177 54.804 62.209 54.868 ;
			RECT	62.345 54.804 62.377 54.868 ;
			RECT	62.513 54.804 62.545 54.868 ;
			RECT	62.681 54.804 62.713 54.868 ;
			RECT	62.849 54.804 62.881 54.868 ;
			RECT	63.017 54.804 63.049 54.868 ;
			RECT	63.185 54.804 63.217 54.868 ;
			RECT	63.353 54.804 63.385 54.868 ;
			RECT	63.521 54.804 63.553 54.868 ;
			RECT	63.689 54.804 63.721 54.868 ;
			RECT	63.857 54.804 63.889 54.868 ;
			RECT	64.025 54.804 64.057 54.868 ;
			RECT	64.193 54.804 64.225 54.868 ;
			RECT	64.361 54.804 64.393 54.868 ;
			RECT	64.529 54.804 64.561 54.868 ;
			RECT	64.697 54.804 64.729 54.868 ;
			RECT	64.865 54.804 64.897 54.868 ;
			RECT	65.033 54.804 65.065 54.868 ;
			RECT	65.201 54.804 65.233 54.868 ;
			RECT	65.369 54.804 65.401 54.868 ;
			RECT	65.537 54.804 65.569 54.868 ;
			RECT	65.705 54.804 65.737 54.868 ;
			RECT	65.873 54.804 65.905 54.868 ;
			RECT	66.041 54.804 66.073 54.868 ;
			RECT	66.209 54.804 66.241 54.868 ;
			RECT	66.377 54.804 66.409 54.868 ;
			RECT	66.545 54.804 66.577 54.868 ;
			RECT	66.713 54.804 66.745 54.868 ;
			RECT	66.881 54.804 66.913 54.868 ;
			RECT	67.049 54.804 67.081 54.868 ;
			RECT	67.217 54.804 67.249 54.868 ;
			RECT	67.385 54.804 67.417 54.868 ;
			RECT	67.553 54.804 67.585 54.868 ;
			RECT	67.721 54.804 67.753 54.868 ;
			RECT	67.889 54.804 67.921 54.868 ;
			RECT	68.057 54.804 68.089 54.868 ;
			RECT	68.225 54.804 68.257 54.868 ;
			RECT	68.393 54.804 68.425 54.868 ;
			RECT	68.561 54.804 68.593 54.868 ;
			RECT	68.729 54.804 68.761 54.868 ;
			RECT	68.897 54.804 68.929 54.868 ;
			RECT	69.065 54.804 69.097 54.868 ;
			RECT	69.233 54.804 69.265 54.868 ;
			RECT	69.401 54.804 69.433 54.868 ;
			RECT	69.569 54.804 69.601 54.868 ;
			RECT	69.737 54.804 69.769 54.868 ;
			RECT	69.905 54.804 69.937 54.868 ;
			RECT	70.073 54.804 70.105 54.868 ;
			RECT	70.241 54.804 70.273 54.868 ;
			RECT	70.409 54.804 70.441 54.868 ;
			RECT	70.577 54.804 70.609 54.868 ;
			RECT	70.745 54.804 70.777 54.868 ;
			RECT	70.913 54.804 70.945 54.868 ;
			RECT	71.081 54.804 71.113 54.868 ;
			RECT	71.249 54.804 71.281 54.868 ;
			RECT	71.417 54.804 71.449 54.868 ;
			RECT	71.585 54.804 71.617 54.868 ;
			RECT	71.753 54.804 71.785 54.868 ;
			RECT	71.921 54.804 71.953 54.868 ;
			RECT	72.089 54.804 72.121 54.868 ;
			RECT	72.257 54.804 72.289 54.868 ;
			RECT	72.425 54.804 72.457 54.868 ;
			RECT	72.593 54.804 72.625 54.868 ;
			RECT	72.761 54.804 72.793 54.868 ;
			RECT	72.929 54.804 72.961 54.868 ;
			RECT	73.097 54.804 73.129 54.868 ;
			RECT	73.265 54.804 73.297 54.868 ;
			RECT	73.433 54.804 73.465 54.868 ;
			RECT	73.601 54.804 73.633 54.868 ;
			RECT	73.769 54.804 73.801 54.868 ;
			RECT	73.937 54.804 73.969 54.868 ;
			RECT	74.105 54.804 74.137 54.868 ;
			RECT	74.273 54.804 74.305 54.868 ;
			RECT	74.441 54.804 74.473 54.868 ;
			RECT	74.609 54.804 74.641 54.868 ;
			RECT	74.777 54.804 74.809 54.868 ;
			RECT	74.945 54.804 74.977 54.868 ;
			RECT	75.113 54.804 75.145 54.868 ;
			RECT	75.281 54.804 75.313 54.868 ;
			RECT	75.449 54.804 75.481 54.868 ;
			RECT	75.617 54.804 75.649 54.868 ;
			RECT	75.785 54.804 75.817 54.868 ;
			RECT	75.953 54.804 75.985 54.868 ;
			RECT	76.121 54.804 76.153 54.868 ;
			RECT	76.289 54.804 76.321 54.868 ;
			RECT	76.457 54.804 76.489 54.868 ;
			RECT	76.625 54.804 76.657 54.868 ;
			RECT	76.793 54.804 76.825 54.868 ;
			RECT	76.961 54.804 76.993 54.868 ;
			RECT	77.129 54.804 77.161 54.868 ;
			RECT	77.297 54.804 77.329 54.868 ;
			RECT	77.465 54.804 77.497 54.868 ;
			RECT	77.633 54.804 77.665 54.868 ;
			RECT	77.801 54.804 77.833 54.868 ;
			RECT	77.969 54.804 78.001 54.868 ;
			RECT	78.137 54.804 78.169 54.868 ;
			RECT	78.305 54.804 78.337 54.868 ;
			RECT	78.473 54.804 78.505 54.868 ;
			RECT	78.641 54.804 78.673 54.868 ;
			RECT	78.809 54.804 78.841 54.868 ;
			RECT	78.977 54.804 79.009 54.868 ;
			RECT	79.145 54.804 79.177 54.868 ;
			RECT	79.313 54.804 79.345 54.868 ;
			RECT	79.481 54.804 79.513 54.868 ;
			RECT	79.649 54.804 79.681 54.868 ;
			RECT	79.817 54.804 79.849 54.868 ;
			RECT	79.985 54.804 80.017 54.868 ;
			RECT	80.153 54.804 80.185 54.868 ;
			RECT	80.321 54.804 80.353 54.868 ;
			RECT	80.489 54.804 80.521 54.868 ;
			RECT	80.657 54.804 80.689 54.868 ;
			RECT	80.825 54.804 80.857 54.868 ;
			RECT	80.993 54.804 81.025 54.868 ;
			RECT	81.161 54.804 81.193 54.868 ;
			RECT	81.329 54.804 81.361 54.868 ;
			RECT	81.497 54.804 81.529 54.868 ;
			RECT	81.665 54.804 81.697 54.868 ;
			RECT	81.833 54.804 81.865 54.868 ;
			RECT	82.001 54.804 82.033 54.868 ;
			RECT	82.169 54.804 82.201 54.868 ;
			RECT	82.337 54.804 82.369 54.868 ;
			RECT	82.505 54.804 82.537 54.868 ;
			RECT	82.673 54.804 82.705 54.868 ;
			RECT	82.841 54.804 82.873 54.868 ;
			RECT	83.009 54.804 83.041 54.868 ;
			RECT	83.177 54.804 83.209 54.868 ;
			RECT	83.345 54.804 83.377 54.868 ;
			RECT	83.513 54.804 83.545 54.868 ;
			RECT	83.681 54.804 83.713 54.868 ;
			RECT	83.849 54.804 83.881 54.868 ;
			RECT	84.017 54.804 84.049 54.868 ;
			RECT	84.185 54.804 84.217 54.868 ;
			RECT	84.353 54.804 84.385 54.868 ;
			RECT	84.521 54.804 84.553 54.868 ;
			RECT	84.689 54.804 84.721 54.868 ;
			RECT	84.857 54.804 84.889 54.868 ;
			RECT	85.025 54.804 85.057 54.868 ;
			RECT	85.193 54.804 85.225 54.868 ;
			RECT	85.361 54.804 85.393 54.868 ;
			RECT	85.529 54.804 85.561 54.868 ;
			RECT	85.697 54.804 85.729 54.868 ;
			RECT	85.865 54.804 85.897 54.868 ;
			RECT	86.033 54.804 86.065 54.868 ;
			RECT	86.201 54.804 86.233 54.868 ;
			RECT	86.369 54.804 86.401 54.868 ;
			RECT	86.537 54.804 86.569 54.868 ;
			RECT	86.705 54.804 86.737 54.868 ;
			RECT	86.873 54.804 86.905 54.868 ;
			RECT	87.041 54.804 87.073 54.868 ;
			RECT	87.209 54.804 87.241 54.868 ;
			RECT	87.377 54.804 87.409 54.868 ;
			RECT	87.545 54.804 87.577 54.868 ;
			RECT	87.713 54.804 87.745 54.868 ;
			RECT	87.881 54.804 87.913 54.868 ;
			RECT	88.049 54.804 88.081 54.868 ;
			RECT	88.217 54.804 88.249 54.868 ;
			RECT	88.385 54.804 88.417 54.868 ;
			RECT	88.553 54.804 88.585 54.868 ;
			RECT	88.721 54.804 88.753 54.868 ;
			RECT	88.889 54.804 88.921 54.868 ;
			RECT	89.057 54.804 89.089 54.868 ;
			RECT	89.225 54.804 89.257 54.868 ;
			RECT	89.393 54.804 89.425 54.868 ;
			RECT	89.561 54.804 89.593 54.868 ;
			RECT	89.729 54.804 89.761 54.868 ;
			RECT	89.897 54.804 89.929 54.868 ;
			RECT	90.065 54.804 90.097 54.868 ;
			RECT	90.233 54.804 90.265 54.868 ;
			RECT	90.401 54.804 90.433 54.868 ;
			RECT	90.569 54.804 90.601 54.868 ;
			RECT	90.737 54.804 90.769 54.868 ;
			RECT	90.905 54.804 90.937 54.868 ;
			RECT	91.073 54.804 91.105 54.868 ;
			RECT	91.241 54.804 91.273 54.868 ;
			RECT	91.409 54.804 91.441 54.868 ;
			RECT	91.577 54.804 91.609 54.868 ;
			RECT	91.745 54.804 91.777 54.868 ;
			RECT	91.913 54.804 91.945 54.868 ;
			RECT	92.081 54.804 92.113 54.868 ;
			RECT	92.249 54.804 92.281 54.868 ;
			RECT	92.417 54.804 92.449 54.868 ;
			RECT	92.585 54.804 92.617 54.868 ;
			RECT	92.753 54.804 92.785 54.868 ;
			RECT	92.921 54.804 92.953 54.868 ;
			RECT	93.089 54.804 93.121 54.868 ;
			RECT	93.257 54.804 93.289 54.868 ;
			RECT	93.425 54.804 93.457 54.868 ;
			RECT	93.593 54.804 93.625 54.868 ;
			RECT	93.761 54.804 93.793 54.868 ;
			RECT	93.929 54.804 93.961 54.868 ;
			RECT	94.097 54.804 94.129 54.868 ;
			RECT	94.265 54.804 94.297 54.868 ;
			RECT	94.433 54.804 94.465 54.868 ;
			RECT	94.601 54.804 94.633 54.868 ;
			RECT	94.769 54.804 94.801 54.868 ;
			RECT	94.937 54.804 94.969 54.868 ;
			RECT	95.105 54.804 95.137 54.868 ;
			RECT	95.273 54.804 95.305 54.868 ;
			RECT	95.441 54.804 95.473 54.868 ;
			RECT	95.609 54.804 95.641 54.868 ;
			RECT	95.777 54.804 95.809 54.868 ;
			RECT	95.945 54.804 95.977 54.868 ;
			RECT	96.113 54.804 96.145 54.868 ;
			RECT	96.281 54.804 96.313 54.868 ;
			RECT	96.449 54.804 96.481 54.868 ;
			RECT	96.617 54.804 96.649 54.868 ;
			RECT	96.785 54.804 96.817 54.868 ;
			RECT	96.953 54.804 96.985 54.868 ;
			RECT	97.121 54.804 97.153 54.868 ;
			RECT	97.289 54.804 97.321 54.868 ;
			RECT	97.457 54.804 97.489 54.868 ;
			RECT	97.625 54.804 97.657 54.868 ;
			RECT	97.793 54.804 97.825 54.868 ;
			RECT	97.961 54.804 97.993 54.868 ;
			RECT	98.129 54.804 98.161 54.868 ;
			RECT	98.297 54.804 98.329 54.868 ;
			RECT	98.465 54.804 98.497 54.868 ;
			RECT	98.633 54.804 98.665 54.868 ;
			RECT	98.801 54.804 98.833 54.868 ;
			RECT	98.969 54.804 99.001 54.868 ;
			RECT	99.137 54.804 99.169 54.868 ;
			RECT	99.305 54.804 99.337 54.868 ;
			RECT	99.473 54.804 99.505 54.868 ;
			RECT	99.641 54.804 99.673 54.868 ;
			RECT	99.809 54.804 99.841 54.868 ;
			RECT	99.977 54.804 100.009 54.868 ;
			RECT	100.145 54.804 100.177 54.868 ;
			RECT	100.313 54.804 100.345 54.868 ;
			RECT	100.481 54.804 100.513 54.868 ;
			RECT	100.649 54.804 100.681 54.868 ;
			RECT	100.817 54.804 100.849 54.868 ;
			RECT	100.985 54.804 101.017 54.868 ;
			RECT	101.153 54.804 101.185 54.868 ;
			RECT	101.321 54.804 101.353 54.868 ;
			RECT	101.489 54.804 101.521 54.868 ;
			RECT	101.657 54.804 101.689 54.868 ;
			RECT	101.825 54.804 101.857 54.868 ;
			RECT	101.993 54.804 102.025 54.868 ;
			RECT	102.123 54.82 102.155 54.852 ;
			RECT	102.245 54.815 102.277 54.847 ;
			RECT	102.375 54.804 102.407 54.868 ;
			RECT	103.795 54.804 103.827 54.868 ;
			RECT	103.925 54.815 103.957 54.847 ;
			RECT	104.047 54.82 104.079 54.852 ;
			RECT	104.177 54.804 104.209 54.868 ;
			RECT	104.345 54.804 104.377 54.868 ;
			RECT	104.513 54.804 104.545 54.868 ;
			RECT	104.681 54.804 104.713 54.868 ;
			RECT	104.849 54.804 104.881 54.868 ;
			RECT	105.017 54.804 105.049 54.868 ;
			RECT	105.185 54.804 105.217 54.868 ;
			RECT	105.353 54.804 105.385 54.868 ;
			RECT	105.521 54.804 105.553 54.868 ;
			RECT	105.689 54.804 105.721 54.868 ;
			RECT	105.857 54.804 105.889 54.868 ;
			RECT	106.025 54.804 106.057 54.868 ;
			RECT	106.193 54.804 106.225 54.868 ;
			RECT	106.361 54.804 106.393 54.868 ;
			RECT	106.529 54.804 106.561 54.868 ;
			RECT	106.697 54.804 106.729 54.868 ;
			RECT	106.865 54.804 106.897 54.868 ;
			RECT	107.033 54.804 107.065 54.868 ;
			RECT	107.201 54.804 107.233 54.868 ;
			RECT	107.369 54.804 107.401 54.868 ;
			RECT	107.537 54.804 107.569 54.868 ;
			RECT	107.705 54.804 107.737 54.868 ;
			RECT	107.873 54.804 107.905 54.868 ;
			RECT	108.041 54.804 108.073 54.868 ;
			RECT	108.209 54.804 108.241 54.868 ;
			RECT	108.377 54.804 108.409 54.868 ;
			RECT	108.545 54.804 108.577 54.868 ;
			RECT	108.713 54.804 108.745 54.868 ;
			RECT	108.881 54.804 108.913 54.868 ;
			RECT	109.049 54.804 109.081 54.868 ;
			RECT	109.217 54.804 109.249 54.868 ;
			RECT	109.385 54.804 109.417 54.868 ;
			RECT	109.553 54.804 109.585 54.868 ;
			RECT	109.721 54.804 109.753 54.868 ;
			RECT	109.889 54.804 109.921 54.868 ;
			RECT	110.057 54.804 110.089 54.868 ;
			RECT	110.225 54.804 110.257 54.868 ;
			RECT	110.393 54.804 110.425 54.868 ;
			RECT	110.561 54.804 110.593 54.868 ;
			RECT	110.729 54.804 110.761 54.868 ;
			RECT	110.897 54.804 110.929 54.868 ;
			RECT	111.065 54.804 111.097 54.868 ;
			RECT	111.233 54.804 111.265 54.868 ;
			RECT	111.401 54.804 111.433 54.868 ;
			RECT	111.569 54.804 111.601 54.868 ;
			RECT	111.737 54.804 111.769 54.868 ;
			RECT	111.905 54.804 111.937 54.868 ;
			RECT	112.073 54.804 112.105 54.868 ;
			RECT	112.241 54.804 112.273 54.868 ;
			RECT	112.409 54.804 112.441 54.868 ;
			RECT	112.577 54.804 112.609 54.868 ;
			RECT	112.745 54.804 112.777 54.868 ;
			RECT	112.913 54.804 112.945 54.868 ;
			RECT	113.081 54.804 113.113 54.868 ;
			RECT	113.249 54.804 113.281 54.868 ;
			RECT	113.417 54.804 113.449 54.868 ;
			RECT	113.585 54.804 113.617 54.868 ;
			RECT	113.753 54.804 113.785 54.868 ;
			RECT	113.921 54.804 113.953 54.868 ;
			RECT	114.089 54.804 114.121 54.868 ;
			RECT	114.257 54.804 114.289 54.868 ;
			RECT	114.425 54.804 114.457 54.868 ;
			RECT	114.593 54.804 114.625 54.868 ;
			RECT	114.761 54.804 114.793 54.868 ;
			RECT	114.929 54.804 114.961 54.868 ;
			RECT	115.097 54.804 115.129 54.868 ;
			RECT	115.265 54.804 115.297 54.868 ;
			RECT	115.433 54.804 115.465 54.868 ;
			RECT	115.601 54.804 115.633 54.868 ;
			RECT	115.769 54.804 115.801 54.868 ;
			RECT	115.937 54.804 115.969 54.868 ;
			RECT	116.105 54.804 116.137 54.868 ;
			RECT	116.273 54.804 116.305 54.868 ;
			RECT	116.441 54.804 116.473 54.868 ;
			RECT	116.609 54.804 116.641 54.868 ;
			RECT	116.777 54.804 116.809 54.868 ;
			RECT	116.945 54.804 116.977 54.868 ;
			RECT	117.113 54.804 117.145 54.868 ;
			RECT	117.281 54.804 117.313 54.868 ;
			RECT	117.449 54.804 117.481 54.868 ;
			RECT	117.617 54.804 117.649 54.868 ;
			RECT	117.785 54.804 117.817 54.868 ;
			RECT	117.953 54.804 117.985 54.868 ;
			RECT	118.121 54.804 118.153 54.868 ;
			RECT	118.289 54.804 118.321 54.868 ;
			RECT	118.457 54.804 118.489 54.868 ;
			RECT	118.625 54.804 118.657 54.868 ;
			RECT	118.793 54.804 118.825 54.868 ;
			RECT	118.961 54.804 118.993 54.868 ;
			RECT	119.129 54.804 119.161 54.868 ;
			RECT	119.297 54.804 119.329 54.868 ;
			RECT	119.465 54.804 119.497 54.868 ;
			RECT	119.633 54.804 119.665 54.868 ;
			RECT	119.801 54.804 119.833 54.868 ;
			RECT	119.969 54.804 120.001 54.868 ;
			RECT	120.137 54.804 120.169 54.868 ;
			RECT	120.305 54.804 120.337 54.868 ;
			RECT	120.473 54.804 120.505 54.868 ;
			RECT	120.641 54.804 120.673 54.868 ;
			RECT	120.809 54.804 120.841 54.868 ;
			RECT	120.977 54.804 121.009 54.868 ;
			RECT	121.145 54.804 121.177 54.868 ;
			RECT	121.313 54.804 121.345 54.868 ;
			RECT	121.481 54.804 121.513 54.868 ;
			RECT	121.649 54.804 121.681 54.868 ;
			RECT	121.817 54.804 121.849 54.868 ;
			RECT	121.985 54.804 122.017 54.868 ;
			RECT	122.153 54.804 122.185 54.868 ;
			RECT	122.321 54.804 122.353 54.868 ;
			RECT	122.489 54.804 122.521 54.868 ;
			RECT	122.657 54.804 122.689 54.868 ;
			RECT	122.825 54.804 122.857 54.868 ;
			RECT	122.993 54.804 123.025 54.868 ;
			RECT	123.161 54.804 123.193 54.868 ;
			RECT	123.329 54.804 123.361 54.868 ;
			RECT	123.497 54.804 123.529 54.868 ;
			RECT	123.665 54.804 123.697 54.868 ;
			RECT	123.833 54.804 123.865 54.868 ;
			RECT	124.001 54.804 124.033 54.868 ;
			RECT	124.169 54.804 124.201 54.868 ;
			RECT	124.337 54.804 124.369 54.868 ;
			RECT	124.505 54.804 124.537 54.868 ;
			RECT	124.673 54.804 124.705 54.868 ;
			RECT	124.841 54.804 124.873 54.868 ;
			RECT	125.009 54.804 125.041 54.868 ;
			RECT	125.177 54.804 125.209 54.868 ;
			RECT	125.345 54.804 125.377 54.868 ;
			RECT	125.513 54.804 125.545 54.868 ;
			RECT	125.681 54.804 125.713 54.868 ;
			RECT	125.849 54.804 125.881 54.868 ;
			RECT	126.017 54.804 126.049 54.868 ;
			RECT	126.185 54.804 126.217 54.868 ;
			RECT	126.353 54.804 126.385 54.868 ;
			RECT	126.521 54.804 126.553 54.868 ;
			RECT	126.689 54.804 126.721 54.868 ;
			RECT	126.857 54.804 126.889 54.868 ;
			RECT	127.025 54.804 127.057 54.868 ;
			RECT	127.193 54.804 127.225 54.868 ;
			RECT	127.361 54.804 127.393 54.868 ;
			RECT	127.529 54.804 127.561 54.868 ;
			RECT	127.697 54.804 127.729 54.868 ;
			RECT	127.865 54.804 127.897 54.868 ;
			RECT	128.033 54.804 128.065 54.868 ;
			RECT	128.201 54.804 128.233 54.868 ;
			RECT	128.369 54.804 128.401 54.868 ;
			RECT	128.537 54.804 128.569 54.868 ;
			RECT	128.705 54.804 128.737 54.868 ;
			RECT	128.873 54.804 128.905 54.868 ;
			RECT	129.041 54.804 129.073 54.868 ;
			RECT	129.209 54.804 129.241 54.868 ;
			RECT	129.377 54.804 129.409 54.868 ;
			RECT	129.545 54.804 129.577 54.868 ;
			RECT	129.713 54.804 129.745 54.868 ;
			RECT	129.881 54.804 129.913 54.868 ;
			RECT	130.049 54.804 130.081 54.868 ;
			RECT	130.217 54.804 130.249 54.868 ;
			RECT	130.385 54.804 130.417 54.868 ;
			RECT	130.553 54.804 130.585 54.868 ;
			RECT	130.721 54.804 130.753 54.868 ;
			RECT	130.889 54.804 130.921 54.868 ;
			RECT	131.057 54.804 131.089 54.868 ;
			RECT	131.225 54.804 131.257 54.868 ;
			RECT	131.393 54.804 131.425 54.868 ;
			RECT	131.561 54.804 131.593 54.868 ;
			RECT	131.729 54.804 131.761 54.868 ;
			RECT	131.897 54.804 131.929 54.868 ;
			RECT	132.065 54.804 132.097 54.868 ;
			RECT	132.233 54.804 132.265 54.868 ;
			RECT	132.401 54.804 132.433 54.868 ;
			RECT	132.569 54.804 132.601 54.868 ;
			RECT	132.737 54.804 132.769 54.868 ;
			RECT	132.905 54.804 132.937 54.868 ;
			RECT	133.073 54.804 133.105 54.868 ;
			RECT	133.241 54.804 133.273 54.868 ;
			RECT	133.409 54.804 133.441 54.868 ;
			RECT	133.577 54.804 133.609 54.868 ;
			RECT	133.745 54.804 133.777 54.868 ;
			RECT	133.913 54.804 133.945 54.868 ;
			RECT	134.081 54.804 134.113 54.868 ;
			RECT	134.249 54.804 134.281 54.868 ;
			RECT	134.417 54.804 134.449 54.868 ;
			RECT	134.585 54.804 134.617 54.868 ;
			RECT	134.753 54.804 134.785 54.868 ;
			RECT	134.921 54.804 134.953 54.868 ;
			RECT	135.089 54.804 135.121 54.868 ;
			RECT	135.257 54.804 135.289 54.868 ;
			RECT	135.425 54.804 135.457 54.868 ;
			RECT	135.593 54.804 135.625 54.868 ;
			RECT	135.761 54.804 135.793 54.868 ;
			RECT	135.929 54.804 135.961 54.868 ;
			RECT	136.097 54.804 136.129 54.868 ;
			RECT	136.265 54.804 136.297 54.868 ;
			RECT	136.433 54.804 136.465 54.868 ;
			RECT	136.601 54.804 136.633 54.868 ;
			RECT	136.769 54.804 136.801 54.868 ;
			RECT	136.937 54.804 136.969 54.868 ;
			RECT	137.105 54.804 137.137 54.868 ;
			RECT	137.273 54.804 137.305 54.868 ;
			RECT	137.441 54.804 137.473 54.868 ;
			RECT	137.609 54.804 137.641 54.868 ;
			RECT	137.777 54.804 137.809 54.868 ;
			RECT	137.945 54.804 137.977 54.868 ;
			RECT	138.113 54.804 138.145 54.868 ;
			RECT	138.281 54.804 138.313 54.868 ;
			RECT	138.449 54.804 138.481 54.868 ;
			RECT	138.617 54.804 138.649 54.868 ;
			RECT	138.785 54.804 138.817 54.868 ;
			RECT	138.953 54.804 138.985 54.868 ;
			RECT	139.121 54.804 139.153 54.868 ;
			RECT	139.289 54.804 139.321 54.868 ;
			RECT	139.457 54.804 139.489 54.868 ;
			RECT	139.625 54.804 139.657 54.868 ;
			RECT	139.793 54.804 139.825 54.868 ;
			RECT	139.961 54.804 139.993 54.868 ;
			RECT	140.129 54.804 140.161 54.868 ;
			RECT	140.297 54.804 140.329 54.868 ;
			RECT	140.465 54.804 140.497 54.868 ;
			RECT	140.633 54.804 140.665 54.868 ;
			RECT	140.801 54.804 140.833 54.868 ;
			RECT	140.969 54.804 141.001 54.868 ;
			RECT	141.137 54.804 141.169 54.868 ;
			RECT	141.305 54.804 141.337 54.868 ;
			RECT	141.473 54.804 141.505 54.868 ;
			RECT	141.641 54.804 141.673 54.868 ;
			RECT	141.809 54.804 141.841 54.868 ;
			RECT	141.977 54.804 142.009 54.868 ;
			RECT	142.145 54.804 142.177 54.868 ;
			RECT	142.313 54.804 142.345 54.868 ;
			RECT	142.481 54.804 142.513 54.868 ;
			RECT	142.649 54.804 142.681 54.868 ;
			RECT	142.817 54.804 142.849 54.868 ;
			RECT	142.985 54.804 143.017 54.868 ;
			RECT	143.153 54.804 143.185 54.868 ;
			RECT	143.321 54.804 143.353 54.868 ;
			RECT	143.489 54.804 143.521 54.868 ;
			RECT	143.657 54.804 143.689 54.868 ;
			RECT	143.825 54.804 143.857 54.868 ;
			RECT	143.993 54.804 144.025 54.868 ;
			RECT	144.161 54.804 144.193 54.868 ;
			RECT	144.329 54.804 144.361 54.868 ;
			RECT	144.497 54.804 144.529 54.868 ;
			RECT	144.665 54.804 144.697 54.868 ;
			RECT	144.833 54.804 144.865 54.868 ;
			RECT	145.001 54.804 145.033 54.868 ;
			RECT	145.169 54.804 145.201 54.868 ;
			RECT	145.337 54.804 145.369 54.868 ;
			RECT	145.505 54.804 145.537 54.868 ;
			RECT	145.673 54.804 145.705 54.868 ;
			RECT	145.841 54.804 145.873 54.868 ;
			RECT	146.009 54.804 146.041 54.868 ;
			RECT	146.177 54.804 146.209 54.868 ;
			RECT	146.345 54.804 146.377 54.868 ;
			RECT	146.513 54.804 146.545 54.868 ;
			RECT	146.681 54.804 146.713 54.868 ;
			RECT	146.849 54.804 146.881 54.868 ;
			RECT	147.017 54.804 147.049 54.868 ;
			RECT	147.185 54.804 147.217 54.868 ;
			RECT	147.316 54.82 147.348 54.852 ;
			RECT	147.437 54.82 147.469 54.852 ;
			RECT	147.567 54.804 147.599 54.868 ;
			RECT	149.879 54.804 149.911 54.868 ;
			RECT	151.13 54.804 151.194 54.868 ;
			RECT	151.81 54.804 151.842 54.868 ;
			RECT	152.249 54.804 152.281 54.868 ;
			RECT	153.56 54.804 153.624 54.868 ;
			RECT	156.601 54.804 156.633 54.868 ;
			RECT	156.731 54.82 156.763 54.852 ;
			RECT	156.852 54.82 156.884 54.852 ;
			RECT	156.983 54.804 157.015 54.868 ;
			RECT	157.151 54.804 157.183 54.868 ;
			RECT	157.319 54.804 157.351 54.868 ;
			RECT	157.487 54.804 157.519 54.868 ;
			RECT	157.655 54.804 157.687 54.868 ;
			RECT	157.823 54.804 157.855 54.868 ;
			RECT	157.991 54.804 158.023 54.868 ;
			RECT	158.159 54.804 158.191 54.868 ;
			RECT	158.327 54.804 158.359 54.868 ;
			RECT	158.495 54.804 158.527 54.868 ;
			RECT	158.663 54.804 158.695 54.868 ;
			RECT	158.831 54.804 158.863 54.868 ;
			RECT	158.999 54.804 159.031 54.868 ;
			RECT	159.167 54.804 159.199 54.868 ;
			RECT	159.335 54.804 159.367 54.868 ;
			RECT	159.503 54.804 159.535 54.868 ;
			RECT	159.671 54.804 159.703 54.868 ;
			RECT	159.839 54.804 159.871 54.868 ;
			RECT	160.007 54.804 160.039 54.868 ;
			RECT	160.175 54.804 160.207 54.868 ;
			RECT	160.343 54.804 160.375 54.868 ;
			RECT	160.511 54.804 160.543 54.868 ;
			RECT	160.679 54.804 160.711 54.868 ;
			RECT	160.847 54.804 160.879 54.868 ;
			RECT	161.015 54.804 161.047 54.868 ;
			RECT	161.183 54.804 161.215 54.868 ;
			RECT	161.351 54.804 161.383 54.868 ;
			RECT	161.519 54.804 161.551 54.868 ;
			RECT	161.687 54.804 161.719 54.868 ;
			RECT	161.855 54.804 161.887 54.868 ;
			RECT	162.023 54.804 162.055 54.868 ;
			RECT	162.191 54.804 162.223 54.868 ;
			RECT	162.359 54.804 162.391 54.868 ;
			RECT	162.527 54.804 162.559 54.868 ;
			RECT	162.695 54.804 162.727 54.868 ;
			RECT	162.863 54.804 162.895 54.868 ;
			RECT	163.031 54.804 163.063 54.868 ;
			RECT	163.199 54.804 163.231 54.868 ;
			RECT	163.367 54.804 163.399 54.868 ;
			RECT	163.535 54.804 163.567 54.868 ;
			RECT	163.703 54.804 163.735 54.868 ;
			RECT	163.871 54.804 163.903 54.868 ;
			RECT	164.039 54.804 164.071 54.868 ;
			RECT	164.207 54.804 164.239 54.868 ;
			RECT	164.375 54.804 164.407 54.868 ;
			RECT	164.543 54.804 164.575 54.868 ;
			RECT	164.711 54.804 164.743 54.868 ;
			RECT	164.879 54.804 164.911 54.868 ;
			RECT	165.047 54.804 165.079 54.868 ;
			RECT	165.215 54.804 165.247 54.868 ;
			RECT	165.383 54.804 165.415 54.868 ;
			RECT	165.551 54.804 165.583 54.868 ;
			RECT	165.719 54.804 165.751 54.868 ;
			RECT	165.887 54.804 165.919 54.868 ;
			RECT	166.055 54.804 166.087 54.868 ;
			RECT	166.223 54.804 166.255 54.868 ;
			RECT	166.391 54.804 166.423 54.868 ;
			RECT	166.559 54.804 166.591 54.868 ;
			RECT	166.727 54.804 166.759 54.868 ;
			RECT	166.895 54.804 166.927 54.868 ;
			RECT	167.063 54.804 167.095 54.868 ;
			RECT	167.231 54.804 167.263 54.868 ;
			RECT	167.399 54.804 167.431 54.868 ;
			RECT	167.567 54.804 167.599 54.868 ;
			RECT	167.735 54.804 167.767 54.868 ;
			RECT	167.903 54.804 167.935 54.868 ;
			RECT	168.071 54.804 168.103 54.868 ;
			RECT	168.239 54.804 168.271 54.868 ;
			RECT	168.407 54.804 168.439 54.868 ;
			RECT	168.575 54.804 168.607 54.868 ;
			RECT	168.743 54.804 168.775 54.868 ;
			RECT	168.911 54.804 168.943 54.868 ;
			RECT	169.079 54.804 169.111 54.868 ;
			RECT	169.247 54.804 169.279 54.868 ;
			RECT	169.415 54.804 169.447 54.868 ;
			RECT	169.583 54.804 169.615 54.868 ;
			RECT	169.751 54.804 169.783 54.868 ;
			RECT	169.919 54.804 169.951 54.868 ;
			RECT	170.087 54.804 170.119 54.868 ;
			RECT	170.255 54.804 170.287 54.868 ;
			RECT	170.423 54.804 170.455 54.868 ;
			RECT	170.591 54.804 170.623 54.868 ;
			RECT	170.759 54.804 170.791 54.868 ;
			RECT	170.927 54.804 170.959 54.868 ;
			RECT	171.095 54.804 171.127 54.868 ;
			RECT	171.263 54.804 171.295 54.868 ;
			RECT	171.431 54.804 171.463 54.868 ;
			RECT	171.599 54.804 171.631 54.868 ;
			RECT	171.767 54.804 171.799 54.868 ;
			RECT	171.935 54.804 171.967 54.868 ;
			RECT	172.103 54.804 172.135 54.868 ;
			RECT	172.271 54.804 172.303 54.868 ;
			RECT	172.439 54.804 172.471 54.868 ;
			RECT	172.607 54.804 172.639 54.868 ;
			RECT	172.775 54.804 172.807 54.868 ;
			RECT	172.943 54.804 172.975 54.868 ;
			RECT	173.111 54.804 173.143 54.868 ;
			RECT	173.279 54.804 173.311 54.868 ;
			RECT	173.447 54.804 173.479 54.868 ;
			RECT	173.615 54.804 173.647 54.868 ;
			RECT	173.783 54.804 173.815 54.868 ;
			RECT	173.951 54.804 173.983 54.868 ;
			RECT	174.119 54.804 174.151 54.868 ;
			RECT	174.287 54.804 174.319 54.868 ;
			RECT	174.455 54.804 174.487 54.868 ;
			RECT	174.623 54.804 174.655 54.868 ;
			RECT	174.791 54.804 174.823 54.868 ;
			RECT	174.959 54.804 174.991 54.868 ;
			RECT	175.127 54.804 175.159 54.868 ;
			RECT	175.295 54.804 175.327 54.868 ;
			RECT	175.463 54.804 175.495 54.868 ;
			RECT	175.631 54.804 175.663 54.868 ;
			RECT	175.799 54.804 175.831 54.868 ;
			RECT	175.967 54.804 175.999 54.868 ;
			RECT	176.135 54.804 176.167 54.868 ;
			RECT	176.303 54.804 176.335 54.868 ;
			RECT	176.471 54.804 176.503 54.868 ;
			RECT	176.639 54.804 176.671 54.868 ;
			RECT	176.807 54.804 176.839 54.868 ;
			RECT	176.975 54.804 177.007 54.868 ;
			RECT	177.143 54.804 177.175 54.868 ;
			RECT	177.311 54.804 177.343 54.868 ;
			RECT	177.479 54.804 177.511 54.868 ;
			RECT	177.647 54.804 177.679 54.868 ;
			RECT	177.815 54.804 177.847 54.868 ;
			RECT	177.983 54.804 178.015 54.868 ;
			RECT	178.151 54.804 178.183 54.868 ;
			RECT	178.319 54.804 178.351 54.868 ;
			RECT	178.487 54.804 178.519 54.868 ;
			RECT	178.655 54.804 178.687 54.868 ;
			RECT	178.823 54.804 178.855 54.868 ;
			RECT	178.991 54.804 179.023 54.868 ;
			RECT	179.159 54.804 179.191 54.868 ;
			RECT	179.327 54.804 179.359 54.868 ;
			RECT	179.495 54.804 179.527 54.868 ;
			RECT	179.663 54.804 179.695 54.868 ;
			RECT	179.831 54.804 179.863 54.868 ;
			RECT	179.999 54.804 180.031 54.868 ;
			RECT	180.167 54.804 180.199 54.868 ;
			RECT	180.335 54.804 180.367 54.868 ;
			RECT	180.503 54.804 180.535 54.868 ;
			RECT	180.671 54.804 180.703 54.868 ;
			RECT	180.839 54.804 180.871 54.868 ;
			RECT	181.007 54.804 181.039 54.868 ;
			RECT	181.175 54.804 181.207 54.868 ;
			RECT	181.343 54.804 181.375 54.868 ;
			RECT	181.511 54.804 181.543 54.868 ;
			RECT	181.679 54.804 181.711 54.868 ;
			RECT	181.847 54.804 181.879 54.868 ;
			RECT	182.015 54.804 182.047 54.868 ;
			RECT	182.183 54.804 182.215 54.868 ;
			RECT	182.351 54.804 182.383 54.868 ;
			RECT	182.519 54.804 182.551 54.868 ;
			RECT	182.687 54.804 182.719 54.868 ;
			RECT	182.855 54.804 182.887 54.868 ;
			RECT	183.023 54.804 183.055 54.868 ;
			RECT	183.191 54.804 183.223 54.868 ;
			RECT	183.359 54.804 183.391 54.868 ;
			RECT	183.527 54.804 183.559 54.868 ;
			RECT	183.695 54.804 183.727 54.868 ;
			RECT	183.863 54.804 183.895 54.868 ;
			RECT	184.031 54.804 184.063 54.868 ;
			RECT	184.199 54.804 184.231 54.868 ;
			RECT	184.367 54.804 184.399 54.868 ;
			RECT	184.535 54.804 184.567 54.868 ;
			RECT	184.703 54.804 184.735 54.868 ;
			RECT	184.871 54.804 184.903 54.868 ;
			RECT	185.039 54.804 185.071 54.868 ;
			RECT	185.207 54.804 185.239 54.868 ;
			RECT	185.375 54.804 185.407 54.868 ;
			RECT	185.543 54.804 185.575 54.868 ;
			RECT	185.711 54.804 185.743 54.868 ;
			RECT	185.879 54.804 185.911 54.868 ;
			RECT	186.047 54.804 186.079 54.868 ;
			RECT	186.215 54.804 186.247 54.868 ;
			RECT	186.383 54.804 186.415 54.868 ;
			RECT	186.551 54.804 186.583 54.868 ;
			RECT	186.719 54.804 186.751 54.868 ;
			RECT	186.887 54.804 186.919 54.868 ;
			RECT	187.055 54.804 187.087 54.868 ;
			RECT	187.223 54.804 187.255 54.868 ;
			RECT	187.391 54.804 187.423 54.868 ;
			RECT	187.559 54.804 187.591 54.868 ;
			RECT	187.727 54.804 187.759 54.868 ;
			RECT	187.895 54.804 187.927 54.868 ;
			RECT	188.063 54.804 188.095 54.868 ;
			RECT	188.231 54.804 188.263 54.868 ;
			RECT	188.399 54.804 188.431 54.868 ;
			RECT	188.567 54.804 188.599 54.868 ;
			RECT	188.735 54.804 188.767 54.868 ;
			RECT	188.903 54.804 188.935 54.868 ;
			RECT	189.071 54.804 189.103 54.868 ;
			RECT	189.239 54.804 189.271 54.868 ;
			RECT	189.407 54.804 189.439 54.868 ;
			RECT	189.575 54.804 189.607 54.868 ;
			RECT	189.743 54.804 189.775 54.868 ;
			RECT	189.911 54.804 189.943 54.868 ;
			RECT	190.079 54.804 190.111 54.868 ;
			RECT	190.247 54.804 190.279 54.868 ;
			RECT	190.415 54.804 190.447 54.868 ;
			RECT	190.583 54.804 190.615 54.868 ;
			RECT	190.751 54.804 190.783 54.868 ;
			RECT	190.919 54.804 190.951 54.868 ;
			RECT	191.087 54.804 191.119 54.868 ;
			RECT	191.255 54.804 191.287 54.868 ;
			RECT	191.423 54.804 191.455 54.868 ;
			RECT	191.591 54.804 191.623 54.868 ;
			RECT	191.759 54.804 191.791 54.868 ;
			RECT	191.927 54.804 191.959 54.868 ;
			RECT	192.095 54.804 192.127 54.868 ;
			RECT	192.263 54.804 192.295 54.868 ;
			RECT	192.431 54.804 192.463 54.868 ;
			RECT	192.599 54.804 192.631 54.868 ;
			RECT	192.767 54.804 192.799 54.868 ;
			RECT	192.935 54.804 192.967 54.868 ;
			RECT	193.103 54.804 193.135 54.868 ;
			RECT	193.271 54.804 193.303 54.868 ;
			RECT	193.439 54.804 193.471 54.868 ;
			RECT	193.607 54.804 193.639 54.868 ;
			RECT	193.775 54.804 193.807 54.868 ;
			RECT	193.943 54.804 193.975 54.868 ;
			RECT	194.111 54.804 194.143 54.868 ;
			RECT	194.279 54.804 194.311 54.868 ;
			RECT	194.447 54.804 194.479 54.868 ;
			RECT	194.615 54.804 194.647 54.868 ;
			RECT	194.783 54.804 194.815 54.868 ;
			RECT	194.951 54.804 194.983 54.868 ;
			RECT	195.119 54.804 195.151 54.868 ;
			RECT	195.287 54.804 195.319 54.868 ;
			RECT	195.455 54.804 195.487 54.868 ;
			RECT	195.623 54.804 195.655 54.868 ;
			RECT	195.791 54.804 195.823 54.868 ;
			RECT	195.959 54.804 195.991 54.868 ;
			RECT	196.127 54.804 196.159 54.868 ;
			RECT	196.295 54.804 196.327 54.868 ;
			RECT	196.463 54.804 196.495 54.868 ;
			RECT	196.631 54.804 196.663 54.868 ;
			RECT	196.799 54.804 196.831 54.868 ;
			RECT	196.967 54.804 196.999 54.868 ;
			RECT	197.135 54.804 197.167 54.868 ;
			RECT	197.303 54.804 197.335 54.868 ;
			RECT	197.471 54.804 197.503 54.868 ;
			RECT	197.639 54.804 197.671 54.868 ;
			RECT	197.807 54.804 197.839 54.868 ;
			RECT	197.975 54.804 198.007 54.868 ;
			RECT	198.143 54.804 198.175 54.868 ;
			RECT	198.311 54.804 198.343 54.868 ;
			RECT	198.479 54.804 198.511 54.868 ;
			RECT	198.647 54.804 198.679 54.868 ;
			RECT	198.815 54.804 198.847 54.868 ;
			RECT	198.983 54.804 199.015 54.868 ;
			RECT	199.151 54.804 199.183 54.868 ;
			RECT	199.319 54.804 199.351 54.868 ;
			RECT	199.487 54.804 199.519 54.868 ;
			RECT	199.655 54.804 199.687 54.868 ;
			RECT	199.823 54.804 199.855 54.868 ;
			RECT	199.991 54.804 200.023 54.868 ;
			RECT	200.121 54.82 200.153 54.852 ;
			RECT	200.243 54.815 200.275 54.847 ;
			RECT	200.373 54.804 200.405 54.868 ;
			RECT	200.9 54.804 200.932 54.868 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 52.856 201.665 52.976 ;
			LAYER	J3 ;
			RECT	0.755 52.884 0.787 52.948 ;
			RECT	1.645 52.884 1.709 52.948 ;
			RECT	2.323 52.884 2.387 52.948 ;
			RECT	3.438 52.884 3.47 52.948 ;
			RECT	3.585 52.884 3.617 52.948 ;
			RECT	4.195 52.884 4.227 52.948 ;
			RECT	4.72 52.884 4.752 52.948 ;
			RECT	4.944 52.884 5.008 52.948 ;
			RECT	5.267 52.884 5.299 52.948 ;
			RECT	5.797 52.884 5.829 52.948 ;
			RECT	5.927 52.895 5.959 52.927 ;
			RECT	6.049 52.9 6.081 52.932 ;
			RECT	6.179 52.884 6.211 52.948 ;
			RECT	6.347 52.884 6.379 52.948 ;
			RECT	6.515 52.884 6.547 52.948 ;
			RECT	6.683 52.884 6.715 52.948 ;
			RECT	6.851 52.884 6.883 52.948 ;
			RECT	7.019 52.884 7.051 52.948 ;
			RECT	7.187 52.884 7.219 52.948 ;
			RECT	7.355 52.884 7.387 52.948 ;
			RECT	7.523 52.884 7.555 52.948 ;
			RECT	7.691 52.884 7.723 52.948 ;
			RECT	7.859 52.884 7.891 52.948 ;
			RECT	8.027 52.884 8.059 52.948 ;
			RECT	8.195 52.884 8.227 52.948 ;
			RECT	8.363 52.884 8.395 52.948 ;
			RECT	8.531 52.884 8.563 52.948 ;
			RECT	8.699 52.884 8.731 52.948 ;
			RECT	8.867 52.884 8.899 52.948 ;
			RECT	9.035 52.884 9.067 52.948 ;
			RECT	9.203 52.884 9.235 52.948 ;
			RECT	9.371 52.884 9.403 52.948 ;
			RECT	9.539 52.884 9.571 52.948 ;
			RECT	9.707 52.884 9.739 52.948 ;
			RECT	9.875 52.884 9.907 52.948 ;
			RECT	10.043 52.884 10.075 52.948 ;
			RECT	10.211 52.884 10.243 52.948 ;
			RECT	10.379 52.884 10.411 52.948 ;
			RECT	10.547 52.884 10.579 52.948 ;
			RECT	10.715 52.884 10.747 52.948 ;
			RECT	10.883 52.884 10.915 52.948 ;
			RECT	11.051 52.884 11.083 52.948 ;
			RECT	11.219 52.884 11.251 52.948 ;
			RECT	11.387 52.884 11.419 52.948 ;
			RECT	11.555 52.884 11.587 52.948 ;
			RECT	11.723 52.884 11.755 52.948 ;
			RECT	11.891 52.884 11.923 52.948 ;
			RECT	12.059 52.884 12.091 52.948 ;
			RECT	12.227 52.884 12.259 52.948 ;
			RECT	12.395 52.884 12.427 52.948 ;
			RECT	12.563 52.884 12.595 52.948 ;
			RECT	12.731 52.884 12.763 52.948 ;
			RECT	12.899 52.884 12.931 52.948 ;
			RECT	13.067 52.884 13.099 52.948 ;
			RECT	13.235 52.884 13.267 52.948 ;
			RECT	13.403 52.884 13.435 52.948 ;
			RECT	13.571 52.884 13.603 52.948 ;
			RECT	13.739 52.884 13.771 52.948 ;
			RECT	13.907 52.884 13.939 52.948 ;
			RECT	14.075 52.884 14.107 52.948 ;
			RECT	14.243 52.884 14.275 52.948 ;
			RECT	14.411 52.884 14.443 52.948 ;
			RECT	14.579 52.884 14.611 52.948 ;
			RECT	14.747 52.884 14.779 52.948 ;
			RECT	14.915 52.884 14.947 52.948 ;
			RECT	15.083 52.884 15.115 52.948 ;
			RECT	15.251 52.884 15.283 52.948 ;
			RECT	15.419 52.884 15.451 52.948 ;
			RECT	15.587 52.884 15.619 52.948 ;
			RECT	15.755 52.884 15.787 52.948 ;
			RECT	15.923 52.884 15.955 52.948 ;
			RECT	16.091 52.884 16.123 52.948 ;
			RECT	16.259 52.884 16.291 52.948 ;
			RECT	16.427 52.884 16.459 52.948 ;
			RECT	16.595 52.884 16.627 52.948 ;
			RECT	16.763 52.884 16.795 52.948 ;
			RECT	16.931 52.884 16.963 52.948 ;
			RECT	17.099 52.884 17.131 52.948 ;
			RECT	17.267 52.884 17.299 52.948 ;
			RECT	17.435 52.884 17.467 52.948 ;
			RECT	17.603 52.884 17.635 52.948 ;
			RECT	17.771 52.884 17.803 52.948 ;
			RECT	17.939 52.884 17.971 52.948 ;
			RECT	18.107 52.884 18.139 52.948 ;
			RECT	18.275 52.884 18.307 52.948 ;
			RECT	18.443 52.884 18.475 52.948 ;
			RECT	18.611 52.884 18.643 52.948 ;
			RECT	18.779 52.884 18.811 52.948 ;
			RECT	18.947 52.884 18.979 52.948 ;
			RECT	19.115 52.884 19.147 52.948 ;
			RECT	19.283 52.884 19.315 52.948 ;
			RECT	19.451 52.884 19.483 52.948 ;
			RECT	19.619 52.884 19.651 52.948 ;
			RECT	19.787 52.884 19.819 52.948 ;
			RECT	19.955 52.884 19.987 52.948 ;
			RECT	20.123 52.884 20.155 52.948 ;
			RECT	20.291 52.884 20.323 52.948 ;
			RECT	20.459 52.884 20.491 52.948 ;
			RECT	20.627 52.884 20.659 52.948 ;
			RECT	20.795 52.884 20.827 52.948 ;
			RECT	20.963 52.884 20.995 52.948 ;
			RECT	21.131 52.884 21.163 52.948 ;
			RECT	21.299 52.884 21.331 52.948 ;
			RECT	21.467 52.884 21.499 52.948 ;
			RECT	21.635 52.884 21.667 52.948 ;
			RECT	21.803 52.884 21.835 52.948 ;
			RECT	21.971 52.884 22.003 52.948 ;
			RECT	22.139 52.884 22.171 52.948 ;
			RECT	22.307 52.884 22.339 52.948 ;
			RECT	22.475 52.884 22.507 52.948 ;
			RECT	22.643 52.884 22.675 52.948 ;
			RECT	22.811 52.884 22.843 52.948 ;
			RECT	22.979 52.884 23.011 52.948 ;
			RECT	23.147 52.884 23.179 52.948 ;
			RECT	23.315 52.884 23.347 52.948 ;
			RECT	23.483 52.884 23.515 52.948 ;
			RECT	23.651 52.884 23.683 52.948 ;
			RECT	23.819 52.884 23.851 52.948 ;
			RECT	23.987 52.884 24.019 52.948 ;
			RECT	24.155 52.884 24.187 52.948 ;
			RECT	24.323 52.884 24.355 52.948 ;
			RECT	24.491 52.884 24.523 52.948 ;
			RECT	24.659 52.884 24.691 52.948 ;
			RECT	24.827 52.884 24.859 52.948 ;
			RECT	24.995 52.884 25.027 52.948 ;
			RECT	25.163 52.884 25.195 52.948 ;
			RECT	25.331 52.884 25.363 52.948 ;
			RECT	25.499 52.884 25.531 52.948 ;
			RECT	25.667 52.884 25.699 52.948 ;
			RECT	25.835 52.884 25.867 52.948 ;
			RECT	26.003 52.884 26.035 52.948 ;
			RECT	26.171 52.884 26.203 52.948 ;
			RECT	26.339 52.884 26.371 52.948 ;
			RECT	26.507 52.884 26.539 52.948 ;
			RECT	26.675 52.884 26.707 52.948 ;
			RECT	26.843 52.884 26.875 52.948 ;
			RECT	27.011 52.884 27.043 52.948 ;
			RECT	27.179 52.884 27.211 52.948 ;
			RECT	27.347 52.884 27.379 52.948 ;
			RECT	27.515 52.884 27.547 52.948 ;
			RECT	27.683 52.884 27.715 52.948 ;
			RECT	27.851 52.884 27.883 52.948 ;
			RECT	28.019 52.884 28.051 52.948 ;
			RECT	28.187 52.884 28.219 52.948 ;
			RECT	28.355 52.884 28.387 52.948 ;
			RECT	28.523 52.884 28.555 52.948 ;
			RECT	28.691 52.884 28.723 52.948 ;
			RECT	28.859 52.884 28.891 52.948 ;
			RECT	29.027 52.884 29.059 52.948 ;
			RECT	29.195 52.884 29.227 52.948 ;
			RECT	29.363 52.884 29.395 52.948 ;
			RECT	29.531 52.884 29.563 52.948 ;
			RECT	29.699 52.884 29.731 52.948 ;
			RECT	29.867 52.884 29.899 52.948 ;
			RECT	30.035 52.884 30.067 52.948 ;
			RECT	30.203 52.884 30.235 52.948 ;
			RECT	30.371 52.884 30.403 52.948 ;
			RECT	30.539 52.884 30.571 52.948 ;
			RECT	30.707 52.884 30.739 52.948 ;
			RECT	30.875 52.884 30.907 52.948 ;
			RECT	31.043 52.884 31.075 52.948 ;
			RECT	31.211 52.884 31.243 52.948 ;
			RECT	31.379 52.884 31.411 52.948 ;
			RECT	31.547 52.884 31.579 52.948 ;
			RECT	31.715 52.884 31.747 52.948 ;
			RECT	31.883 52.884 31.915 52.948 ;
			RECT	32.051 52.884 32.083 52.948 ;
			RECT	32.219 52.884 32.251 52.948 ;
			RECT	32.387 52.884 32.419 52.948 ;
			RECT	32.555 52.884 32.587 52.948 ;
			RECT	32.723 52.884 32.755 52.948 ;
			RECT	32.891 52.884 32.923 52.948 ;
			RECT	33.059 52.884 33.091 52.948 ;
			RECT	33.227 52.884 33.259 52.948 ;
			RECT	33.395 52.884 33.427 52.948 ;
			RECT	33.563 52.884 33.595 52.948 ;
			RECT	33.731 52.884 33.763 52.948 ;
			RECT	33.899 52.884 33.931 52.948 ;
			RECT	34.067 52.884 34.099 52.948 ;
			RECT	34.235 52.884 34.267 52.948 ;
			RECT	34.403 52.884 34.435 52.948 ;
			RECT	34.571 52.884 34.603 52.948 ;
			RECT	34.739 52.884 34.771 52.948 ;
			RECT	34.907 52.884 34.939 52.948 ;
			RECT	35.075 52.884 35.107 52.948 ;
			RECT	35.243 52.884 35.275 52.948 ;
			RECT	35.411 52.884 35.443 52.948 ;
			RECT	35.579 52.884 35.611 52.948 ;
			RECT	35.747 52.884 35.779 52.948 ;
			RECT	35.915 52.884 35.947 52.948 ;
			RECT	36.083 52.884 36.115 52.948 ;
			RECT	36.251 52.884 36.283 52.948 ;
			RECT	36.419 52.884 36.451 52.948 ;
			RECT	36.587 52.884 36.619 52.948 ;
			RECT	36.755 52.884 36.787 52.948 ;
			RECT	36.923 52.884 36.955 52.948 ;
			RECT	37.091 52.884 37.123 52.948 ;
			RECT	37.259 52.884 37.291 52.948 ;
			RECT	37.427 52.884 37.459 52.948 ;
			RECT	37.595 52.884 37.627 52.948 ;
			RECT	37.763 52.884 37.795 52.948 ;
			RECT	37.931 52.884 37.963 52.948 ;
			RECT	38.099 52.884 38.131 52.948 ;
			RECT	38.267 52.884 38.299 52.948 ;
			RECT	38.435 52.884 38.467 52.948 ;
			RECT	38.603 52.884 38.635 52.948 ;
			RECT	38.771 52.884 38.803 52.948 ;
			RECT	38.939 52.884 38.971 52.948 ;
			RECT	39.107 52.884 39.139 52.948 ;
			RECT	39.275 52.884 39.307 52.948 ;
			RECT	39.443 52.884 39.475 52.948 ;
			RECT	39.611 52.884 39.643 52.948 ;
			RECT	39.779 52.884 39.811 52.948 ;
			RECT	39.947 52.884 39.979 52.948 ;
			RECT	40.115 52.884 40.147 52.948 ;
			RECT	40.283 52.884 40.315 52.948 ;
			RECT	40.451 52.884 40.483 52.948 ;
			RECT	40.619 52.884 40.651 52.948 ;
			RECT	40.787 52.884 40.819 52.948 ;
			RECT	40.955 52.884 40.987 52.948 ;
			RECT	41.123 52.884 41.155 52.948 ;
			RECT	41.291 52.884 41.323 52.948 ;
			RECT	41.459 52.884 41.491 52.948 ;
			RECT	41.627 52.884 41.659 52.948 ;
			RECT	41.795 52.884 41.827 52.948 ;
			RECT	41.963 52.884 41.995 52.948 ;
			RECT	42.131 52.884 42.163 52.948 ;
			RECT	42.299 52.884 42.331 52.948 ;
			RECT	42.467 52.884 42.499 52.948 ;
			RECT	42.635 52.884 42.667 52.948 ;
			RECT	42.803 52.884 42.835 52.948 ;
			RECT	42.971 52.884 43.003 52.948 ;
			RECT	43.139 52.884 43.171 52.948 ;
			RECT	43.307 52.884 43.339 52.948 ;
			RECT	43.475 52.884 43.507 52.948 ;
			RECT	43.643 52.884 43.675 52.948 ;
			RECT	43.811 52.884 43.843 52.948 ;
			RECT	43.979 52.884 44.011 52.948 ;
			RECT	44.147 52.884 44.179 52.948 ;
			RECT	44.315 52.884 44.347 52.948 ;
			RECT	44.483 52.884 44.515 52.948 ;
			RECT	44.651 52.884 44.683 52.948 ;
			RECT	44.819 52.884 44.851 52.948 ;
			RECT	44.987 52.884 45.019 52.948 ;
			RECT	45.155 52.884 45.187 52.948 ;
			RECT	45.323 52.884 45.355 52.948 ;
			RECT	45.491 52.884 45.523 52.948 ;
			RECT	45.659 52.884 45.691 52.948 ;
			RECT	45.827 52.884 45.859 52.948 ;
			RECT	45.995 52.884 46.027 52.948 ;
			RECT	46.163 52.884 46.195 52.948 ;
			RECT	46.331 52.884 46.363 52.948 ;
			RECT	46.499 52.884 46.531 52.948 ;
			RECT	46.667 52.884 46.699 52.948 ;
			RECT	46.835 52.884 46.867 52.948 ;
			RECT	47.003 52.884 47.035 52.948 ;
			RECT	47.171 52.884 47.203 52.948 ;
			RECT	47.339 52.884 47.371 52.948 ;
			RECT	47.507 52.884 47.539 52.948 ;
			RECT	47.675 52.884 47.707 52.948 ;
			RECT	47.843 52.884 47.875 52.948 ;
			RECT	48.011 52.884 48.043 52.948 ;
			RECT	48.179 52.884 48.211 52.948 ;
			RECT	48.347 52.884 48.379 52.948 ;
			RECT	48.515 52.884 48.547 52.948 ;
			RECT	48.683 52.884 48.715 52.948 ;
			RECT	48.851 52.884 48.883 52.948 ;
			RECT	49.019 52.884 49.051 52.948 ;
			RECT	49.187 52.884 49.219 52.948 ;
			RECT	49.318 52.9 49.35 52.932 ;
			RECT	49.439 52.9 49.471 52.932 ;
			RECT	49.569 52.884 49.601 52.948 ;
			RECT	51.881 52.884 51.913 52.948 ;
			RECT	53.132 52.884 53.196 52.948 ;
			RECT	53.812 52.884 53.844 52.948 ;
			RECT	54.251 52.884 54.283 52.948 ;
			RECT	55.562 52.884 55.626 52.948 ;
			RECT	58.603 52.884 58.635 52.948 ;
			RECT	58.733 52.9 58.765 52.932 ;
			RECT	58.854 52.9 58.886 52.932 ;
			RECT	58.985 52.884 59.017 52.948 ;
			RECT	59.153 52.884 59.185 52.948 ;
			RECT	59.321 52.884 59.353 52.948 ;
			RECT	59.489 52.884 59.521 52.948 ;
			RECT	59.657 52.884 59.689 52.948 ;
			RECT	59.825 52.884 59.857 52.948 ;
			RECT	59.993 52.884 60.025 52.948 ;
			RECT	60.161 52.884 60.193 52.948 ;
			RECT	60.329 52.884 60.361 52.948 ;
			RECT	60.497 52.884 60.529 52.948 ;
			RECT	60.665 52.884 60.697 52.948 ;
			RECT	60.833 52.884 60.865 52.948 ;
			RECT	61.001 52.884 61.033 52.948 ;
			RECT	61.169 52.884 61.201 52.948 ;
			RECT	61.337 52.884 61.369 52.948 ;
			RECT	61.505 52.884 61.537 52.948 ;
			RECT	61.673 52.884 61.705 52.948 ;
			RECT	61.841 52.884 61.873 52.948 ;
			RECT	62.009 52.884 62.041 52.948 ;
			RECT	62.177 52.884 62.209 52.948 ;
			RECT	62.345 52.884 62.377 52.948 ;
			RECT	62.513 52.884 62.545 52.948 ;
			RECT	62.681 52.884 62.713 52.948 ;
			RECT	62.849 52.884 62.881 52.948 ;
			RECT	63.017 52.884 63.049 52.948 ;
			RECT	63.185 52.884 63.217 52.948 ;
			RECT	63.353 52.884 63.385 52.948 ;
			RECT	63.521 52.884 63.553 52.948 ;
			RECT	63.689 52.884 63.721 52.948 ;
			RECT	63.857 52.884 63.889 52.948 ;
			RECT	64.025 52.884 64.057 52.948 ;
			RECT	64.193 52.884 64.225 52.948 ;
			RECT	64.361 52.884 64.393 52.948 ;
			RECT	64.529 52.884 64.561 52.948 ;
			RECT	64.697 52.884 64.729 52.948 ;
			RECT	64.865 52.884 64.897 52.948 ;
			RECT	65.033 52.884 65.065 52.948 ;
			RECT	65.201 52.884 65.233 52.948 ;
			RECT	65.369 52.884 65.401 52.948 ;
			RECT	65.537 52.884 65.569 52.948 ;
			RECT	65.705 52.884 65.737 52.948 ;
			RECT	65.873 52.884 65.905 52.948 ;
			RECT	66.041 52.884 66.073 52.948 ;
			RECT	66.209 52.884 66.241 52.948 ;
			RECT	66.377 52.884 66.409 52.948 ;
			RECT	66.545 52.884 66.577 52.948 ;
			RECT	66.713 52.884 66.745 52.948 ;
			RECT	66.881 52.884 66.913 52.948 ;
			RECT	67.049 52.884 67.081 52.948 ;
			RECT	67.217 52.884 67.249 52.948 ;
			RECT	67.385 52.884 67.417 52.948 ;
			RECT	67.553 52.884 67.585 52.948 ;
			RECT	67.721 52.884 67.753 52.948 ;
			RECT	67.889 52.884 67.921 52.948 ;
			RECT	68.057 52.884 68.089 52.948 ;
			RECT	68.225 52.884 68.257 52.948 ;
			RECT	68.393 52.884 68.425 52.948 ;
			RECT	68.561 52.884 68.593 52.948 ;
			RECT	68.729 52.884 68.761 52.948 ;
			RECT	68.897 52.884 68.929 52.948 ;
			RECT	69.065 52.884 69.097 52.948 ;
			RECT	69.233 52.884 69.265 52.948 ;
			RECT	69.401 52.884 69.433 52.948 ;
			RECT	69.569 52.884 69.601 52.948 ;
			RECT	69.737 52.884 69.769 52.948 ;
			RECT	69.905 52.884 69.937 52.948 ;
			RECT	70.073 52.884 70.105 52.948 ;
			RECT	70.241 52.884 70.273 52.948 ;
			RECT	70.409 52.884 70.441 52.948 ;
			RECT	70.577 52.884 70.609 52.948 ;
			RECT	70.745 52.884 70.777 52.948 ;
			RECT	70.913 52.884 70.945 52.948 ;
			RECT	71.081 52.884 71.113 52.948 ;
			RECT	71.249 52.884 71.281 52.948 ;
			RECT	71.417 52.884 71.449 52.948 ;
			RECT	71.585 52.884 71.617 52.948 ;
			RECT	71.753 52.884 71.785 52.948 ;
			RECT	71.921 52.884 71.953 52.948 ;
			RECT	72.089 52.884 72.121 52.948 ;
			RECT	72.257 52.884 72.289 52.948 ;
			RECT	72.425 52.884 72.457 52.948 ;
			RECT	72.593 52.884 72.625 52.948 ;
			RECT	72.761 52.884 72.793 52.948 ;
			RECT	72.929 52.884 72.961 52.948 ;
			RECT	73.097 52.884 73.129 52.948 ;
			RECT	73.265 52.884 73.297 52.948 ;
			RECT	73.433 52.884 73.465 52.948 ;
			RECT	73.601 52.884 73.633 52.948 ;
			RECT	73.769 52.884 73.801 52.948 ;
			RECT	73.937 52.884 73.969 52.948 ;
			RECT	74.105 52.884 74.137 52.948 ;
			RECT	74.273 52.884 74.305 52.948 ;
			RECT	74.441 52.884 74.473 52.948 ;
			RECT	74.609 52.884 74.641 52.948 ;
			RECT	74.777 52.884 74.809 52.948 ;
			RECT	74.945 52.884 74.977 52.948 ;
			RECT	75.113 52.884 75.145 52.948 ;
			RECT	75.281 52.884 75.313 52.948 ;
			RECT	75.449 52.884 75.481 52.948 ;
			RECT	75.617 52.884 75.649 52.948 ;
			RECT	75.785 52.884 75.817 52.948 ;
			RECT	75.953 52.884 75.985 52.948 ;
			RECT	76.121 52.884 76.153 52.948 ;
			RECT	76.289 52.884 76.321 52.948 ;
			RECT	76.457 52.884 76.489 52.948 ;
			RECT	76.625 52.884 76.657 52.948 ;
			RECT	76.793 52.884 76.825 52.948 ;
			RECT	76.961 52.884 76.993 52.948 ;
			RECT	77.129 52.884 77.161 52.948 ;
			RECT	77.297 52.884 77.329 52.948 ;
			RECT	77.465 52.884 77.497 52.948 ;
			RECT	77.633 52.884 77.665 52.948 ;
			RECT	77.801 52.884 77.833 52.948 ;
			RECT	77.969 52.884 78.001 52.948 ;
			RECT	78.137 52.884 78.169 52.948 ;
			RECT	78.305 52.884 78.337 52.948 ;
			RECT	78.473 52.884 78.505 52.948 ;
			RECT	78.641 52.884 78.673 52.948 ;
			RECT	78.809 52.884 78.841 52.948 ;
			RECT	78.977 52.884 79.009 52.948 ;
			RECT	79.145 52.884 79.177 52.948 ;
			RECT	79.313 52.884 79.345 52.948 ;
			RECT	79.481 52.884 79.513 52.948 ;
			RECT	79.649 52.884 79.681 52.948 ;
			RECT	79.817 52.884 79.849 52.948 ;
			RECT	79.985 52.884 80.017 52.948 ;
			RECT	80.153 52.884 80.185 52.948 ;
			RECT	80.321 52.884 80.353 52.948 ;
			RECT	80.489 52.884 80.521 52.948 ;
			RECT	80.657 52.884 80.689 52.948 ;
			RECT	80.825 52.884 80.857 52.948 ;
			RECT	80.993 52.884 81.025 52.948 ;
			RECT	81.161 52.884 81.193 52.948 ;
			RECT	81.329 52.884 81.361 52.948 ;
			RECT	81.497 52.884 81.529 52.948 ;
			RECT	81.665 52.884 81.697 52.948 ;
			RECT	81.833 52.884 81.865 52.948 ;
			RECT	82.001 52.884 82.033 52.948 ;
			RECT	82.169 52.884 82.201 52.948 ;
			RECT	82.337 52.884 82.369 52.948 ;
			RECT	82.505 52.884 82.537 52.948 ;
			RECT	82.673 52.884 82.705 52.948 ;
			RECT	82.841 52.884 82.873 52.948 ;
			RECT	83.009 52.884 83.041 52.948 ;
			RECT	83.177 52.884 83.209 52.948 ;
			RECT	83.345 52.884 83.377 52.948 ;
			RECT	83.513 52.884 83.545 52.948 ;
			RECT	83.681 52.884 83.713 52.948 ;
			RECT	83.849 52.884 83.881 52.948 ;
			RECT	84.017 52.884 84.049 52.948 ;
			RECT	84.185 52.884 84.217 52.948 ;
			RECT	84.353 52.884 84.385 52.948 ;
			RECT	84.521 52.884 84.553 52.948 ;
			RECT	84.689 52.884 84.721 52.948 ;
			RECT	84.857 52.884 84.889 52.948 ;
			RECT	85.025 52.884 85.057 52.948 ;
			RECT	85.193 52.884 85.225 52.948 ;
			RECT	85.361 52.884 85.393 52.948 ;
			RECT	85.529 52.884 85.561 52.948 ;
			RECT	85.697 52.884 85.729 52.948 ;
			RECT	85.865 52.884 85.897 52.948 ;
			RECT	86.033 52.884 86.065 52.948 ;
			RECT	86.201 52.884 86.233 52.948 ;
			RECT	86.369 52.884 86.401 52.948 ;
			RECT	86.537 52.884 86.569 52.948 ;
			RECT	86.705 52.884 86.737 52.948 ;
			RECT	86.873 52.884 86.905 52.948 ;
			RECT	87.041 52.884 87.073 52.948 ;
			RECT	87.209 52.884 87.241 52.948 ;
			RECT	87.377 52.884 87.409 52.948 ;
			RECT	87.545 52.884 87.577 52.948 ;
			RECT	87.713 52.884 87.745 52.948 ;
			RECT	87.881 52.884 87.913 52.948 ;
			RECT	88.049 52.884 88.081 52.948 ;
			RECT	88.217 52.884 88.249 52.948 ;
			RECT	88.385 52.884 88.417 52.948 ;
			RECT	88.553 52.884 88.585 52.948 ;
			RECT	88.721 52.884 88.753 52.948 ;
			RECT	88.889 52.884 88.921 52.948 ;
			RECT	89.057 52.884 89.089 52.948 ;
			RECT	89.225 52.884 89.257 52.948 ;
			RECT	89.393 52.884 89.425 52.948 ;
			RECT	89.561 52.884 89.593 52.948 ;
			RECT	89.729 52.884 89.761 52.948 ;
			RECT	89.897 52.884 89.929 52.948 ;
			RECT	90.065 52.884 90.097 52.948 ;
			RECT	90.233 52.884 90.265 52.948 ;
			RECT	90.401 52.884 90.433 52.948 ;
			RECT	90.569 52.884 90.601 52.948 ;
			RECT	90.737 52.884 90.769 52.948 ;
			RECT	90.905 52.884 90.937 52.948 ;
			RECT	91.073 52.884 91.105 52.948 ;
			RECT	91.241 52.884 91.273 52.948 ;
			RECT	91.409 52.884 91.441 52.948 ;
			RECT	91.577 52.884 91.609 52.948 ;
			RECT	91.745 52.884 91.777 52.948 ;
			RECT	91.913 52.884 91.945 52.948 ;
			RECT	92.081 52.884 92.113 52.948 ;
			RECT	92.249 52.884 92.281 52.948 ;
			RECT	92.417 52.884 92.449 52.948 ;
			RECT	92.585 52.884 92.617 52.948 ;
			RECT	92.753 52.884 92.785 52.948 ;
			RECT	92.921 52.884 92.953 52.948 ;
			RECT	93.089 52.884 93.121 52.948 ;
			RECT	93.257 52.884 93.289 52.948 ;
			RECT	93.425 52.884 93.457 52.948 ;
			RECT	93.593 52.884 93.625 52.948 ;
			RECT	93.761 52.884 93.793 52.948 ;
			RECT	93.929 52.884 93.961 52.948 ;
			RECT	94.097 52.884 94.129 52.948 ;
			RECT	94.265 52.884 94.297 52.948 ;
			RECT	94.433 52.884 94.465 52.948 ;
			RECT	94.601 52.884 94.633 52.948 ;
			RECT	94.769 52.884 94.801 52.948 ;
			RECT	94.937 52.884 94.969 52.948 ;
			RECT	95.105 52.884 95.137 52.948 ;
			RECT	95.273 52.884 95.305 52.948 ;
			RECT	95.441 52.884 95.473 52.948 ;
			RECT	95.609 52.884 95.641 52.948 ;
			RECT	95.777 52.884 95.809 52.948 ;
			RECT	95.945 52.884 95.977 52.948 ;
			RECT	96.113 52.884 96.145 52.948 ;
			RECT	96.281 52.884 96.313 52.948 ;
			RECT	96.449 52.884 96.481 52.948 ;
			RECT	96.617 52.884 96.649 52.948 ;
			RECT	96.785 52.884 96.817 52.948 ;
			RECT	96.953 52.884 96.985 52.948 ;
			RECT	97.121 52.884 97.153 52.948 ;
			RECT	97.289 52.884 97.321 52.948 ;
			RECT	97.457 52.884 97.489 52.948 ;
			RECT	97.625 52.884 97.657 52.948 ;
			RECT	97.793 52.884 97.825 52.948 ;
			RECT	97.961 52.884 97.993 52.948 ;
			RECT	98.129 52.884 98.161 52.948 ;
			RECT	98.297 52.884 98.329 52.948 ;
			RECT	98.465 52.884 98.497 52.948 ;
			RECT	98.633 52.884 98.665 52.948 ;
			RECT	98.801 52.884 98.833 52.948 ;
			RECT	98.969 52.884 99.001 52.948 ;
			RECT	99.137 52.884 99.169 52.948 ;
			RECT	99.305 52.884 99.337 52.948 ;
			RECT	99.473 52.884 99.505 52.948 ;
			RECT	99.641 52.884 99.673 52.948 ;
			RECT	99.809 52.884 99.841 52.948 ;
			RECT	99.977 52.884 100.009 52.948 ;
			RECT	100.145 52.884 100.177 52.948 ;
			RECT	100.313 52.884 100.345 52.948 ;
			RECT	100.481 52.884 100.513 52.948 ;
			RECT	100.649 52.884 100.681 52.948 ;
			RECT	100.817 52.884 100.849 52.948 ;
			RECT	100.985 52.884 101.017 52.948 ;
			RECT	101.153 52.884 101.185 52.948 ;
			RECT	101.321 52.884 101.353 52.948 ;
			RECT	101.489 52.884 101.521 52.948 ;
			RECT	101.657 52.884 101.689 52.948 ;
			RECT	101.825 52.884 101.857 52.948 ;
			RECT	101.993 52.884 102.025 52.948 ;
			RECT	102.123 52.9 102.155 52.932 ;
			RECT	102.245 52.895 102.277 52.927 ;
			RECT	102.375 52.884 102.407 52.948 ;
			RECT	103.795 52.884 103.827 52.948 ;
			RECT	103.925 52.895 103.957 52.927 ;
			RECT	104.047 52.9 104.079 52.932 ;
			RECT	104.177 52.884 104.209 52.948 ;
			RECT	104.345 52.884 104.377 52.948 ;
			RECT	104.513 52.884 104.545 52.948 ;
			RECT	104.681 52.884 104.713 52.948 ;
			RECT	104.849 52.884 104.881 52.948 ;
			RECT	105.017 52.884 105.049 52.948 ;
			RECT	105.185 52.884 105.217 52.948 ;
			RECT	105.353 52.884 105.385 52.948 ;
			RECT	105.521 52.884 105.553 52.948 ;
			RECT	105.689 52.884 105.721 52.948 ;
			RECT	105.857 52.884 105.889 52.948 ;
			RECT	106.025 52.884 106.057 52.948 ;
			RECT	106.193 52.884 106.225 52.948 ;
			RECT	106.361 52.884 106.393 52.948 ;
			RECT	106.529 52.884 106.561 52.948 ;
			RECT	106.697 52.884 106.729 52.948 ;
			RECT	106.865 52.884 106.897 52.948 ;
			RECT	107.033 52.884 107.065 52.948 ;
			RECT	107.201 52.884 107.233 52.948 ;
			RECT	107.369 52.884 107.401 52.948 ;
			RECT	107.537 52.884 107.569 52.948 ;
			RECT	107.705 52.884 107.737 52.948 ;
			RECT	107.873 52.884 107.905 52.948 ;
			RECT	108.041 52.884 108.073 52.948 ;
			RECT	108.209 52.884 108.241 52.948 ;
			RECT	108.377 52.884 108.409 52.948 ;
			RECT	108.545 52.884 108.577 52.948 ;
			RECT	108.713 52.884 108.745 52.948 ;
			RECT	108.881 52.884 108.913 52.948 ;
			RECT	109.049 52.884 109.081 52.948 ;
			RECT	109.217 52.884 109.249 52.948 ;
			RECT	109.385 52.884 109.417 52.948 ;
			RECT	109.553 52.884 109.585 52.948 ;
			RECT	109.721 52.884 109.753 52.948 ;
			RECT	109.889 52.884 109.921 52.948 ;
			RECT	110.057 52.884 110.089 52.948 ;
			RECT	110.225 52.884 110.257 52.948 ;
			RECT	110.393 52.884 110.425 52.948 ;
			RECT	110.561 52.884 110.593 52.948 ;
			RECT	110.729 52.884 110.761 52.948 ;
			RECT	110.897 52.884 110.929 52.948 ;
			RECT	111.065 52.884 111.097 52.948 ;
			RECT	111.233 52.884 111.265 52.948 ;
			RECT	111.401 52.884 111.433 52.948 ;
			RECT	111.569 52.884 111.601 52.948 ;
			RECT	111.737 52.884 111.769 52.948 ;
			RECT	111.905 52.884 111.937 52.948 ;
			RECT	112.073 52.884 112.105 52.948 ;
			RECT	112.241 52.884 112.273 52.948 ;
			RECT	112.409 52.884 112.441 52.948 ;
			RECT	112.577 52.884 112.609 52.948 ;
			RECT	112.745 52.884 112.777 52.948 ;
			RECT	112.913 52.884 112.945 52.948 ;
			RECT	113.081 52.884 113.113 52.948 ;
			RECT	113.249 52.884 113.281 52.948 ;
			RECT	113.417 52.884 113.449 52.948 ;
			RECT	113.585 52.884 113.617 52.948 ;
			RECT	113.753 52.884 113.785 52.948 ;
			RECT	113.921 52.884 113.953 52.948 ;
			RECT	114.089 52.884 114.121 52.948 ;
			RECT	114.257 52.884 114.289 52.948 ;
			RECT	114.425 52.884 114.457 52.948 ;
			RECT	114.593 52.884 114.625 52.948 ;
			RECT	114.761 52.884 114.793 52.948 ;
			RECT	114.929 52.884 114.961 52.948 ;
			RECT	115.097 52.884 115.129 52.948 ;
			RECT	115.265 52.884 115.297 52.948 ;
			RECT	115.433 52.884 115.465 52.948 ;
			RECT	115.601 52.884 115.633 52.948 ;
			RECT	115.769 52.884 115.801 52.948 ;
			RECT	115.937 52.884 115.969 52.948 ;
			RECT	116.105 52.884 116.137 52.948 ;
			RECT	116.273 52.884 116.305 52.948 ;
			RECT	116.441 52.884 116.473 52.948 ;
			RECT	116.609 52.884 116.641 52.948 ;
			RECT	116.777 52.884 116.809 52.948 ;
			RECT	116.945 52.884 116.977 52.948 ;
			RECT	117.113 52.884 117.145 52.948 ;
			RECT	117.281 52.884 117.313 52.948 ;
			RECT	117.449 52.884 117.481 52.948 ;
			RECT	117.617 52.884 117.649 52.948 ;
			RECT	117.785 52.884 117.817 52.948 ;
			RECT	117.953 52.884 117.985 52.948 ;
			RECT	118.121 52.884 118.153 52.948 ;
			RECT	118.289 52.884 118.321 52.948 ;
			RECT	118.457 52.884 118.489 52.948 ;
			RECT	118.625 52.884 118.657 52.948 ;
			RECT	118.793 52.884 118.825 52.948 ;
			RECT	118.961 52.884 118.993 52.948 ;
			RECT	119.129 52.884 119.161 52.948 ;
			RECT	119.297 52.884 119.329 52.948 ;
			RECT	119.465 52.884 119.497 52.948 ;
			RECT	119.633 52.884 119.665 52.948 ;
			RECT	119.801 52.884 119.833 52.948 ;
			RECT	119.969 52.884 120.001 52.948 ;
			RECT	120.137 52.884 120.169 52.948 ;
			RECT	120.305 52.884 120.337 52.948 ;
			RECT	120.473 52.884 120.505 52.948 ;
			RECT	120.641 52.884 120.673 52.948 ;
			RECT	120.809 52.884 120.841 52.948 ;
			RECT	120.977 52.884 121.009 52.948 ;
			RECT	121.145 52.884 121.177 52.948 ;
			RECT	121.313 52.884 121.345 52.948 ;
			RECT	121.481 52.884 121.513 52.948 ;
			RECT	121.649 52.884 121.681 52.948 ;
			RECT	121.817 52.884 121.849 52.948 ;
			RECT	121.985 52.884 122.017 52.948 ;
			RECT	122.153 52.884 122.185 52.948 ;
			RECT	122.321 52.884 122.353 52.948 ;
			RECT	122.489 52.884 122.521 52.948 ;
			RECT	122.657 52.884 122.689 52.948 ;
			RECT	122.825 52.884 122.857 52.948 ;
			RECT	122.993 52.884 123.025 52.948 ;
			RECT	123.161 52.884 123.193 52.948 ;
			RECT	123.329 52.884 123.361 52.948 ;
			RECT	123.497 52.884 123.529 52.948 ;
			RECT	123.665 52.884 123.697 52.948 ;
			RECT	123.833 52.884 123.865 52.948 ;
			RECT	124.001 52.884 124.033 52.948 ;
			RECT	124.169 52.884 124.201 52.948 ;
			RECT	124.337 52.884 124.369 52.948 ;
			RECT	124.505 52.884 124.537 52.948 ;
			RECT	124.673 52.884 124.705 52.948 ;
			RECT	124.841 52.884 124.873 52.948 ;
			RECT	125.009 52.884 125.041 52.948 ;
			RECT	125.177 52.884 125.209 52.948 ;
			RECT	125.345 52.884 125.377 52.948 ;
			RECT	125.513 52.884 125.545 52.948 ;
			RECT	125.681 52.884 125.713 52.948 ;
			RECT	125.849 52.884 125.881 52.948 ;
			RECT	126.017 52.884 126.049 52.948 ;
			RECT	126.185 52.884 126.217 52.948 ;
			RECT	126.353 52.884 126.385 52.948 ;
			RECT	126.521 52.884 126.553 52.948 ;
			RECT	126.689 52.884 126.721 52.948 ;
			RECT	126.857 52.884 126.889 52.948 ;
			RECT	127.025 52.884 127.057 52.948 ;
			RECT	127.193 52.884 127.225 52.948 ;
			RECT	127.361 52.884 127.393 52.948 ;
			RECT	127.529 52.884 127.561 52.948 ;
			RECT	127.697 52.884 127.729 52.948 ;
			RECT	127.865 52.884 127.897 52.948 ;
			RECT	128.033 52.884 128.065 52.948 ;
			RECT	128.201 52.884 128.233 52.948 ;
			RECT	128.369 52.884 128.401 52.948 ;
			RECT	128.537 52.884 128.569 52.948 ;
			RECT	128.705 52.884 128.737 52.948 ;
			RECT	128.873 52.884 128.905 52.948 ;
			RECT	129.041 52.884 129.073 52.948 ;
			RECT	129.209 52.884 129.241 52.948 ;
			RECT	129.377 52.884 129.409 52.948 ;
			RECT	129.545 52.884 129.577 52.948 ;
			RECT	129.713 52.884 129.745 52.948 ;
			RECT	129.881 52.884 129.913 52.948 ;
			RECT	130.049 52.884 130.081 52.948 ;
			RECT	130.217 52.884 130.249 52.948 ;
			RECT	130.385 52.884 130.417 52.948 ;
			RECT	130.553 52.884 130.585 52.948 ;
			RECT	130.721 52.884 130.753 52.948 ;
			RECT	130.889 52.884 130.921 52.948 ;
			RECT	131.057 52.884 131.089 52.948 ;
			RECT	131.225 52.884 131.257 52.948 ;
			RECT	131.393 52.884 131.425 52.948 ;
			RECT	131.561 52.884 131.593 52.948 ;
			RECT	131.729 52.884 131.761 52.948 ;
			RECT	131.897 52.884 131.929 52.948 ;
			RECT	132.065 52.884 132.097 52.948 ;
			RECT	132.233 52.884 132.265 52.948 ;
			RECT	132.401 52.884 132.433 52.948 ;
			RECT	132.569 52.884 132.601 52.948 ;
			RECT	132.737 52.884 132.769 52.948 ;
			RECT	132.905 52.884 132.937 52.948 ;
			RECT	133.073 52.884 133.105 52.948 ;
			RECT	133.241 52.884 133.273 52.948 ;
			RECT	133.409 52.884 133.441 52.948 ;
			RECT	133.577 52.884 133.609 52.948 ;
			RECT	133.745 52.884 133.777 52.948 ;
			RECT	133.913 52.884 133.945 52.948 ;
			RECT	134.081 52.884 134.113 52.948 ;
			RECT	134.249 52.884 134.281 52.948 ;
			RECT	134.417 52.884 134.449 52.948 ;
			RECT	134.585 52.884 134.617 52.948 ;
			RECT	134.753 52.884 134.785 52.948 ;
			RECT	134.921 52.884 134.953 52.948 ;
			RECT	135.089 52.884 135.121 52.948 ;
			RECT	135.257 52.884 135.289 52.948 ;
			RECT	135.425 52.884 135.457 52.948 ;
			RECT	135.593 52.884 135.625 52.948 ;
			RECT	135.761 52.884 135.793 52.948 ;
			RECT	135.929 52.884 135.961 52.948 ;
			RECT	136.097 52.884 136.129 52.948 ;
			RECT	136.265 52.884 136.297 52.948 ;
			RECT	136.433 52.884 136.465 52.948 ;
			RECT	136.601 52.884 136.633 52.948 ;
			RECT	136.769 52.884 136.801 52.948 ;
			RECT	136.937 52.884 136.969 52.948 ;
			RECT	137.105 52.884 137.137 52.948 ;
			RECT	137.273 52.884 137.305 52.948 ;
			RECT	137.441 52.884 137.473 52.948 ;
			RECT	137.609 52.884 137.641 52.948 ;
			RECT	137.777 52.884 137.809 52.948 ;
			RECT	137.945 52.884 137.977 52.948 ;
			RECT	138.113 52.884 138.145 52.948 ;
			RECT	138.281 52.884 138.313 52.948 ;
			RECT	138.449 52.884 138.481 52.948 ;
			RECT	138.617 52.884 138.649 52.948 ;
			RECT	138.785 52.884 138.817 52.948 ;
			RECT	138.953 52.884 138.985 52.948 ;
			RECT	139.121 52.884 139.153 52.948 ;
			RECT	139.289 52.884 139.321 52.948 ;
			RECT	139.457 52.884 139.489 52.948 ;
			RECT	139.625 52.884 139.657 52.948 ;
			RECT	139.793 52.884 139.825 52.948 ;
			RECT	139.961 52.884 139.993 52.948 ;
			RECT	140.129 52.884 140.161 52.948 ;
			RECT	140.297 52.884 140.329 52.948 ;
			RECT	140.465 52.884 140.497 52.948 ;
			RECT	140.633 52.884 140.665 52.948 ;
			RECT	140.801 52.884 140.833 52.948 ;
			RECT	140.969 52.884 141.001 52.948 ;
			RECT	141.137 52.884 141.169 52.948 ;
			RECT	141.305 52.884 141.337 52.948 ;
			RECT	141.473 52.884 141.505 52.948 ;
			RECT	141.641 52.884 141.673 52.948 ;
			RECT	141.809 52.884 141.841 52.948 ;
			RECT	141.977 52.884 142.009 52.948 ;
			RECT	142.145 52.884 142.177 52.948 ;
			RECT	142.313 52.884 142.345 52.948 ;
			RECT	142.481 52.884 142.513 52.948 ;
			RECT	142.649 52.884 142.681 52.948 ;
			RECT	142.817 52.884 142.849 52.948 ;
			RECT	142.985 52.884 143.017 52.948 ;
			RECT	143.153 52.884 143.185 52.948 ;
			RECT	143.321 52.884 143.353 52.948 ;
			RECT	143.489 52.884 143.521 52.948 ;
			RECT	143.657 52.884 143.689 52.948 ;
			RECT	143.825 52.884 143.857 52.948 ;
			RECT	143.993 52.884 144.025 52.948 ;
			RECT	144.161 52.884 144.193 52.948 ;
			RECT	144.329 52.884 144.361 52.948 ;
			RECT	144.497 52.884 144.529 52.948 ;
			RECT	144.665 52.884 144.697 52.948 ;
			RECT	144.833 52.884 144.865 52.948 ;
			RECT	145.001 52.884 145.033 52.948 ;
			RECT	145.169 52.884 145.201 52.948 ;
			RECT	145.337 52.884 145.369 52.948 ;
			RECT	145.505 52.884 145.537 52.948 ;
			RECT	145.673 52.884 145.705 52.948 ;
			RECT	145.841 52.884 145.873 52.948 ;
			RECT	146.009 52.884 146.041 52.948 ;
			RECT	146.177 52.884 146.209 52.948 ;
			RECT	146.345 52.884 146.377 52.948 ;
			RECT	146.513 52.884 146.545 52.948 ;
			RECT	146.681 52.884 146.713 52.948 ;
			RECT	146.849 52.884 146.881 52.948 ;
			RECT	147.017 52.884 147.049 52.948 ;
			RECT	147.185 52.884 147.217 52.948 ;
			RECT	147.316 52.9 147.348 52.932 ;
			RECT	147.437 52.9 147.469 52.932 ;
			RECT	147.567 52.884 147.599 52.948 ;
			RECT	149.879 52.884 149.911 52.948 ;
			RECT	151.13 52.884 151.194 52.948 ;
			RECT	151.81 52.884 151.842 52.948 ;
			RECT	152.249 52.884 152.281 52.948 ;
			RECT	153.56 52.884 153.624 52.948 ;
			RECT	156.601 52.884 156.633 52.948 ;
			RECT	156.731 52.9 156.763 52.932 ;
			RECT	156.852 52.9 156.884 52.932 ;
			RECT	156.983 52.884 157.015 52.948 ;
			RECT	157.151 52.884 157.183 52.948 ;
			RECT	157.319 52.884 157.351 52.948 ;
			RECT	157.487 52.884 157.519 52.948 ;
			RECT	157.655 52.884 157.687 52.948 ;
			RECT	157.823 52.884 157.855 52.948 ;
			RECT	157.991 52.884 158.023 52.948 ;
			RECT	158.159 52.884 158.191 52.948 ;
			RECT	158.327 52.884 158.359 52.948 ;
			RECT	158.495 52.884 158.527 52.948 ;
			RECT	158.663 52.884 158.695 52.948 ;
			RECT	158.831 52.884 158.863 52.948 ;
			RECT	158.999 52.884 159.031 52.948 ;
			RECT	159.167 52.884 159.199 52.948 ;
			RECT	159.335 52.884 159.367 52.948 ;
			RECT	159.503 52.884 159.535 52.948 ;
			RECT	159.671 52.884 159.703 52.948 ;
			RECT	159.839 52.884 159.871 52.948 ;
			RECT	160.007 52.884 160.039 52.948 ;
			RECT	160.175 52.884 160.207 52.948 ;
			RECT	160.343 52.884 160.375 52.948 ;
			RECT	160.511 52.884 160.543 52.948 ;
			RECT	160.679 52.884 160.711 52.948 ;
			RECT	160.847 52.884 160.879 52.948 ;
			RECT	161.015 52.884 161.047 52.948 ;
			RECT	161.183 52.884 161.215 52.948 ;
			RECT	161.351 52.884 161.383 52.948 ;
			RECT	161.519 52.884 161.551 52.948 ;
			RECT	161.687 52.884 161.719 52.948 ;
			RECT	161.855 52.884 161.887 52.948 ;
			RECT	162.023 52.884 162.055 52.948 ;
			RECT	162.191 52.884 162.223 52.948 ;
			RECT	162.359 52.884 162.391 52.948 ;
			RECT	162.527 52.884 162.559 52.948 ;
			RECT	162.695 52.884 162.727 52.948 ;
			RECT	162.863 52.884 162.895 52.948 ;
			RECT	163.031 52.884 163.063 52.948 ;
			RECT	163.199 52.884 163.231 52.948 ;
			RECT	163.367 52.884 163.399 52.948 ;
			RECT	163.535 52.884 163.567 52.948 ;
			RECT	163.703 52.884 163.735 52.948 ;
			RECT	163.871 52.884 163.903 52.948 ;
			RECT	164.039 52.884 164.071 52.948 ;
			RECT	164.207 52.884 164.239 52.948 ;
			RECT	164.375 52.884 164.407 52.948 ;
			RECT	164.543 52.884 164.575 52.948 ;
			RECT	164.711 52.884 164.743 52.948 ;
			RECT	164.879 52.884 164.911 52.948 ;
			RECT	165.047 52.884 165.079 52.948 ;
			RECT	165.215 52.884 165.247 52.948 ;
			RECT	165.383 52.884 165.415 52.948 ;
			RECT	165.551 52.884 165.583 52.948 ;
			RECT	165.719 52.884 165.751 52.948 ;
			RECT	165.887 52.884 165.919 52.948 ;
			RECT	166.055 52.884 166.087 52.948 ;
			RECT	166.223 52.884 166.255 52.948 ;
			RECT	166.391 52.884 166.423 52.948 ;
			RECT	166.559 52.884 166.591 52.948 ;
			RECT	166.727 52.884 166.759 52.948 ;
			RECT	166.895 52.884 166.927 52.948 ;
			RECT	167.063 52.884 167.095 52.948 ;
			RECT	167.231 52.884 167.263 52.948 ;
			RECT	167.399 52.884 167.431 52.948 ;
			RECT	167.567 52.884 167.599 52.948 ;
			RECT	167.735 52.884 167.767 52.948 ;
			RECT	167.903 52.884 167.935 52.948 ;
			RECT	168.071 52.884 168.103 52.948 ;
			RECT	168.239 52.884 168.271 52.948 ;
			RECT	168.407 52.884 168.439 52.948 ;
			RECT	168.575 52.884 168.607 52.948 ;
			RECT	168.743 52.884 168.775 52.948 ;
			RECT	168.911 52.884 168.943 52.948 ;
			RECT	169.079 52.884 169.111 52.948 ;
			RECT	169.247 52.884 169.279 52.948 ;
			RECT	169.415 52.884 169.447 52.948 ;
			RECT	169.583 52.884 169.615 52.948 ;
			RECT	169.751 52.884 169.783 52.948 ;
			RECT	169.919 52.884 169.951 52.948 ;
			RECT	170.087 52.884 170.119 52.948 ;
			RECT	170.255 52.884 170.287 52.948 ;
			RECT	170.423 52.884 170.455 52.948 ;
			RECT	170.591 52.884 170.623 52.948 ;
			RECT	170.759 52.884 170.791 52.948 ;
			RECT	170.927 52.884 170.959 52.948 ;
			RECT	171.095 52.884 171.127 52.948 ;
			RECT	171.263 52.884 171.295 52.948 ;
			RECT	171.431 52.884 171.463 52.948 ;
			RECT	171.599 52.884 171.631 52.948 ;
			RECT	171.767 52.884 171.799 52.948 ;
			RECT	171.935 52.884 171.967 52.948 ;
			RECT	172.103 52.884 172.135 52.948 ;
			RECT	172.271 52.884 172.303 52.948 ;
			RECT	172.439 52.884 172.471 52.948 ;
			RECT	172.607 52.884 172.639 52.948 ;
			RECT	172.775 52.884 172.807 52.948 ;
			RECT	172.943 52.884 172.975 52.948 ;
			RECT	173.111 52.884 173.143 52.948 ;
			RECT	173.279 52.884 173.311 52.948 ;
			RECT	173.447 52.884 173.479 52.948 ;
			RECT	173.615 52.884 173.647 52.948 ;
			RECT	173.783 52.884 173.815 52.948 ;
			RECT	173.951 52.884 173.983 52.948 ;
			RECT	174.119 52.884 174.151 52.948 ;
			RECT	174.287 52.884 174.319 52.948 ;
			RECT	174.455 52.884 174.487 52.948 ;
			RECT	174.623 52.884 174.655 52.948 ;
			RECT	174.791 52.884 174.823 52.948 ;
			RECT	174.959 52.884 174.991 52.948 ;
			RECT	175.127 52.884 175.159 52.948 ;
			RECT	175.295 52.884 175.327 52.948 ;
			RECT	175.463 52.884 175.495 52.948 ;
			RECT	175.631 52.884 175.663 52.948 ;
			RECT	175.799 52.884 175.831 52.948 ;
			RECT	175.967 52.884 175.999 52.948 ;
			RECT	176.135 52.884 176.167 52.948 ;
			RECT	176.303 52.884 176.335 52.948 ;
			RECT	176.471 52.884 176.503 52.948 ;
			RECT	176.639 52.884 176.671 52.948 ;
			RECT	176.807 52.884 176.839 52.948 ;
			RECT	176.975 52.884 177.007 52.948 ;
			RECT	177.143 52.884 177.175 52.948 ;
			RECT	177.311 52.884 177.343 52.948 ;
			RECT	177.479 52.884 177.511 52.948 ;
			RECT	177.647 52.884 177.679 52.948 ;
			RECT	177.815 52.884 177.847 52.948 ;
			RECT	177.983 52.884 178.015 52.948 ;
			RECT	178.151 52.884 178.183 52.948 ;
			RECT	178.319 52.884 178.351 52.948 ;
			RECT	178.487 52.884 178.519 52.948 ;
			RECT	178.655 52.884 178.687 52.948 ;
			RECT	178.823 52.884 178.855 52.948 ;
			RECT	178.991 52.884 179.023 52.948 ;
			RECT	179.159 52.884 179.191 52.948 ;
			RECT	179.327 52.884 179.359 52.948 ;
			RECT	179.495 52.884 179.527 52.948 ;
			RECT	179.663 52.884 179.695 52.948 ;
			RECT	179.831 52.884 179.863 52.948 ;
			RECT	179.999 52.884 180.031 52.948 ;
			RECT	180.167 52.884 180.199 52.948 ;
			RECT	180.335 52.884 180.367 52.948 ;
			RECT	180.503 52.884 180.535 52.948 ;
			RECT	180.671 52.884 180.703 52.948 ;
			RECT	180.839 52.884 180.871 52.948 ;
			RECT	181.007 52.884 181.039 52.948 ;
			RECT	181.175 52.884 181.207 52.948 ;
			RECT	181.343 52.884 181.375 52.948 ;
			RECT	181.511 52.884 181.543 52.948 ;
			RECT	181.679 52.884 181.711 52.948 ;
			RECT	181.847 52.884 181.879 52.948 ;
			RECT	182.015 52.884 182.047 52.948 ;
			RECT	182.183 52.884 182.215 52.948 ;
			RECT	182.351 52.884 182.383 52.948 ;
			RECT	182.519 52.884 182.551 52.948 ;
			RECT	182.687 52.884 182.719 52.948 ;
			RECT	182.855 52.884 182.887 52.948 ;
			RECT	183.023 52.884 183.055 52.948 ;
			RECT	183.191 52.884 183.223 52.948 ;
			RECT	183.359 52.884 183.391 52.948 ;
			RECT	183.527 52.884 183.559 52.948 ;
			RECT	183.695 52.884 183.727 52.948 ;
			RECT	183.863 52.884 183.895 52.948 ;
			RECT	184.031 52.884 184.063 52.948 ;
			RECT	184.199 52.884 184.231 52.948 ;
			RECT	184.367 52.884 184.399 52.948 ;
			RECT	184.535 52.884 184.567 52.948 ;
			RECT	184.703 52.884 184.735 52.948 ;
			RECT	184.871 52.884 184.903 52.948 ;
			RECT	185.039 52.884 185.071 52.948 ;
			RECT	185.207 52.884 185.239 52.948 ;
			RECT	185.375 52.884 185.407 52.948 ;
			RECT	185.543 52.884 185.575 52.948 ;
			RECT	185.711 52.884 185.743 52.948 ;
			RECT	185.879 52.884 185.911 52.948 ;
			RECT	186.047 52.884 186.079 52.948 ;
			RECT	186.215 52.884 186.247 52.948 ;
			RECT	186.383 52.884 186.415 52.948 ;
			RECT	186.551 52.884 186.583 52.948 ;
			RECT	186.719 52.884 186.751 52.948 ;
			RECT	186.887 52.884 186.919 52.948 ;
			RECT	187.055 52.884 187.087 52.948 ;
			RECT	187.223 52.884 187.255 52.948 ;
			RECT	187.391 52.884 187.423 52.948 ;
			RECT	187.559 52.884 187.591 52.948 ;
			RECT	187.727 52.884 187.759 52.948 ;
			RECT	187.895 52.884 187.927 52.948 ;
			RECT	188.063 52.884 188.095 52.948 ;
			RECT	188.231 52.884 188.263 52.948 ;
			RECT	188.399 52.884 188.431 52.948 ;
			RECT	188.567 52.884 188.599 52.948 ;
			RECT	188.735 52.884 188.767 52.948 ;
			RECT	188.903 52.884 188.935 52.948 ;
			RECT	189.071 52.884 189.103 52.948 ;
			RECT	189.239 52.884 189.271 52.948 ;
			RECT	189.407 52.884 189.439 52.948 ;
			RECT	189.575 52.884 189.607 52.948 ;
			RECT	189.743 52.884 189.775 52.948 ;
			RECT	189.911 52.884 189.943 52.948 ;
			RECT	190.079 52.884 190.111 52.948 ;
			RECT	190.247 52.884 190.279 52.948 ;
			RECT	190.415 52.884 190.447 52.948 ;
			RECT	190.583 52.884 190.615 52.948 ;
			RECT	190.751 52.884 190.783 52.948 ;
			RECT	190.919 52.884 190.951 52.948 ;
			RECT	191.087 52.884 191.119 52.948 ;
			RECT	191.255 52.884 191.287 52.948 ;
			RECT	191.423 52.884 191.455 52.948 ;
			RECT	191.591 52.884 191.623 52.948 ;
			RECT	191.759 52.884 191.791 52.948 ;
			RECT	191.927 52.884 191.959 52.948 ;
			RECT	192.095 52.884 192.127 52.948 ;
			RECT	192.263 52.884 192.295 52.948 ;
			RECT	192.431 52.884 192.463 52.948 ;
			RECT	192.599 52.884 192.631 52.948 ;
			RECT	192.767 52.884 192.799 52.948 ;
			RECT	192.935 52.884 192.967 52.948 ;
			RECT	193.103 52.884 193.135 52.948 ;
			RECT	193.271 52.884 193.303 52.948 ;
			RECT	193.439 52.884 193.471 52.948 ;
			RECT	193.607 52.884 193.639 52.948 ;
			RECT	193.775 52.884 193.807 52.948 ;
			RECT	193.943 52.884 193.975 52.948 ;
			RECT	194.111 52.884 194.143 52.948 ;
			RECT	194.279 52.884 194.311 52.948 ;
			RECT	194.447 52.884 194.479 52.948 ;
			RECT	194.615 52.884 194.647 52.948 ;
			RECT	194.783 52.884 194.815 52.948 ;
			RECT	194.951 52.884 194.983 52.948 ;
			RECT	195.119 52.884 195.151 52.948 ;
			RECT	195.287 52.884 195.319 52.948 ;
			RECT	195.455 52.884 195.487 52.948 ;
			RECT	195.623 52.884 195.655 52.948 ;
			RECT	195.791 52.884 195.823 52.948 ;
			RECT	195.959 52.884 195.991 52.948 ;
			RECT	196.127 52.884 196.159 52.948 ;
			RECT	196.295 52.884 196.327 52.948 ;
			RECT	196.463 52.884 196.495 52.948 ;
			RECT	196.631 52.884 196.663 52.948 ;
			RECT	196.799 52.884 196.831 52.948 ;
			RECT	196.967 52.884 196.999 52.948 ;
			RECT	197.135 52.884 197.167 52.948 ;
			RECT	197.303 52.884 197.335 52.948 ;
			RECT	197.471 52.884 197.503 52.948 ;
			RECT	197.639 52.884 197.671 52.948 ;
			RECT	197.807 52.884 197.839 52.948 ;
			RECT	197.975 52.884 198.007 52.948 ;
			RECT	198.143 52.884 198.175 52.948 ;
			RECT	198.311 52.884 198.343 52.948 ;
			RECT	198.479 52.884 198.511 52.948 ;
			RECT	198.647 52.884 198.679 52.948 ;
			RECT	198.815 52.884 198.847 52.948 ;
			RECT	198.983 52.884 199.015 52.948 ;
			RECT	199.151 52.884 199.183 52.948 ;
			RECT	199.319 52.884 199.351 52.948 ;
			RECT	199.487 52.884 199.519 52.948 ;
			RECT	199.655 52.884 199.687 52.948 ;
			RECT	199.823 52.884 199.855 52.948 ;
			RECT	199.991 52.884 200.023 52.948 ;
			RECT	200.121 52.9 200.153 52.932 ;
			RECT	200.243 52.895 200.275 52.927 ;
			RECT	200.373 52.884 200.405 52.948 ;
			RECT	200.9 52.884 200.932 52.948 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 50.936 201.665 51.056 ;
			LAYER	J3 ;
			RECT	0.755 50.964 0.787 51.028 ;
			RECT	1.645 50.964 1.709 51.028 ;
			RECT	2.323 50.964 2.387 51.028 ;
			RECT	3.438 50.964 3.47 51.028 ;
			RECT	3.585 50.964 3.617 51.028 ;
			RECT	4.195 50.964 4.227 51.028 ;
			RECT	4.72 50.964 4.752 51.028 ;
			RECT	4.944 50.964 5.008 51.028 ;
			RECT	5.267 50.964 5.299 51.028 ;
			RECT	5.797 50.964 5.829 51.028 ;
			RECT	5.927 50.975 5.959 51.007 ;
			RECT	6.049 50.98 6.081 51.012 ;
			RECT	6.179 50.964 6.211 51.028 ;
			RECT	6.347 50.964 6.379 51.028 ;
			RECT	6.515 50.964 6.547 51.028 ;
			RECT	6.683 50.964 6.715 51.028 ;
			RECT	6.851 50.964 6.883 51.028 ;
			RECT	7.019 50.964 7.051 51.028 ;
			RECT	7.187 50.964 7.219 51.028 ;
			RECT	7.355 50.964 7.387 51.028 ;
			RECT	7.523 50.964 7.555 51.028 ;
			RECT	7.691 50.964 7.723 51.028 ;
			RECT	7.859 50.964 7.891 51.028 ;
			RECT	8.027 50.964 8.059 51.028 ;
			RECT	8.195 50.964 8.227 51.028 ;
			RECT	8.363 50.964 8.395 51.028 ;
			RECT	8.531 50.964 8.563 51.028 ;
			RECT	8.699 50.964 8.731 51.028 ;
			RECT	8.867 50.964 8.899 51.028 ;
			RECT	9.035 50.964 9.067 51.028 ;
			RECT	9.203 50.964 9.235 51.028 ;
			RECT	9.371 50.964 9.403 51.028 ;
			RECT	9.539 50.964 9.571 51.028 ;
			RECT	9.707 50.964 9.739 51.028 ;
			RECT	9.875 50.964 9.907 51.028 ;
			RECT	10.043 50.964 10.075 51.028 ;
			RECT	10.211 50.964 10.243 51.028 ;
			RECT	10.379 50.964 10.411 51.028 ;
			RECT	10.547 50.964 10.579 51.028 ;
			RECT	10.715 50.964 10.747 51.028 ;
			RECT	10.883 50.964 10.915 51.028 ;
			RECT	11.051 50.964 11.083 51.028 ;
			RECT	11.219 50.964 11.251 51.028 ;
			RECT	11.387 50.964 11.419 51.028 ;
			RECT	11.555 50.964 11.587 51.028 ;
			RECT	11.723 50.964 11.755 51.028 ;
			RECT	11.891 50.964 11.923 51.028 ;
			RECT	12.059 50.964 12.091 51.028 ;
			RECT	12.227 50.964 12.259 51.028 ;
			RECT	12.395 50.964 12.427 51.028 ;
			RECT	12.563 50.964 12.595 51.028 ;
			RECT	12.731 50.964 12.763 51.028 ;
			RECT	12.899 50.964 12.931 51.028 ;
			RECT	13.067 50.964 13.099 51.028 ;
			RECT	13.235 50.964 13.267 51.028 ;
			RECT	13.403 50.964 13.435 51.028 ;
			RECT	13.571 50.964 13.603 51.028 ;
			RECT	13.739 50.964 13.771 51.028 ;
			RECT	13.907 50.964 13.939 51.028 ;
			RECT	14.075 50.964 14.107 51.028 ;
			RECT	14.243 50.964 14.275 51.028 ;
			RECT	14.411 50.964 14.443 51.028 ;
			RECT	14.579 50.964 14.611 51.028 ;
			RECT	14.747 50.964 14.779 51.028 ;
			RECT	14.915 50.964 14.947 51.028 ;
			RECT	15.083 50.964 15.115 51.028 ;
			RECT	15.251 50.964 15.283 51.028 ;
			RECT	15.419 50.964 15.451 51.028 ;
			RECT	15.587 50.964 15.619 51.028 ;
			RECT	15.755 50.964 15.787 51.028 ;
			RECT	15.923 50.964 15.955 51.028 ;
			RECT	16.091 50.964 16.123 51.028 ;
			RECT	16.259 50.964 16.291 51.028 ;
			RECT	16.427 50.964 16.459 51.028 ;
			RECT	16.595 50.964 16.627 51.028 ;
			RECT	16.763 50.964 16.795 51.028 ;
			RECT	16.931 50.964 16.963 51.028 ;
			RECT	17.099 50.964 17.131 51.028 ;
			RECT	17.267 50.964 17.299 51.028 ;
			RECT	17.435 50.964 17.467 51.028 ;
			RECT	17.603 50.964 17.635 51.028 ;
			RECT	17.771 50.964 17.803 51.028 ;
			RECT	17.939 50.964 17.971 51.028 ;
			RECT	18.107 50.964 18.139 51.028 ;
			RECT	18.275 50.964 18.307 51.028 ;
			RECT	18.443 50.964 18.475 51.028 ;
			RECT	18.611 50.964 18.643 51.028 ;
			RECT	18.779 50.964 18.811 51.028 ;
			RECT	18.947 50.964 18.979 51.028 ;
			RECT	19.115 50.964 19.147 51.028 ;
			RECT	19.283 50.964 19.315 51.028 ;
			RECT	19.451 50.964 19.483 51.028 ;
			RECT	19.619 50.964 19.651 51.028 ;
			RECT	19.787 50.964 19.819 51.028 ;
			RECT	19.955 50.964 19.987 51.028 ;
			RECT	20.123 50.964 20.155 51.028 ;
			RECT	20.291 50.964 20.323 51.028 ;
			RECT	20.459 50.964 20.491 51.028 ;
			RECT	20.627 50.964 20.659 51.028 ;
			RECT	20.795 50.964 20.827 51.028 ;
			RECT	20.963 50.964 20.995 51.028 ;
			RECT	21.131 50.964 21.163 51.028 ;
			RECT	21.299 50.964 21.331 51.028 ;
			RECT	21.467 50.964 21.499 51.028 ;
			RECT	21.635 50.964 21.667 51.028 ;
			RECT	21.803 50.964 21.835 51.028 ;
			RECT	21.971 50.964 22.003 51.028 ;
			RECT	22.139 50.964 22.171 51.028 ;
			RECT	22.307 50.964 22.339 51.028 ;
			RECT	22.475 50.964 22.507 51.028 ;
			RECT	22.643 50.964 22.675 51.028 ;
			RECT	22.811 50.964 22.843 51.028 ;
			RECT	22.979 50.964 23.011 51.028 ;
			RECT	23.147 50.964 23.179 51.028 ;
			RECT	23.315 50.964 23.347 51.028 ;
			RECT	23.483 50.964 23.515 51.028 ;
			RECT	23.651 50.964 23.683 51.028 ;
			RECT	23.819 50.964 23.851 51.028 ;
			RECT	23.987 50.964 24.019 51.028 ;
			RECT	24.155 50.964 24.187 51.028 ;
			RECT	24.323 50.964 24.355 51.028 ;
			RECT	24.491 50.964 24.523 51.028 ;
			RECT	24.659 50.964 24.691 51.028 ;
			RECT	24.827 50.964 24.859 51.028 ;
			RECT	24.995 50.964 25.027 51.028 ;
			RECT	25.163 50.964 25.195 51.028 ;
			RECT	25.331 50.964 25.363 51.028 ;
			RECT	25.499 50.964 25.531 51.028 ;
			RECT	25.667 50.964 25.699 51.028 ;
			RECT	25.835 50.964 25.867 51.028 ;
			RECT	26.003 50.964 26.035 51.028 ;
			RECT	26.171 50.964 26.203 51.028 ;
			RECT	26.339 50.964 26.371 51.028 ;
			RECT	26.507 50.964 26.539 51.028 ;
			RECT	26.675 50.964 26.707 51.028 ;
			RECT	26.843 50.964 26.875 51.028 ;
			RECT	27.011 50.964 27.043 51.028 ;
			RECT	27.179 50.964 27.211 51.028 ;
			RECT	27.347 50.964 27.379 51.028 ;
			RECT	27.515 50.964 27.547 51.028 ;
			RECT	27.683 50.964 27.715 51.028 ;
			RECT	27.851 50.964 27.883 51.028 ;
			RECT	28.019 50.964 28.051 51.028 ;
			RECT	28.187 50.964 28.219 51.028 ;
			RECT	28.355 50.964 28.387 51.028 ;
			RECT	28.523 50.964 28.555 51.028 ;
			RECT	28.691 50.964 28.723 51.028 ;
			RECT	28.859 50.964 28.891 51.028 ;
			RECT	29.027 50.964 29.059 51.028 ;
			RECT	29.195 50.964 29.227 51.028 ;
			RECT	29.363 50.964 29.395 51.028 ;
			RECT	29.531 50.964 29.563 51.028 ;
			RECT	29.699 50.964 29.731 51.028 ;
			RECT	29.867 50.964 29.899 51.028 ;
			RECT	30.035 50.964 30.067 51.028 ;
			RECT	30.203 50.964 30.235 51.028 ;
			RECT	30.371 50.964 30.403 51.028 ;
			RECT	30.539 50.964 30.571 51.028 ;
			RECT	30.707 50.964 30.739 51.028 ;
			RECT	30.875 50.964 30.907 51.028 ;
			RECT	31.043 50.964 31.075 51.028 ;
			RECT	31.211 50.964 31.243 51.028 ;
			RECT	31.379 50.964 31.411 51.028 ;
			RECT	31.547 50.964 31.579 51.028 ;
			RECT	31.715 50.964 31.747 51.028 ;
			RECT	31.883 50.964 31.915 51.028 ;
			RECT	32.051 50.964 32.083 51.028 ;
			RECT	32.219 50.964 32.251 51.028 ;
			RECT	32.387 50.964 32.419 51.028 ;
			RECT	32.555 50.964 32.587 51.028 ;
			RECT	32.723 50.964 32.755 51.028 ;
			RECT	32.891 50.964 32.923 51.028 ;
			RECT	33.059 50.964 33.091 51.028 ;
			RECT	33.227 50.964 33.259 51.028 ;
			RECT	33.395 50.964 33.427 51.028 ;
			RECT	33.563 50.964 33.595 51.028 ;
			RECT	33.731 50.964 33.763 51.028 ;
			RECT	33.899 50.964 33.931 51.028 ;
			RECT	34.067 50.964 34.099 51.028 ;
			RECT	34.235 50.964 34.267 51.028 ;
			RECT	34.403 50.964 34.435 51.028 ;
			RECT	34.571 50.964 34.603 51.028 ;
			RECT	34.739 50.964 34.771 51.028 ;
			RECT	34.907 50.964 34.939 51.028 ;
			RECT	35.075 50.964 35.107 51.028 ;
			RECT	35.243 50.964 35.275 51.028 ;
			RECT	35.411 50.964 35.443 51.028 ;
			RECT	35.579 50.964 35.611 51.028 ;
			RECT	35.747 50.964 35.779 51.028 ;
			RECT	35.915 50.964 35.947 51.028 ;
			RECT	36.083 50.964 36.115 51.028 ;
			RECT	36.251 50.964 36.283 51.028 ;
			RECT	36.419 50.964 36.451 51.028 ;
			RECT	36.587 50.964 36.619 51.028 ;
			RECT	36.755 50.964 36.787 51.028 ;
			RECT	36.923 50.964 36.955 51.028 ;
			RECT	37.091 50.964 37.123 51.028 ;
			RECT	37.259 50.964 37.291 51.028 ;
			RECT	37.427 50.964 37.459 51.028 ;
			RECT	37.595 50.964 37.627 51.028 ;
			RECT	37.763 50.964 37.795 51.028 ;
			RECT	37.931 50.964 37.963 51.028 ;
			RECT	38.099 50.964 38.131 51.028 ;
			RECT	38.267 50.964 38.299 51.028 ;
			RECT	38.435 50.964 38.467 51.028 ;
			RECT	38.603 50.964 38.635 51.028 ;
			RECT	38.771 50.964 38.803 51.028 ;
			RECT	38.939 50.964 38.971 51.028 ;
			RECT	39.107 50.964 39.139 51.028 ;
			RECT	39.275 50.964 39.307 51.028 ;
			RECT	39.443 50.964 39.475 51.028 ;
			RECT	39.611 50.964 39.643 51.028 ;
			RECT	39.779 50.964 39.811 51.028 ;
			RECT	39.947 50.964 39.979 51.028 ;
			RECT	40.115 50.964 40.147 51.028 ;
			RECT	40.283 50.964 40.315 51.028 ;
			RECT	40.451 50.964 40.483 51.028 ;
			RECT	40.619 50.964 40.651 51.028 ;
			RECT	40.787 50.964 40.819 51.028 ;
			RECT	40.955 50.964 40.987 51.028 ;
			RECT	41.123 50.964 41.155 51.028 ;
			RECT	41.291 50.964 41.323 51.028 ;
			RECT	41.459 50.964 41.491 51.028 ;
			RECT	41.627 50.964 41.659 51.028 ;
			RECT	41.795 50.964 41.827 51.028 ;
			RECT	41.963 50.964 41.995 51.028 ;
			RECT	42.131 50.964 42.163 51.028 ;
			RECT	42.299 50.964 42.331 51.028 ;
			RECT	42.467 50.964 42.499 51.028 ;
			RECT	42.635 50.964 42.667 51.028 ;
			RECT	42.803 50.964 42.835 51.028 ;
			RECT	42.971 50.964 43.003 51.028 ;
			RECT	43.139 50.964 43.171 51.028 ;
			RECT	43.307 50.964 43.339 51.028 ;
			RECT	43.475 50.964 43.507 51.028 ;
			RECT	43.643 50.964 43.675 51.028 ;
			RECT	43.811 50.964 43.843 51.028 ;
			RECT	43.979 50.964 44.011 51.028 ;
			RECT	44.147 50.964 44.179 51.028 ;
			RECT	44.315 50.964 44.347 51.028 ;
			RECT	44.483 50.964 44.515 51.028 ;
			RECT	44.651 50.964 44.683 51.028 ;
			RECT	44.819 50.964 44.851 51.028 ;
			RECT	44.987 50.964 45.019 51.028 ;
			RECT	45.155 50.964 45.187 51.028 ;
			RECT	45.323 50.964 45.355 51.028 ;
			RECT	45.491 50.964 45.523 51.028 ;
			RECT	45.659 50.964 45.691 51.028 ;
			RECT	45.827 50.964 45.859 51.028 ;
			RECT	45.995 50.964 46.027 51.028 ;
			RECT	46.163 50.964 46.195 51.028 ;
			RECT	46.331 50.964 46.363 51.028 ;
			RECT	46.499 50.964 46.531 51.028 ;
			RECT	46.667 50.964 46.699 51.028 ;
			RECT	46.835 50.964 46.867 51.028 ;
			RECT	47.003 50.964 47.035 51.028 ;
			RECT	47.171 50.964 47.203 51.028 ;
			RECT	47.339 50.964 47.371 51.028 ;
			RECT	47.507 50.964 47.539 51.028 ;
			RECT	47.675 50.964 47.707 51.028 ;
			RECT	47.843 50.964 47.875 51.028 ;
			RECT	48.011 50.964 48.043 51.028 ;
			RECT	48.179 50.964 48.211 51.028 ;
			RECT	48.347 50.964 48.379 51.028 ;
			RECT	48.515 50.964 48.547 51.028 ;
			RECT	48.683 50.964 48.715 51.028 ;
			RECT	48.851 50.964 48.883 51.028 ;
			RECT	49.019 50.964 49.051 51.028 ;
			RECT	49.187 50.964 49.219 51.028 ;
			RECT	49.318 50.98 49.35 51.012 ;
			RECT	49.439 50.98 49.471 51.012 ;
			RECT	49.569 50.964 49.601 51.028 ;
			RECT	51.881 50.964 51.913 51.028 ;
			RECT	53.132 50.964 53.196 51.028 ;
			RECT	53.812 50.964 53.844 51.028 ;
			RECT	54.251 50.964 54.283 51.028 ;
			RECT	55.562 50.964 55.626 51.028 ;
			RECT	58.603 50.964 58.635 51.028 ;
			RECT	58.733 50.98 58.765 51.012 ;
			RECT	58.854 50.98 58.886 51.012 ;
			RECT	58.985 50.964 59.017 51.028 ;
			RECT	59.153 50.964 59.185 51.028 ;
			RECT	59.321 50.964 59.353 51.028 ;
			RECT	59.489 50.964 59.521 51.028 ;
			RECT	59.657 50.964 59.689 51.028 ;
			RECT	59.825 50.964 59.857 51.028 ;
			RECT	59.993 50.964 60.025 51.028 ;
			RECT	60.161 50.964 60.193 51.028 ;
			RECT	60.329 50.964 60.361 51.028 ;
			RECT	60.497 50.964 60.529 51.028 ;
			RECT	60.665 50.964 60.697 51.028 ;
			RECT	60.833 50.964 60.865 51.028 ;
			RECT	61.001 50.964 61.033 51.028 ;
			RECT	61.169 50.964 61.201 51.028 ;
			RECT	61.337 50.964 61.369 51.028 ;
			RECT	61.505 50.964 61.537 51.028 ;
			RECT	61.673 50.964 61.705 51.028 ;
			RECT	61.841 50.964 61.873 51.028 ;
			RECT	62.009 50.964 62.041 51.028 ;
			RECT	62.177 50.964 62.209 51.028 ;
			RECT	62.345 50.964 62.377 51.028 ;
			RECT	62.513 50.964 62.545 51.028 ;
			RECT	62.681 50.964 62.713 51.028 ;
			RECT	62.849 50.964 62.881 51.028 ;
			RECT	63.017 50.964 63.049 51.028 ;
			RECT	63.185 50.964 63.217 51.028 ;
			RECT	63.353 50.964 63.385 51.028 ;
			RECT	63.521 50.964 63.553 51.028 ;
			RECT	63.689 50.964 63.721 51.028 ;
			RECT	63.857 50.964 63.889 51.028 ;
			RECT	64.025 50.964 64.057 51.028 ;
			RECT	64.193 50.964 64.225 51.028 ;
			RECT	64.361 50.964 64.393 51.028 ;
			RECT	64.529 50.964 64.561 51.028 ;
			RECT	64.697 50.964 64.729 51.028 ;
			RECT	64.865 50.964 64.897 51.028 ;
			RECT	65.033 50.964 65.065 51.028 ;
			RECT	65.201 50.964 65.233 51.028 ;
			RECT	65.369 50.964 65.401 51.028 ;
			RECT	65.537 50.964 65.569 51.028 ;
			RECT	65.705 50.964 65.737 51.028 ;
			RECT	65.873 50.964 65.905 51.028 ;
			RECT	66.041 50.964 66.073 51.028 ;
			RECT	66.209 50.964 66.241 51.028 ;
			RECT	66.377 50.964 66.409 51.028 ;
			RECT	66.545 50.964 66.577 51.028 ;
			RECT	66.713 50.964 66.745 51.028 ;
			RECT	66.881 50.964 66.913 51.028 ;
			RECT	67.049 50.964 67.081 51.028 ;
			RECT	67.217 50.964 67.249 51.028 ;
			RECT	67.385 50.964 67.417 51.028 ;
			RECT	67.553 50.964 67.585 51.028 ;
			RECT	67.721 50.964 67.753 51.028 ;
			RECT	67.889 50.964 67.921 51.028 ;
			RECT	68.057 50.964 68.089 51.028 ;
			RECT	68.225 50.964 68.257 51.028 ;
			RECT	68.393 50.964 68.425 51.028 ;
			RECT	68.561 50.964 68.593 51.028 ;
			RECT	68.729 50.964 68.761 51.028 ;
			RECT	68.897 50.964 68.929 51.028 ;
			RECT	69.065 50.964 69.097 51.028 ;
			RECT	69.233 50.964 69.265 51.028 ;
			RECT	69.401 50.964 69.433 51.028 ;
			RECT	69.569 50.964 69.601 51.028 ;
			RECT	69.737 50.964 69.769 51.028 ;
			RECT	69.905 50.964 69.937 51.028 ;
			RECT	70.073 50.964 70.105 51.028 ;
			RECT	70.241 50.964 70.273 51.028 ;
			RECT	70.409 50.964 70.441 51.028 ;
			RECT	70.577 50.964 70.609 51.028 ;
			RECT	70.745 50.964 70.777 51.028 ;
			RECT	70.913 50.964 70.945 51.028 ;
			RECT	71.081 50.964 71.113 51.028 ;
			RECT	71.249 50.964 71.281 51.028 ;
			RECT	71.417 50.964 71.449 51.028 ;
			RECT	71.585 50.964 71.617 51.028 ;
			RECT	71.753 50.964 71.785 51.028 ;
			RECT	71.921 50.964 71.953 51.028 ;
			RECT	72.089 50.964 72.121 51.028 ;
			RECT	72.257 50.964 72.289 51.028 ;
			RECT	72.425 50.964 72.457 51.028 ;
			RECT	72.593 50.964 72.625 51.028 ;
			RECT	72.761 50.964 72.793 51.028 ;
			RECT	72.929 50.964 72.961 51.028 ;
			RECT	73.097 50.964 73.129 51.028 ;
			RECT	73.265 50.964 73.297 51.028 ;
			RECT	73.433 50.964 73.465 51.028 ;
			RECT	73.601 50.964 73.633 51.028 ;
			RECT	73.769 50.964 73.801 51.028 ;
			RECT	73.937 50.964 73.969 51.028 ;
			RECT	74.105 50.964 74.137 51.028 ;
			RECT	74.273 50.964 74.305 51.028 ;
			RECT	74.441 50.964 74.473 51.028 ;
			RECT	74.609 50.964 74.641 51.028 ;
			RECT	74.777 50.964 74.809 51.028 ;
			RECT	74.945 50.964 74.977 51.028 ;
			RECT	75.113 50.964 75.145 51.028 ;
			RECT	75.281 50.964 75.313 51.028 ;
			RECT	75.449 50.964 75.481 51.028 ;
			RECT	75.617 50.964 75.649 51.028 ;
			RECT	75.785 50.964 75.817 51.028 ;
			RECT	75.953 50.964 75.985 51.028 ;
			RECT	76.121 50.964 76.153 51.028 ;
			RECT	76.289 50.964 76.321 51.028 ;
			RECT	76.457 50.964 76.489 51.028 ;
			RECT	76.625 50.964 76.657 51.028 ;
			RECT	76.793 50.964 76.825 51.028 ;
			RECT	76.961 50.964 76.993 51.028 ;
			RECT	77.129 50.964 77.161 51.028 ;
			RECT	77.297 50.964 77.329 51.028 ;
			RECT	77.465 50.964 77.497 51.028 ;
			RECT	77.633 50.964 77.665 51.028 ;
			RECT	77.801 50.964 77.833 51.028 ;
			RECT	77.969 50.964 78.001 51.028 ;
			RECT	78.137 50.964 78.169 51.028 ;
			RECT	78.305 50.964 78.337 51.028 ;
			RECT	78.473 50.964 78.505 51.028 ;
			RECT	78.641 50.964 78.673 51.028 ;
			RECT	78.809 50.964 78.841 51.028 ;
			RECT	78.977 50.964 79.009 51.028 ;
			RECT	79.145 50.964 79.177 51.028 ;
			RECT	79.313 50.964 79.345 51.028 ;
			RECT	79.481 50.964 79.513 51.028 ;
			RECT	79.649 50.964 79.681 51.028 ;
			RECT	79.817 50.964 79.849 51.028 ;
			RECT	79.985 50.964 80.017 51.028 ;
			RECT	80.153 50.964 80.185 51.028 ;
			RECT	80.321 50.964 80.353 51.028 ;
			RECT	80.489 50.964 80.521 51.028 ;
			RECT	80.657 50.964 80.689 51.028 ;
			RECT	80.825 50.964 80.857 51.028 ;
			RECT	80.993 50.964 81.025 51.028 ;
			RECT	81.161 50.964 81.193 51.028 ;
			RECT	81.329 50.964 81.361 51.028 ;
			RECT	81.497 50.964 81.529 51.028 ;
			RECT	81.665 50.964 81.697 51.028 ;
			RECT	81.833 50.964 81.865 51.028 ;
			RECT	82.001 50.964 82.033 51.028 ;
			RECT	82.169 50.964 82.201 51.028 ;
			RECT	82.337 50.964 82.369 51.028 ;
			RECT	82.505 50.964 82.537 51.028 ;
			RECT	82.673 50.964 82.705 51.028 ;
			RECT	82.841 50.964 82.873 51.028 ;
			RECT	83.009 50.964 83.041 51.028 ;
			RECT	83.177 50.964 83.209 51.028 ;
			RECT	83.345 50.964 83.377 51.028 ;
			RECT	83.513 50.964 83.545 51.028 ;
			RECT	83.681 50.964 83.713 51.028 ;
			RECT	83.849 50.964 83.881 51.028 ;
			RECT	84.017 50.964 84.049 51.028 ;
			RECT	84.185 50.964 84.217 51.028 ;
			RECT	84.353 50.964 84.385 51.028 ;
			RECT	84.521 50.964 84.553 51.028 ;
			RECT	84.689 50.964 84.721 51.028 ;
			RECT	84.857 50.964 84.889 51.028 ;
			RECT	85.025 50.964 85.057 51.028 ;
			RECT	85.193 50.964 85.225 51.028 ;
			RECT	85.361 50.964 85.393 51.028 ;
			RECT	85.529 50.964 85.561 51.028 ;
			RECT	85.697 50.964 85.729 51.028 ;
			RECT	85.865 50.964 85.897 51.028 ;
			RECT	86.033 50.964 86.065 51.028 ;
			RECT	86.201 50.964 86.233 51.028 ;
			RECT	86.369 50.964 86.401 51.028 ;
			RECT	86.537 50.964 86.569 51.028 ;
			RECT	86.705 50.964 86.737 51.028 ;
			RECT	86.873 50.964 86.905 51.028 ;
			RECT	87.041 50.964 87.073 51.028 ;
			RECT	87.209 50.964 87.241 51.028 ;
			RECT	87.377 50.964 87.409 51.028 ;
			RECT	87.545 50.964 87.577 51.028 ;
			RECT	87.713 50.964 87.745 51.028 ;
			RECT	87.881 50.964 87.913 51.028 ;
			RECT	88.049 50.964 88.081 51.028 ;
			RECT	88.217 50.964 88.249 51.028 ;
			RECT	88.385 50.964 88.417 51.028 ;
			RECT	88.553 50.964 88.585 51.028 ;
			RECT	88.721 50.964 88.753 51.028 ;
			RECT	88.889 50.964 88.921 51.028 ;
			RECT	89.057 50.964 89.089 51.028 ;
			RECT	89.225 50.964 89.257 51.028 ;
			RECT	89.393 50.964 89.425 51.028 ;
			RECT	89.561 50.964 89.593 51.028 ;
			RECT	89.729 50.964 89.761 51.028 ;
			RECT	89.897 50.964 89.929 51.028 ;
			RECT	90.065 50.964 90.097 51.028 ;
			RECT	90.233 50.964 90.265 51.028 ;
			RECT	90.401 50.964 90.433 51.028 ;
			RECT	90.569 50.964 90.601 51.028 ;
			RECT	90.737 50.964 90.769 51.028 ;
			RECT	90.905 50.964 90.937 51.028 ;
			RECT	91.073 50.964 91.105 51.028 ;
			RECT	91.241 50.964 91.273 51.028 ;
			RECT	91.409 50.964 91.441 51.028 ;
			RECT	91.577 50.964 91.609 51.028 ;
			RECT	91.745 50.964 91.777 51.028 ;
			RECT	91.913 50.964 91.945 51.028 ;
			RECT	92.081 50.964 92.113 51.028 ;
			RECT	92.249 50.964 92.281 51.028 ;
			RECT	92.417 50.964 92.449 51.028 ;
			RECT	92.585 50.964 92.617 51.028 ;
			RECT	92.753 50.964 92.785 51.028 ;
			RECT	92.921 50.964 92.953 51.028 ;
			RECT	93.089 50.964 93.121 51.028 ;
			RECT	93.257 50.964 93.289 51.028 ;
			RECT	93.425 50.964 93.457 51.028 ;
			RECT	93.593 50.964 93.625 51.028 ;
			RECT	93.761 50.964 93.793 51.028 ;
			RECT	93.929 50.964 93.961 51.028 ;
			RECT	94.097 50.964 94.129 51.028 ;
			RECT	94.265 50.964 94.297 51.028 ;
			RECT	94.433 50.964 94.465 51.028 ;
			RECT	94.601 50.964 94.633 51.028 ;
			RECT	94.769 50.964 94.801 51.028 ;
			RECT	94.937 50.964 94.969 51.028 ;
			RECT	95.105 50.964 95.137 51.028 ;
			RECT	95.273 50.964 95.305 51.028 ;
			RECT	95.441 50.964 95.473 51.028 ;
			RECT	95.609 50.964 95.641 51.028 ;
			RECT	95.777 50.964 95.809 51.028 ;
			RECT	95.945 50.964 95.977 51.028 ;
			RECT	96.113 50.964 96.145 51.028 ;
			RECT	96.281 50.964 96.313 51.028 ;
			RECT	96.449 50.964 96.481 51.028 ;
			RECT	96.617 50.964 96.649 51.028 ;
			RECT	96.785 50.964 96.817 51.028 ;
			RECT	96.953 50.964 96.985 51.028 ;
			RECT	97.121 50.964 97.153 51.028 ;
			RECT	97.289 50.964 97.321 51.028 ;
			RECT	97.457 50.964 97.489 51.028 ;
			RECT	97.625 50.964 97.657 51.028 ;
			RECT	97.793 50.964 97.825 51.028 ;
			RECT	97.961 50.964 97.993 51.028 ;
			RECT	98.129 50.964 98.161 51.028 ;
			RECT	98.297 50.964 98.329 51.028 ;
			RECT	98.465 50.964 98.497 51.028 ;
			RECT	98.633 50.964 98.665 51.028 ;
			RECT	98.801 50.964 98.833 51.028 ;
			RECT	98.969 50.964 99.001 51.028 ;
			RECT	99.137 50.964 99.169 51.028 ;
			RECT	99.305 50.964 99.337 51.028 ;
			RECT	99.473 50.964 99.505 51.028 ;
			RECT	99.641 50.964 99.673 51.028 ;
			RECT	99.809 50.964 99.841 51.028 ;
			RECT	99.977 50.964 100.009 51.028 ;
			RECT	100.145 50.964 100.177 51.028 ;
			RECT	100.313 50.964 100.345 51.028 ;
			RECT	100.481 50.964 100.513 51.028 ;
			RECT	100.649 50.964 100.681 51.028 ;
			RECT	100.817 50.964 100.849 51.028 ;
			RECT	100.985 50.964 101.017 51.028 ;
			RECT	101.153 50.964 101.185 51.028 ;
			RECT	101.321 50.964 101.353 51.028 ;
			RECT	101.489 50.964 101.521 51.028 ;
			RECT	101.657 50.964 101.689 51.028 ;
			RECT	101.825 50.964 101.857 51.028 ;
			RECT	101.993 50.964 102.025 51.028 ;
			RECT	102.123 50.98 102.155 51.012 ;
			RECT	102.245 50.975 102.277 51.007 ;
			RECT	102.375 50.964 102.407 51.028 ;
			RECT	103.795 50.964 103.827 51.028 ;
			RECT	103.925 50.975 103.957 51.007 ;
			RECT	104.047 50.98 104.079 51.012 ;
			RECT	104.177 50.964 104.209 51.028 ;
			RECT	104.345 50.964 104.377 51.028 ;
			RECT	104.513 50.964 104.545 51.028 ;
			RECT	104.681 50.964 104.713 51.028 ;
			RECT	104.849 50.964 104.881 51.028 ;
			RECT	105.017 50.964 105.049 51.028 ;
			RECT	105.185 50.964 105.217 51.028 ;
			RECT	105.353 50.964 105.385 51.028 ;
			RECT	105.521 50.964 105.553 51.028 ;
			RECT	105.689 50.964 105.721 51.028 ;
			RECT	105.857 50.964 105.889 51.028 ;
			RECT	106.025 50.964 106.057 51.028 ;
			RECT	106.193 50.964 106.225 51.028 ;
			RECT	106.361 50.964 106.393 51.028 ;
			RECT	106.529 50.964 106.561 51.028 ;
			RECT	106.697 50.964 106.729 51.028 ;
			RECT	106.865 50.964 106.897 51.028 ;
			RECT	107.033 50.964 107.065 51.028 ;
			RECT	107.201 50.964 107.233 51.028 ;
			RECT	107.369 50.964 107.401 51.028 ;
			RECT	107.537 50.964 107.569 51.028 ;
			RECT	107.705 50.964 107.737 51.028 ;
			RECT	107.873 50.964 107.905 51.028 ;
			RECT	108.041 50.964 108.073 51.028 ;
			RECT	108.209 50.964 108.241 51.028 ;
			RECT	108.377 50.964 108.409 51.028 ;
			RECT	108.545 50.964 108.577 51.028 ;
			RECT	108.713 50.964 108.745 51.028 ;
			RECT	108.881 50.964 108.913 51.028 ;
			RECT	109.049 50.964 109.081 51.028 ;
			RECT	109.217 50.964 109.249 51.028 ;
			RECT	109.385 50.964 109.417 51.028 ;
			RECT	109.553 50.964 109.585 51.028 ;
			RECT	109.721 50.964 109.753 51.028 ;
			RECT	109.889 50.964 109.921 51.028 ;
			RECT	110.057 50.964 110.089 51.028 ;
			RECT	110.225 50.964 110.257 51.028 ;
			RECT	110.393 50.964 110.425 51.028 ;
			RECT	110.561 50.964 110.593 51.028 ;
			RECT	110.729 50.964 110.761 51.028 ;
			RECT	110.897 50.964 110.929 51.028 ;
			RECT	111.065 50.964 111.097 51.028 ;
			RECT	111.233 50.964 111.265 51.028 ;
			RECT	111.401 50.964 111.433 51.028 ;
			RECT	111.569 50.964 111.601 51.028 ;
			RECT	111.737 50.964 111.769 51.028 ;
			RECT	111.905 50.964 111.937 51.028 ;
			RECT	112.073 50.964 112.105 51.028 ;
			RECT	112.241 50.964 112.273 51.028 ;
			RECT	112.409 50.964 112.441 51.028 ;
			RECT	112.577 50.964 112.609 51.028 ;
			RECT	112.745 50.964 112.777 51.028 ;
			RECT	112.913 50.964 112.945 51.028 ;
			RECT	113.081 50.964 113.113 51.028 ;
			RECT	113.249 50.964 113.281 51.028 ;
			RECT	113.417 50.964 113.449 51.028 ;
			RECT	113.585 50.964 113.617 51.028 ;
			RECT	113.753 50.964 113.785 51.028 ;
			RECT	113.921 50.964 113.953 51.028 ;
			RECT	114.089 50.964 114.121 51.028 ;
			RECT	114.257 50.964 114.289 51.028 ;
			RECT	114.425 50.964 114.457 51.028 ;
			RECT	114.593 50.964 114.625 51.028 ;
			RECT	114.761 50.964 114.793 51.028 ;
			RECT	114.929 50.964 114.961 51.028 ;
			RECT	115.097 50.964 115.129 51.028 ;
			RECT	115.265 50.964 115.297 51.028 ;
			RECT	115.433 50.964 115.465 51.028 ;
			RECT	115.601 50.964 115.633 51.028 ;
			RECT	115.769 50.964 115.801 51.028 ;
			RECT	115.937 50.964 115.969 51.028 ;
			RECT	116.105 50.964 116.137 51.028 ;
			RECT	116.273 50.964 116.305 51.028 ;
			RECT	116.441 50.964 116.473 51.028 ;
			RECT	116.609 50.964 116.641 51.028 ;
			RECT	116.777 50.964 116.809 51.028 ;
			RECT	116.945 50.964 116.977 51.028 ;
			RECT	117.113 50.964 117.145 51.028 ;
			RECT	117.281 50.964 117.313 51.028 ;
			RECT	117.449 50.964 117.481 51.028 ;
			RECT	117.617 50.964 117.649 51.028 ;
			RECT	117.785 50.964 117.817 51.028 ;
			RECT	117.953 50.964 117.985 51.028 ;
			RECT	118.121 50.964 118.153 51.028 ;
			RECT	118.289 50.964 118.321 51.028 ;
			RECT	118.457 50.964 118.489 51.028 ;
			RECT	118.625 50.964 118.657 51.028 ;
			RECT	118.793 50.964 118.825 51.028 ;
			RECT	118.961 50.964 118.993 51.028 ;
			RECT	119.129 50.964 119.161 51.028 ;
			RECT	119.297 50.964 119.329 51.028 ;
			RECT	119.465 50.964 119.497 51.028 ;
			RECT	119.633 50.964 119.665 51.028 ;
			RECT	119.801 50.964 119.833 51.028 ;
			RECT	119.969 50.964 120.001 51.028 ;
			RECT	120.137 50.964 120.169 51.028 ;
			RECT	120.305 50.964 120.337 51.028 ;
			RECT	120.473 50.964 120.505 51.028 ;
			RECT	120.641 50.964 120.673 51.028 ;
			RECT	120.809 50.964 120.841 51.028 ;
			RECT	120.977 50.964 121.009 51.028 ;
			RECT	121.145 50.964 121.177 51.028 ;
			RECT	121.313 50.964 121.345 51.028 ;
			RECT	121.481 50.964 121.513 51.028 ;
			RECT	121.649 50.964 121.681 51.028 ;
			RECT	121.817 50.964 121.849 51.028 ;
			RECT	121.985 50.964 122.017 51.028 ;
			RECT	122.153 50.964 122.185 51.028 ;
			RECT	122.321 50.964 122.353 51.028 ;
			RECT	122.489 50.964 122.521 51.028 ;
			RECT	122.657 50.964 122.689 51.028 ;
			RECT	122.825 50.964 122.857 51.028 ;
			RECT	122.993 50.964 123.025 51.028 ;
			RECT	123.161 50.964 123.193 51.028 ;
			RECT	123.329 50.964 123.361 51.028 ;
			RECT	123.497 50.964 123.529 51.028 ;
			RECT	123.665 50.964 123.697 51.028 ;
			RECT	123.833 50.964 123.865 51.028 ;
			RECT	124.001 50.964 124.033 51.028 ;
			RECT	124.169 50.964 124.201 51.028 ;
			RECT	124.337 50.964 124.369 51.028 ;
			RECT	124.505 50.964 124.537 51.028 ;
			RECT	124.673 50.964 124.705 51.028 ;
			RECT	124.841 50.964 124.873 51.028 ;
			RECT	125.009 50.964 125.041 51.028 ;
			RECT	125.177 50.964 125.209 51.028 ;
			RECT	125.345 50.964 125.377 51.028 ;
			RECT	125.513 50.964 125.545 51.028 ;
			RECT	125.681 50.964 125.713 51.028 ;
			RECT	125.849 50.964 125.881 51.028 ;
			RECT	126.017 50.964 126.049 51.028 ;
			RECT	126.185 50.964 126.217 51.028 ;
			RECT	126.353 50.964 126.385 51.028 ;
			RECT	126.521 50.964 126.553 51.028 ;
			RECT	126.689 50.964 126.721 51.028 ;
			RECT	126.857 50.964 126.889 51.028 ;
			RECT	127.025 50.964 127.057 51.028 ;
			RECT	127.193 50.964 127.225 51.028 ;
			RECT	127.361 50.964 127.393 51.028 ;
			RECT	127.529 50.964 127.561 51.028 ;
			RECT	127.697 50.964 127.729 51.028 ;
			RECT	127.865 50.964 127.897 51.028 ;
			RECT	128.033 50.964 128.065 51.028 ;
			RECT	128.201 50.964 128.233 51.028 ;
			RECT	128.369 50.964 128.401 51.028 ;
			RECT	128.537 50.964 128.569 51.028 ;
			RECT	128.705 50.964 128.737 51.028 ;
			RECT	128.873 50.964 128.905 51.028 ;
			RECT	129.041 50.964 129.073 51.028 ;
			RECT	129.209 50.964 129.241 51.028 ;
			RECT	129.377 50.964 129.409 51.028 ;
			RECT	129.545 50.964 129.577 51.028 ;
			RECT	129.713 50.964 129.745 51.028 ;
			RECT	129.881 50.964 129.913 51.028 ;
			RECT	130.049 50.964 130.081 51.028 ;
			RECT	130.217 50.964 130.249 51.028 ;
			RECT	130.385 50.964 130.417 51.028 ;
			RECT	130.553 50.964 130.585 51.028 ;
			RECT	130.721 50.964 130.753 51.028 ;
			RECT	130.889 50.964 130.921 51.028 ;
			RECT	131.057 50.964 131.089 51.028 ;
			RECT	131.225 50.964 131.257 51.028 ;
			RECT	131.393 50.964 131.425 51.028 ;
			RECT	131.561 50.964 131.593 51.028 ;
			RECT	131.729 50.964 131.761 51.028 ;
			RECT	131.897 50.964 131.929 51.028 ;
			RECT	132.065 50.964 132.097 51.028 ;
			RECT	132.233 50.964 132.265 51.028 ;
			RECT	132.401 50.964 132.433 51.028 ;
			RECT	132.569 50.964 132.601 51.028 ;
			RECT	132.737 50.964 132.769 51.028 ;
			RECT	132.905 50.964 132.937 51.028 ;
			RECT	133.073 50.964 133.105 51.028 ;
			RECT	133.241 50.964 133.273 51.028 ;
			RECT	133.409 50.964 133.441 51.028 ;
			RECT	133.577 50.964 133.609 51.028 ;
			RECT	133.745 50.964 133.777 51.028 ;
			RECT	133.913 50.964 133.945 51.028 ;
			RECT	134.081 50.964 134.113 51.028 ;
			RECT	134.249 50.964 134.281 51.028 ;
			RECT	134.417 50.964 134.449 51.028 ;
			RECT	134.585 50.964 134.617 51.028 ;
			RECT	134.753 50.964 134.785 51.028 ;
			RECT	134.921 50.964 134.953 51.028 ;
			RECT	135.089 50.964 135.121 51.028 ;
			RECT	135.257 50.964 135.289 51.028 ;
			RECT	135.425 50.964 135.457 51.028 ;
			RECT	135.593 50.964 135.625 51.028 ;
			RECT	135.761 50.964 135.793 51.028 ;
			RECT	135.929 50.964 135.961 51.028 ;
			RECT	136.097 50.964 136.129 51.028 ;
			RECT	136.265 50.964 136.297 51.028 ;
			RECT	136.433 50.964 136.465 51.028 ;
			RECT	136.601 50.964 136.633 51.028 ;
			RECT	136.769 50.964 136.801 51.028 ;
			RECT	136.937 50.964 136.969 51.028 ;
			RECT	137.105 50.964 137.137 51.028 ;
			RECT	137.273 50.964 137.305 51.028 ;
			RECT	137.441 50.964 137.473 51.028 ;
			RECT	137.609 50.964 137.641 51.028 ;
			RECT	137.777 50.964 137.809 51.028 ;
			RECT	137.945 50.964 137.977 51.028 ;
			RECT	138.113 50.964 138.145 51.028 ;
			RECT	138.281 50.964 138.313 51.028 ;
			RECT	138.449 50.964 138.481 51.028 ;
			RECT	138.617 50.964 138.649 51.028 ;
			RECT	138.785 50.964 138.817 51.028 ;
			RECT	138.953 50.964 138.985 51.028 ;
			RECT	139.121 50.964 139.153 51.028 ;
			RECT	139.289 50.964 139.321 51.028 ;
			RECT	139.457 50.964 139.489 51.028 ;
			RECT	139.625 50.964 139.657 51.028 ;
			RECT	139.793 50.964 139.825 51.028 ;
			RECT	139.961 50.964 139.993 51.028 ;
			RECT	140.129 50.964 140.161 51.028 ;
			RECT	140.297 50.964 140.329 51.028 ;
			RECT	140.465 50.964 140.497 51.028 ;
			RECT	140.633 50.964 140.665 51.028 ;
			RECT	140.801 50.964 140.833 51.028 ;
			RECT	140.969 50.964 141.001 51.028 ;
			RECT	141.137 50.964 141.169 51.028 ;
			RECT	141.305 50.964 141.337 51.028 ;
			RECT	141.473 50.964 141.505 51.028 ;
			RECT	141.641 50.964 141.673 51.028 ;
			RECT	141.809 50.964 141.841 51.028 ;
			RECT	141.977 50.964 142.009 51.028 ;
			RECT	142.145 50.964 142.177 51.028 ;
			RECT	142.313 50.964 142.345 51.028 ;
			RECT	142.481 50.964 142.513 51.028 ;
			RECT	142.649 50.964 142.681 51.028 ;
			RECT	142.817 50.964 142.849 51.028 ;
			RECT	142.985 50.964 143.017 51.028 ;
			RECT	143.153 50.964 143.185 51.028 ;
			RECT	143.321 50.964 143.353 51.028 ;
			RECT	143.489 50.964 143.521 51.028 ;
			RECT	143.657 50.964 143.689 51.028 ;
			RECT	143.825 50.964 143.857 51.028 ;
			RECT	143.993 50.964 144.025 51.028 ;
			RECT	144.161 50.964 144.193 51.028 ;
			RECT	144.329 50.964 144.361 51.028 ;
			RECT	144.497 50.964 144.529 51.028 ;
			RECT	144.665 50.964 144.697 51.028 ;
			RECT	144.833 50.964 144.865 51.028 ;
			RECT	145.001 50.964 145.033 51.028 ;
			RECT	145.169 50.964 145.201 51.028 ;
			RECT	145.337 50.964 145.369 51.028 ;
			RECT	145.505 50.964 145.537 51.028 ;
			RECT	145.673 50.964 145.705 51.028 ;
			RECT	145.841 50.964 145.873 51.028 ;
			RECT	146.009 50.964 146.041 51.028 ;
			RECT	146.177 50.964 146.209 51.028 ;
			RECT	146.345 50.964 146.377 51.028 ;
			RECT	146.513 50.964 146.545 51.028 ;
			RECT	146.681 50.964 146.713 51.028 ;
			RECT	146.849 50.964 146.881 51.028 ;
			RECT	147.017 50.964 147.049 51.028 ;
			RECT	147.185 50.964 147.217 51.028 ;
			RECT	147.316 50.98 147.348 51.012 ;
			RECT	147.437 50.98 147.469 51.012 ;
			RECT	147.567 50.964 147.599 51.028 ;
			RECT	149.879 50.964 149.911 51.028 ;
			RECT	151.13 50.964 151.194 51.028 ;
			RECT	151.81 50.964 151.842 51.028 ;
			RECT	152.249 50.964 152.281 51.028 ;
			RECT	153.56 50.964 153.624 51.028 ;
			RECT	156.601 50.964 156.633 51.028 ;
			RECT	156.731 50.98 156.763 51.012 ;
			RECT	156.852 50.98 156.884 51.012 ;
			RECT	156.983 50.964 157.015 51.028 ;
			RECT	157.151 50.964 157.183 51.028 ;
			RECT	157.319 50.964 157.351 51.028 ;
			RECT	157.487 50.964 157.519 51.028 ;
			RECT	157.655 50.964 157.687 51.028 ;
			RECT	157.823 50.964 157.855 51.028 ;
			RECT	157.991 50.964 158.023 51.028 ;
			RECT	158.159 50.964 158.191 51.028 ;
			RECT	158.327 50.964 158.359 51.028 ;
			RECT	158.495 50.964 158.527 51.028 ;
			RECT	158.663 50.964 158.695 51.028 ;
			RECT	158.831 50.964 158.863 51.028 ;
			RECT	158.999 50.964 159.031 51.028 ;
			RECT	159.167 50.964 159.199 51.028 ;
			RECT	159.335 50.964 159.367 51.028 ;
			RECT	159.503 50.964 159.535 51.028 ;
			RECT	159.671 50.964 159.703 51.028 ;
			RECT	159.839 50.964 159.871 51.028 ;
			RECT	160.007 50.964 160.039 51.028 ;
			RECT	160.175 50.964 160.207 51.028 ;
			RECT	160.343 50.964 160.375 51.028 ;
			RECT	160.511 50.964 160.543 51.028 ;
			RECT	160.679 50.964 160.711 51.028 ;
			RECT	160.847 50.964 160.879 51.028 ;
			RECT	161.015 50.964 161.047 51.028 ;
			RECT	161.183 50.964 161.215 51.028 ;
			RECT	161.351 50.964 161.383 51.028 ;
			RECT	161.519 50.964 161.551 51.028 ;
			RECT	161.687 50.964 161.719 51.028 ;
			RECT	161.855 50.964 161.887 51.028 ;
			RECT	162.023 50.964 162.055 51.028 ;
			RECT	162.191 50.964 162.223 51.028 ;
			RECT	162.359 50.964 162.391 51.028 ;
			RECT	162.527 50.964 162.559 51.028 ;
			RECT	162.695 50.964 162.727 51.028 ;
			RECT	162.863 50.964 162.895 51.028 ;
			RECT	163.031 50.964 163.063 51.028 ;
			RECT	163.199 50.964 163.231 51.028 ;
			RECT	163.367 50.964 163.399 51.028 ;
			RECT	163.535 50.964 163.567 51.028 ;
			RECT	163.703 50.964 163.735 51.028 ;
			RECT	163.871 50.964 163.903 51.028 ;
			RECT	164.039 50.964 164.071 51.028 ;
			RECT	164.207 50.964 164.239 51.028 ;
			RECT	164.375 50.964 164.407 51.028 ;
			RECT	164.543 50.964 164.575 51.028 ;
			RECT	164.711 50.964 164.743 51.028 ;
			RECT	164.879 50.964 164.911 51.028 ;
			RECT	165.047 50.964 165.079 51.028 ;
			RECT	165.215 50.964 165.247 51.028 ;
			RECT	165.383 50.964 165.415 51.028 ;
			RECT	165.551 50.964 165.583 51.028 ;
			RECT	165.719 50.964 165.751 51.028 ;
			RECT	165.887 50.964 165.919 51.028 ;
			RECT	166.055 50.964 166.087 51.028 ;
			RECT	166.223 50.964 166.255 51.028 ;
			RECT	166.391 50.964 166.423 51.028 ;
			RECT	166.559 50.964 166.591 51.028 ;
			RECT	166.727 50.964 166.759 51.028 ;
			RECT	166.895 50.964 166.927 51.028 ;
			RECT	167.063 50.964 167.095 51.028 ;
			RECT	167.231 50.964 167.263 51.028 ;
			RECT	167.399 50.964 167.431 51.028 ;
			RECT	167.567 50.964 167.599 51.028 ;
			RECT	167.735 50.964 167.767 51.028 ;
			RECT	167.903 50.964 167.935 51.028 ;
			RECT	168.071 50.964 168.103 51.028 ;
			RECT	168.239 50.964 168.271 51.028 ;
			RECT	168.407 50.964 168.439 51.028 ;
			RECT	168.575 50.964 168.607 51.028 ;
			RECT	168.743 50.964 168.775 51.028 ;
			RECT	168.911 50.964 168.943 51.028 ;
			RECT	169.079 50.964 169.111 51.028 ;
			RECT	169.247 50.964 169.279 51.028 ;
			RECT	169.415 50.964 169.447 51.028 ;
			RECT	169.583 50.964 169.615 51.028 ;
			RECT	169.751 50.964 169.783 51.028 ;
			RECT	169.919 50.964 169.951 51.028 ;
			RECT	170.087 50.964 170.119 51.028 ;
			RECT	170.255 50.964 170.287 51.028 ;
			RECT	170.423 50.964 170.455 51.028 ;
			RECT	170.591 50.964 170.623 51.028 ;
			RECT	170.759 50.964 170.791 51.028 ;
			RECT	170.927 50.964 170.959 51.028 ;
			RECT	171.095 50.964 171.127 51.028 ;
			RECT	171.263 50.964 171.295 51.028 ;
			RECT	171.431 50.964 171.463 51.028 ;
			RECT	171.599 50.964 171.631 51.028 ;
			RECT	171.767 50.964 171.799 51.028 ;
			RECT	171.935 50.964 171.967 51.028 ;
			RECT	172.103 50.964 172.135 51.028 ;
			RECT	172.271 50.964 172.303 51.028 ;
			RECT	172.439 50.964 172.471 51.028 ;
			RECT	172.607 50.964 172.639 51.028 ;
			RECT	172.775 50.964 172.807 51.028 ;
			RECT	172.943 50.964 172.975 51.028 ;
			RECT	173.111 50.964 173.143 51.028 ;
			RECT	173.279 50.964 173.311 51.028 ;
			RECT	173.447 50.964 173.479 51.028 ;
			RECT	173.615 50.964 173.647 51.028 ;
			RECT	173.783 50.964 173.815 51.028 ;
			RECT	173.951 50.964 173.983 51.028 ;
			RECT	174.119 50.964 174.151 51.028 ;
			RECT	174.287 50.964 174.319 51.028 ;
			RECT	174.455 50.964 174.487 51.028 ;
			RECT	174.623 50.964 174.655 51.028 ;
			RECT	174.791 50.964 174.823 51.028 ;
			RECT	174.959 50.964 174.991 51.028 ;
			RECT	175.127 50.964 175.159 51.028 ;
			RECT	175.295 50.964 175.327 51.028 ;
			RECT	175.463 50.964 175.495 51.028 ;
			RECT	175.631 50.964 175.663 51.028 ;
			RECT	175.799 50.964 175.831 51.028 ;
			RECT	175.967 50.964 175.999 51.028 ;
			RECT	176.135 50.964 176.167 51.028 ;
			RECT	176.303 50.964 176.335 51.028 ;
			RECT	176.471 50.964 176.503 51.028 ;
			RECT	176.639 50.964 176.671 51.028 ;
			RECT	176.807 50.964 176.839 51.028 ;
			RECT	176.975 50.964 177.007 51.028 ;
			RECT	177.143 50.964 177.175 51.028 ;
			RECT	177.311 50.964 177.343 51.028 ;
			RECT	177.479 50.964 177.511 51.028 ;
			RECT	177.647 50.964 177.679 51.028 ;
			RECT	177.815 50.964 177.847 51.028 ;
			RECT	177.983 50.964 178.015 51.028 ;
			RECT	178.151 50.964 178.183 51.028 ;
			RECT	178.319 50.964 178.351 51.028 ;
			RECT	178.487 50.964 178.519 51.028 ;
			RECT	178.655 50.964 178.687 51.028 ;
			RECT	178.823 50.964 178.855 51.028 ;
			RECT	178.991 50.964 179.023 51.028 ;
			RECT	179.159 50.964 179.191 51.028 ;
			RECT	179.327 50.964 179.359 51.028 ;
			RECT	179.495 50.964 179.527 51.028 ;
			RECT	179.663 50.964 179.695 51.028 ;
			RECT	179.831 50.964 179.863 51.028 ;
			RECT	179.999 50.964 180.031 51.028 ;
			RECT	180.167 50.964 180.199 51.028 ;
			RECT	180.335 50.964 180.367 51.028 ;
			RECT	180.503 50.964 180.535 51.028 ;
			RECT	180.671 50.964 180.703 51.028 ;
			RECT	180.839 50.964 180.871 51.028 ;
			RECT	181.007 50.964 181.039 51.028 ;
			RECT	181.175 50.964 181.207 51.028 ;
			RECT	181.343 50.964 181.375 51.028 ;
			RECT	181.511 50.964 181.543 51.028 ;
			RECT	181.679 50.964 181.711 51.028 ;
			RECT	181.847 50.964 181.879 51.028 ;
			RECT	182.015 50.964 182.047 51.028 ;
			RECT	182.183 50.964 182.215 51.028 ;
			RECT	182.351 50.964 182.383 51.028 ;
			RECT	182.519 50.964 182.551 51.028 ;
			RECT	182.687 50.964 182.719 51.028 ;
			RECT	182.855 50.964 182.887 51.028 ;
			RECT	183.023 50.964 183.055 51.028 ;
			RECT	183.191 50.964 183.223 51.028 ;
			RECT	183.359 50.964 183.391 51.028 ;
			RECT	183.527 50.964 183.559 51.028 ;
			RECT	183.695 50.964 183.727 51.028 ;
			RECT	183.863 50.964 183.895 51.028 ;
			RECT	184.031 50.964 184.063 51.028 ;
			RECT	184.199 50.964 184.231 51.028 ;
			RECT	184.367 50.964 184.399 51.028 ;
			RECT	184.535 50.964 184.567 51.028 ;
			RECT	184.703 50.964 184.735 51.028 ;
			RECT	184.871 50.964 184.903 51.028 ;
			RECT	185.039 50.964 185.071 51.028 ;
			RECT	185.207 50.964 185.239 51.028 ;
			RECT	185.375 50.964 185.407 51.028 ;
			RECT	185.543 50.964 185.575 51.028 ;
			RECT	185.711 50.964 185.743 51.028 ;
			RECT	185.879 50.964 185.911 51.028 ;
			RECT	186.047 50.964 186.079 51.028 ;
			RECT	186.215 50.964 186.247 51.028 ;
			RECT	186.383 50.964 186.415 51.028 ;
			RECT	186.551 50.964 186.583 51.028 ;
			RECT	186.719 50.964 186.751 51.028 ;
			RECT	186.887 50.964 186.919 51.028 ;
			RECT	187.055 50.964 187.087 51.028 ;
			RECT	187.223 50.964 187.255 51.028 ;
			RECT	187.391 50.964 187.423 51.028 ;
			RECT	187.559 50.964 187.591 51.028 ;
			RECT	187.727 50.964 187.759 51.028 ;
			RECT	187.895 50.964 187.927 51.028 ;
			RECT	188.063 50.964 188.095 51.028 ;
			RECT	188.231 50.964 188.263 51.028 ;
			RECT	188.399 50.964 188.431 51.028 ;
			RECT	188.567 50.964 188.599 51.028 ;
			RECT	188.735 50.964 188.767 51.028 ;
			RECT	188.903 50.964 188.935 51.028 ;
			RECT	189.071 50.964 189.103 51.028 ;
			RECT	189.239 50.964 189.271 51.028 ;
			RECT	189.407 50.964 189.439 51.028 ;
			RECT	189.575 50.964 189.607 51.028 ;
			RECT	189.743 50.964 189.775 51.028 ;
			RECT	189.911 50.964 189.943 51.028 ;
			RECT	190.079 50.964 190.111 51.028 ;
			RECT	190.247 50.964 190.279 51.028 ;
			RECT	190.415 50.964 190.447 51.028 ;
			RECT	190.583 50.964 190.615 51.028 ;
			RECT	190.751 50.964 190.783 51.028 ;
			RECT	190.919 50.964 190.951 51.028 ;
			RECT	191.087 50.964 191.119 51.028 ;
			RECT	191.255 50.964 191.287 51.028 ;
			RECT	191.423 50.964 191.455 51.028 ;
			RECT	191.591 50.964 191.623 51.028 ;
			RECT	191.759 50.964 191.791 51.028 ;
			RECT	191.927 50.964 191.959 51.028 ;
			RECT	192.095 50.964 192.127 51.028 ;
			RECT	192.263 50.964 192.295 51.028 ;
			RECT	192.431 50.964 192.463 51.028 ;
			RECT	192.599 50.964 192.631 51.028 ;
			RECT	192.767 50.964 192.799 51.028 ;
			RECT	192.935 50.964 192.967 51.028 ;
			RECT	193.103 50.964 193.135 51.028 ;
			RECT	193.271 50.964 193.303 51.028 ;
			RECT	193.439 50.964 193.471 51.028 ;
			RECT	193.607 50.964 193.639 51.028 ;
			RECT	193.775 50.964 193.807 51.028 ;
			RECT	193.943 50.964 193.975 51.028 ;
			RECT	194.111 50.964 194.143 51.028 ;
			RECT	194.279 50.964 194.311 51.028 ;
			RECT	194.447 50.964 194.479 51.028 ;
			RECT	194.615 50.964 194.647 51.028 ;
			RECT	194.783 50.964 194.815 51.028 ;
			RECT	194.951 50.964 194.983 51.028 ;
			RECT	195.119 50.964 195.151 51.028 ;
			RECT	195.287 50.964 195.319 51.028 ;
			RECT	195.455 50.964 195.487 51.028 ;
			RECT	195.623 50.964 195.655 51.028 ;
			RECT	195.791 50.964 195.823 51.028 ;
			RECT	195.959 50.964 195.991 51.028 ;
			RECT	196.127 50.964 196.159 51.028 ;
			RECT	196.295 50.964 196.327 51.028 ;
			RECT	196.463 50.964 196.495 51.028 ;
			RECT	196.631 50.964 196.663 51.028 ;
			RECT	196.799 50.964 196.831 51.028 ;
			RECT	196.967 50.964 196.999 51.028 ;
			RECT	197.135 50.964 197.167 51.028 ;
			RECT	197.303 50.964 197.335 51.028 ;
			RECT	197.471 50.964 197.503 51.028 ;
			RECT	197.639 50.964 197.671 51.028 ;
			RECT	197.807 50.964 197.839 51.028 ;
			RECT	197.975 50.964 198.007 51.028 ;
			RECT	198.143 50.964 198.175 51.028 ;
			RECT	198.311 50.964 198.343 51.028 ;
			RECT	198.479 50.964 198.511 51.028 ;
			RECT	198.647 50.964 198.679 51.028 ;
			RECT	198.815 50.964 198.847 51.028 ;
			RECT	198.983 50.964 199.015 51.028 ;
			RECT	199.151 50.964 199.183 51.028 ;
			RECT	199.319 50.964 199.351 51.028 ;
			RECT	199.487 50.964 199.519 51.028 ;
			RECT	199.655 50.964 199.687 51.028 ;
			RECT	199.823 50.964 199.855 51.028 ;
			RECT	199.991 50.964 200.023 51.028 ;
			RECT	200.121 50.98 200.153 51.012 ;
			RECT	200.243 50.975 200.275 51.007 ;
			RECT	200.373 50.964 200.405 51.028 ;
			RECT	200.9 50.964 200.932 51.028 ;
		END

		PORT
			LAYER	C4 ;
			RECT	0.294 77.816 201.665 77.936 ;
			LAYER	J3 ;
			RECT	0.755 77.844 0.787 77.908 ;
			RECT	1.645 77.844 1.709 77.908 ;
			RECT	2.323 77.844 2.387 77.908 ;
			RECT	3.438 77.844 3.47 77.908 ;
			RECT	3.585 77.844 3.617 77.908 ;
			RECT	4.195 77.844 4.227 77.908 ;
			RECT	4.72 77.844 4.752 77.908 ;
			RECT	4.944 77.844 5.008 77.908 ;
			RECT	5.267 77.844 5.299 77.908 ;
			RECT	5.797 77.844 5.829 77.908 ;
			RECT	5.927 77.855 5.959 77.887 ;
			RECT	6.049 77.86 6.081 77.892 ;
			RECT	6.179 77.844 6.211 77.908 ;
			RECT	6.347 77.844 6.379 77.908 ;
			RECT	6.515 77.844 6.547 77.908 ;
			RECT	6.683 77.844 6.715 77.908 ;
			RECT	6.851 77.844 6.883 77.908 ;
			RECT	7.019 77.844 7.051 77.908 ;
			RECT	7.187 77.844 7.219 77.908 ;
			RECT	7.355 77.844 7.387 77.908 ;
			RECT	7.523 77.844 7.555 77.908 ;
			RECT	7.691 77.844 7.723 77.908 ;
			RECT	7.859 77.844 7.891 77.908 ;
			RECT	8.027 77.844 8.059 77.908 ;
			RECT	8.195 77.844 8.227 77.908 ;
			RECT	8.363 77.844 8.395 77.908 ;
			RECT	8.531 77.844 8.563 77.908 ;
			RECT	8.699 77.844 8.731 77.908 ;
			RECT	8.867 77.844 8.899 77.908 ;
			RECT	9.035 77.844 9.067 77.908 ;
			RECT	9.203 77.844 9.235 77.908 ;
			RECT	9.371 77.844 9.403 77.908 ;
			RECT	9.539 77.844 9.571 77.908 ;
			RECT	9.707 77.844 9.739 77.908 ;
			RECT	9.875 77.844 9.907 77.908 ;
			RECT	10.043 77.844 10.075 77.908 ;
			RECT	10.211 77.844 10.243 77.908 ;
			RECT	10.379 77.844 10.411 77.908 ;
			RECT	10.547 77.844 10.579 77.908 ;
			RECT	10.715 77.844 10.747 77.908 ;
			RECT	10.883 77.844 10.915 77.908 ;
			RECT	11.051 77.844 11.083 77.908 ;
			RECT	11.219 77.844 11.251 77.908 ;
			RECT	11.387 77.844 11.419 77.908 ;
			RECT	11.555 77.844 11.587 77.908 ;
			RECT	11.723 77.844 11.755 77.908 ;
			RECT	11.891 77.844 11.923 77.908 ;
			RECT	12.059 77.844 12.091 77.908 ;
			RECT	12.227 77.844 12.259 77.908 ;
			RECT	12.395 77.844 12.427 77.908 ;
			RECT	12.563 77.844 12.595 77.908 ;
			RECT	12.731 77.844 12.763 77.908 ;
			RECT	12.899 77.844 12.931 77.908 ;
			RECT	13.067 77.844 13.099 77.908 ;
			RECT	13.235 77.844 13.267 77.908 ;
			RECT	13.403 77.844 13.435 77.908 ;
			RECT	13.571 77.844 13.603 77.908 ;
			RECT	13.739 77.844 13.771 77.908 ;
			RECT	13.907 77.844 13.939 77.908 ;
			RECT	14.075 77.844 14.107 77.908 ;
			RECT	14.243 77.844 14.275 77.908 ;
			RECT	14.411 77.844 14.443 77.908 ;
			RECT	14.579 77.844 14.611 77.908 ;
			RECT	14.747 77.844 14.779 77.908 ;
			RECT	14.915 77.844 14.947 77.908 ;
			RECT	15.083 77.844 15.115 77.908 ;
			RECT	15.251 77.844 15.283 77.908 ;
			RECT	15.419 77.844 15.451 77.908 ;
			RECT	15.587 77.844 15.619 77.908 ;
			RECT	15.755 77.844 15.787 77.908 ;
			RECT	15.923 77.844 15.955 77.908 ;
			RECT	16.091 77.844 16.123 77.908 ;
			RECT	16.259 77.844 16.291 77.908 ;
			RECT	16.427 77.844 16.459 77.908 ;
			RECT	16.595 77.844 16.627 77.908 ;
			RECT	16.763 77.844 16.795 77.908 ;
			RECT	16.931 77.844 16.963 77.908 ;
			RECT	17.099 77.844 17.131 77.908 ;
			RECT	17.267 77.844 17.299 77.908 ;
			RECT	17.435 77.844 17.467 77.908 ;
			RECT	17.603 77.844 17.635 77.908 ;
			RECT	17.771 77.844 17.803 77.908 ;
			RECT	17.939 77.844 17.971 77.908 ;
			RECT	18.107 77.844 18.139 77.908 ;
			RECT	18.275 77.844 18.307 77.908 ;
			RECT	18.443 77.844 18.475 77.908 ;
			RECT	18.611 77.844 18.643 77.908 ;
			RECT	18.779 77.844 18.811 77.908 ;
			RECT	18.947 77.844 18.979 77.908 ;
			RECT	19.115 77.844 19.147 77.908 ;
			RECT	19.283 77.844 19.315 77.908 ;
			RECT	19.451 77.844 19.483 77.908 ;
			RECT	19.619 77.844 19.651 77.908 ;
			RECT	19.787 77.844 19.819 77.908 ;
			RECT	19.955 77.844 19.987 77.908 ;
			RECT	20.123 77.844 20.155 77.908 ;
			RECT	20.291 77.844 20.323 77.908 ;
			RECT	20.459 77.844 20.491 77.908 ;
			RECT	20.627 77.844 20.659 77.908 ;
			RECT	20.795 77.844 20.827 77.908 ;
			RECT	20.963 77.844 20.995 77.908 ;
			RECT	21.131 77.844 21.163 77.908 ;
			RECT	21.299 77.844 21.331 77.908 ;
			RECT	21.467 77.844 21.499 77.908 ;
			RECT	21.635 77.844 21.667 77.908 ;
			RECT	21.803 77.844 21.835 77.908 ;
			RECT	21.971 77.844 22.003 77.908 ;
			RECT	22.139 77.844 22.171 77.908 ;
			RECT	22.307 77.844 22.339 77.908 ;
			RECT	22.475 77.844 22.507 77.908 ;
			RECT	22.643 77.844 22.675 77.908 ;
			RECT	22.811 77.844 22.843 77.908 ;
			RECT	22.979 77.844 23.011 77.908 ;
			RECT	23.147 77.844 23.179 77.908 ;
			RECT	23.315 77.844 23.347 77.908 ;
			RECT	23.483 77.844 23.515 77.908 ;
			RECT	23.651 77.844 23.683 77.908 ;
			RECT	23.819 77.844 23.851 77.908 ;
			RECT	23.987 77.844 24.019 77.908 ;
			RECT	24.155 77.844 24.187 77.908 ;
			RECT	24.323 77.844 24.355 77.908 ;
			RECT	24.491 77.844 24.523 77.908 ;
			RECT	24.659 77.844 24.691 77.908 ;
			RECT	24.827 77.844 24.859 77.908 ;
			RECT	24.995 77.844 25.027 77.908 ;
			RECT	25.163 77.844 25.195 77.908 ;
			RECT	25.331 77.844 25.363 77.908 ;
			RECT	25.499 77.844 25.531 77.908 ;
			RECT	25.667 77.844 25.699 77.908 ;
			RECT	25.835 77.844 25.867 77.908 ;
			RECT	26.003 77.844 26.035 77.908 ;
			RECT	26.171 77.844 26.203 77.908 ;
			RECT	26.339 77.844 26.371 77.908 ;
			RECT	26.507 77.844 26.539 77.908 ;
			RECT	26.675 77.844 26.707 77.908 ;
			RECT	26.843 77.844 26.875 77.908 ;
			RECT	27.011 77.844 27.043 77.908 ;
			RECT	27.179 77.844 27.211 77.908 ;
			RECT	27.347 77.844 27.379 77.908 ;
			RECT	27.515 77.844 27.547 77.908 ;
			RECT	27.683 77.844 27.715 77.908 ;
			RECT	27.851 77.844 27.883 77.908 ;
			RECT	28.019 77.844 28.051 77.908 ;
			RECT	28.187 77.844 28.219 77.908 ;
			RECT	28.355 77.844 28.387 77.908 ;
			RECT	28.523 77.844 28.555 77.908 ;
			RECT	28.691 77.844 28.723 77.908 ;
			RECT	28.859 77.844 28.891 77.908 ;
			RECT	29.027 77.844 29.059 77.908 ;
			RECT	29.195 77.844 29.227 77.908 ;
			RECT	29.363 77.844 29.395 77.908 ;
			RECT	29.531 77.844 29.563 77.908 ;
			RECT	29.699 77.844 29.731 77.908 ;
			RECT	29.867 77.844 29.899 77.908 ;
			RECT	30.035 77.844 30.067 77.908 ;
			RECT	30.203 77.844 30.235 77.908 ;
			RECT	30.371 77.844 30.403 77.908 ;
			RECT	30.539 77.844 30.571 77.908 ;
			RECT	30.707 77.844 30.739 77.908 ;
			RECT	30.875 77.844 30.907 77.908 ;
			RECT	31.043 77.844 31.075 77.908 ;
			RECT	31.211 77.844 31.243 77.908 ;
			RECT	31.379 77.844 31.411 77.908 ;
			RECT	31.547 77.844 31.579 77.908 ;
			RECT	31.715 77.844 31.747 77.908 ;
			RECT	31.883 77.844 31.915 77.908 ;
			RECT	32.051 77.844 32.083 77.908 ;
			RECT	32.219 77.844 32.251 77.908 ;
			RECT	32.387 77.844 32.419 77.908 ;
			RECT	32.555 77.844 32.587 77.908 ;
			RECT	32.723 77.844 32.755 77.908 ;
			RECT	32.891 77.844 32.923 77.908 ;
			RECT	33.059 77.844 33.091 77.908 ;
			RECT	33.227 77.844 33.259 77.908 ;
			RECT	33.395 77.844 33.427 77.908 ;
			RECT	33.563 77.844 33.595 77.908 ;
			RECT	33.731 77.844 33.763 77.908 ;
			RECT	33.899 77.844 33.931 77.908 ;
			RECT	34.067 77.844 34.099 77.908 ;
			RECT	34.235 77.844 34.267 77.908 ;
			RECT	34.403 77.844 34.435 77.908 ;
			RECT	34.571 77.844 34.603 77.908 ;
			RECT	34.739 77.844 34.771 77.908 ;
			RECT	34.907 77.844 34.939 77.908 ;
			RECT	35.075 77.844 35.107 77.908 ;
			RECT	35.243 77.844 35.275 77.908 ;
			RECT	35.411 77.844 35.443 77.908 ;
			RECT	35.579 77.844 35.611 77.908 ;
			RECT	35.747 77.844 35.779 77.908 ;
			RECT	35.915 77.844 35.947 77.908 ;
			RECT	36.083 77.844 36.115 77.908 ;
			RECT	36.251 77.844 36.283 77.908 ;
			RECT	36.419 77.844 36.451 77.908 ;
			RECT	36.587 77.844 36.619 77.908 ;
			RECT	36.755 77.844 36.787 77.908 ;
			RECT	36.923 77.844 36.955 77.908 ;
			RECT	37.091 77.844 37.123 77.908 ;
			RECT	37.259 77.844 37.291 77.908 ;
			RECT	37.427 77.844 37.459 77.908 ;
			RECT	37.595 77.844 37.627 77.908 ;
			RECT	37.763 77.844 37.795 77.908 ;
			RECT	37.931 77.844 37.963 77.908 ;
			RECT	38.099 77.844 38.131 77.908 ;
			RECT	38.267 77.844 38.299 77.908 ;
			RECT	38.435 77.844 38.467 77.908 ;
			RECT	38.603 77.844 38.635 77.908 ;
			RECT	38.771 77.844 38.803 77.908 ;
			RECT	38.939 77.844 38.971 77.908 ;
			RECT	39.107 77.844 39.139 77.908 ;
			RECT	39.275 77.844 39.307 77.908 ;
			RECT	39.443 77.844 39.475 77.908 ;
			RECT	39.611 77.844 39.643 77.908 ;
			RECT	39.779 77.844 39.811 77.908 ;
			RECT	39.947 77.844 39.979 77.908 ;
			RECT	40.115 77.844 40.147 77.908 ;
			RECT	40.283 77.844 40.315 77.908 ;
			RECT	40.451 77.844 40.483 77.908 ;
			RECT	40.619 77.844 40.651 77.908 ;
			RECT	40.787 77.844 40.819 77.908 ;
			RECT	40.955 77.844 40.987 77.908 ;
			RECT	41.123 77.844 41.155 77.908 ;
			RECT	41.291 77.844 41.323 77.908 ;
			RECT	41.459 77.844 41.491 77.908 ;
			RECT	41.627 77.844 41.659 77.908 ;
			RECT	41.795 77.844 41.827 77.908 ;
			RECT	41.963 77.844 41.995 77.908 ;
			RECT	42.131 77.844 42.163 77.908 ;
			RECT	42.299 77.844 42.331 77.908 ;
			RECT	42.467 77.844 42.499 77.908 ;
			RECT	42.635 77.844 42.667 77.908 ;
			RECT	42.803 77.844 42.835 77.908 ;
			RECT	42.971 77.844 43.003 77.908 ;
			RECT	43.139 77.844 43.171 77.908 ;
			RECT	43.307 77.844 43.339 77.908 ;
			RECT	43.475 77.844 43.507 77.908 ;
			RECT	43.643 77.844 43.675 77.908 ;
			RECT	43.811 77.844 43.843 77.908 ;
			RECT	43.979 77.844 44.011 77.908 ;
			RECT	44.147 77.844 44.179 77.908 ;
			RECT	44.315 77.844 44.347 77.908 ;
			RECT	44.483 77.844 44.515 77.908 ;
			RECT	44.651 77.844 44.683 77.908 ;
			RECT	44.819 77.844 44.851 77.908 ;
			RECT	44.987 77.844 45.019 77.908 ;
			RECT	45.155 77.844 45.187 77.908 ;
			RECT	45.323 77.844 45.355 77.908 ;
			RECT	45.491 77.844 45.523 77.908 ;
			RECT	45.659 77.844 45.691 77.908 ;
			RECT	45.827 77.844 45.859 77.908 ;
			RECT	45.995 77.844 46.027 77.908 ;
			RECT	46.163 77.844 46.195 77.908 ;
			RECT	46.331 77.844 46.363 77.908 ;
			RECT	46.499 77.844 46.531 77.908 ;
			RECT	46.667 77.844 46.699 77.908 ;
			RECT	46.835 77.844 46.867 77.908 ;
			RECT	47.003 77.844 47.035 77.908 ;
			RECT	47.171 77.844 47.203 77.908 ;
			RECT	47.339 77.844 47.371 77.908 ;
			RECT	47.507 77.844 47.539 77.908 ;
			RECT	47.675 77.844 47.707 77.908 ;
			RECT	47.843 77.844 47.875 77.908 ;
			RECT	48.011 77.844 48.043 77.908 ;
			RECT	48.179 77.844 48.211 77.908 ;
			RECT	48.347 77.844 48.379 77.908 ;
			RECT	48.515 77.844 48.547 77.908 ;
			RECT	48.683 77.844 48.715 77.908 ;
			RECT	48.851 77.844 48.883 77.908 ;
			RECT	49.019 77.844 49.051 77.908 ;
			RECT	49.187 77.844 49.219 77.908 ;
			RECT	49.318 77.86 49.35 77.892 ;
			RECT	49.439 77.86 49.471 77.892 ;
			RECT	49.569 77.844 49.601 77.908 ;
			RECT	51.881 77.844 51.913 77.908 ;
			RECT	53.132 77.844 53.196 77.908 ;
			RECT	53.812 77.844 53.844 77.908 ;
			RECT	54.251 77.844 54.283 77.908 ;
			RECT	55.562 77.844 55.626 77.908 ;
			RECT	58.603 77.844 58.635 77.908 ;
			RECT	58.733 77.86 58.765 77.892 ;
			RECT	58.854 77.86 58.886 77.892 ;
			RECT	58.985 77.844 59.017 77.908 ;
			RECT	59.153 77.844 59.185 77.908 ;
			RECT	59.321 77.844 59.353 77.908 ;
			RECT	59.489 77.844 59.521 77.908 ;
			RECT	59.657 77.844 59.689 77.908 ;
			RECT	59.825 77.844 59.857 77.908 ;
			RECT	59.993 77.844 60.025 77.908 ;
			RECT	60.161 77.844 60.193 77.908 ;
			RECT	60.329 77.844 60.361 77.908 ;
			RECT	60.497 77.844 60.529 77.908 ;
			RECT	60.665 77.844 60.697 77.908 ;
			RECT	60.833 77.844 60.865 77.908 ;
			RECT	61.001 77.844 61.033 77.908 ;
			RECT	61.169 77.844 61.201 77.908 ;
			RECT	61.337 77.844 61.369 77.908 ;
			RECT	61.505 77.844 61.537 77.908 ;
			RECT	61.673 77.844 61.705 77.908 ;
			RECT	61.841 77.844 61.873 77.908 ;
			RECT	62.009 77.844 62.041 77.908 ;
			RECT	62.177 77.844 62.209 77.908 ;
			RECT	62.345 77.844 62.377 77.908 ;
			RECT	62.513 77.844 62.545 77.908 ;
			RECT	62.681 77.844 62.713 77.908 ;
			RECT	62.849 77.844 62.881 77.908 ;
			RECT	63.017 77.844 63.049 77.908 ;
			RECT	63.185 77.844 63.217 77.908 ;
			RECT	63.353 77.844 63.385 77.908 ;
			RECT	63.521 77.844 63.553 77.908 ;
			RECT	63.689 77.844 63.721 77.908 ;
			RECT	63.857 77.844 63.889 77.908 ;
			RECT	64.025 77.844 64.057 77.908 ;
			RECT	64.193 77.844 64.225 77.908 ;
			RECT	64.361 77.844 64.393 77.908 ;
			RECT	64.529 77.844 64.561 77.908 ;
			RECT	64.697 77.844 64.729 77.908 ;
			RECT	64.865 77.844 64.897 77.908 ;
			RECT	65.033 77.844 65.065 77.908 ;
			RECT	65.201 77.844 65.233 77.908 ;
			RECT	65.369 77.844 65.401 77.908 ;
			RECT	65.537 77.844 65.569 77.908 ;
			RECT	65.705 77.844 65.737 77.908 ;
			RECT	65.873 77.844 65.905 77.908 ;
			RECT	66.041 77.844 66.073 77.908 ;
			RECT	66.209 77.844 66.241 77.908 ;
			RECT	66.377 77.844 66.409 77.908 ;
			RECT	66.545 77.844 66.577 77.908 ;
			RECT	66.713 77.844 66.745 77.908 ;
			RECT	66.881 77.844 66.913 77.908 ;
			RECT	67.049 77.844 67.081 77.908 ;
			RECT	67.217 77.844 67.249 77.908 ;
			RECT	67.385 77.844 67.417 77.908 ;
			RECT	67.553 77.844 67.585 77.908 ;
			RECT	67.721 77.844 67.753 77.908 ;
			RECT	67.889 77.844 67.921 77.908 ;
			RECT	68.057 77.844 68.089 77.908 ;
			RECT	68.225 77.844 68.257 77.908 ;
			RECT	68.393 77.844 68.425 77.908 ;
			RECT	68.561 77.844 68.593 77.908 ;
			RECT	68.729 77.844 68.761 77.908 ;
			RECT	68.897 77.844 68.929 77.908 ;
			RECT	69.065 77.844 69.097 77.908 ;
			RECT	69.233 77.844 69.265 77.908 ;
			RECT	69.401 77.844 69.433 77.908 ;
			RECT	69.569 77.844 69.601 77.908 ;
			RECT	69.737 77.844 69.769 77.908 ;
			RECT	69.905 77.844 69.937 77.908 ;
			RECT	70.073 77.844 70.105 77.908 ;
			RECT	70.241 77.844 70.273 77.908 ;
			RECT	70.409 77.844 70.441 77.908 ;
			RECT	70.577 77.844 70.609 77.908 ;
			RECT	70.745 77.844 70.777 77.908 ;
			RECT	70.913 77.844 70.945 77.908 ;
			RECT	71.081 77.844 71.113 77.908 ;
			RECT	71.249 77.844 71.281 77.908 ;
			RECT	71.417 77.844 71.449 77.908 ;
			RECT	71.585 77.844 71.617 77.908 ;
			RECT	71.753 77.844 71.785 77.908 ;
			RECT	71.921 77.844 71.953 77.908 ;
			RECT	72.089 77.844 72.121 77.908 ;
			RECT	72.257 77.844 72.289 77.908 ;
			RECT	72.425 77.844 72.457 77.908 ;
			RECT	72.593 77.844 72.625 77.908 ;
			RECT	72.761 77.844 72.793 77.908 ;
			RECT	72.929 77.844 72.961 77.908 ;
			RECT	73.097 77.844 73.129 77.908 ;
			RECT	73.265 77.844 73.297 77.908 ;
			RECT	73.433 77.844 73.465 77.908 ;
			RECT	73.601 77.844 73.633 77.908 ;
			RECT	73.769 77.844 73.801 77.908 ;
			RECT	73.937 77.844 73.969 77.908 ;
			RECT	74.105 77.844 74.137 77.908 ;
			RECT	74.273 77.844 74.305 77.908 ;
			RECT	74.441 77.844 74.473 77.908 ;
			RECT	74.609 77.844 74.641 77.908 ;
			RECT	74.777 77.844 74.809 77.908 ;
			RECT	74.945 77.844 74.977 77.908 ;
			RECT	75.113 77.844 75.145 77.908 ;
			RECT	75.281 77.844 75.313 77.908 ;
			RECT	75.449 77.844 75.481 77.908 ;
			RECT	75.617 77.844 75.649 77.908 ;
			RECT	75.785 77.844 75.817 77.908 ;
			RECT	75.953 77.844 75.985 77.908 ;
			RECT	76.121 77.844 76.153 77.908 ;
			RECT	76.289 77.844 76.321 77.908 ;
			RECT	76.457 77.844 76.489 77.908 ;
			RECT	76.625 77.844 76.657 77.908 ;
			RECT	76.793 77.844 76.825 77.908 ;
			RECT	76.961 77.844 76.993 77.908 ;
			RECT	77.129 77.844 77.161 77.908 ;
			RECT	77.297 77.844 77.329 77.908 ;
			RECT	77.465 77.844 77.497 77.908 ;
			RECT	77.633 77.844 77.665 77.908 ;
			RECT	77.801 77.844 77.833 77.908 ;
			RECT	77.969 77.844 78.001 77.908 ;
			RECT	78.137 77.844 78.169 77.908 ;
			RECT	78.305 77.844 78.337 77.908 ;
			RECT	78.473 77.844 78.505 77.908 ;
			RECT	78.641 77.844 78.673 77.908 ;
			RECT	78.809 77.844 78.841 77.908 ;
			RECT	78.977 77.844 79.009 77.908 ;
			RECT	79.145 77.844 79.177 77.908 ;
			RECT	79.313 77.844 79.345 77.908 ;
			RECT	79.481 77.844 79.513 77.908 ;
			RECT	79.649 77.844 79.681 77.908 ;
			RECT	79.817 77.844 79.849 77.908 ;
			RECT	79.985 77.844 80.017 77.908 ;
			RECT	80.153 77.844 80.185 77.908 ;
			RECT	80.321 77.844 80.353 77.908 ;
			RECT	80.489 77.844 80.521 77.908 ;
			RECT	80.657 77.844 80.689 77.908 ;
			RECT	80.825 77.844 80.857 77.908 ;
			RECT	80.993 77.844 81.025 77.908 ;
			RECT	81.161 77.844 81.193 77.908 ;
			RECT	81.329 77.844 81.361 77.908 ;
			RECT	81.497 77.844 81.529 77.908 ;
			RECT	81.665 77.844 81.697 77.908 ;
			RECT	81.833 77.844 81.865 77.908 ;
			RECT	82.001 77.844 82.033 77.908 ;
			RECT	82.169 77.844 82.201 77.908 ;
			RECT	82.337 77.844 82.369 77.908 ;
			RECT	82.505 77.844 82.537 77.908 ;
			RECT	82.673 77.844 82.705 77.908 ;
			RECT	82.841 77.844 82.873 77.908 ;
			RECT	83.009 77.844 83.041 77.908 ;
			RECT	83.177 77.844 83.209 77.908 ;
			RECT	83.345 77.844 83.377 77.908 ;
			RECT	83.513 77.844 83.545 77.908 ;
			RECT	83.681 77.844 83.713 77.908 ;
			RECT	83.849 77.844 83.881 77.908 ;
			RECT	84.017 77.844 84.049 77.908 ;
			RECT	84.185 77.844 84.217 77.908 ;
			RECT	84.353 77.844 84.385 77.908 ;
			RECT	84.521 77.844 84.553 77.908 ;
			RECT	84.689 77.844 84.721 77.908 ;
			RECT	84.857 77.844 84.889 77.908 ;
			RECT	85.025 77.844 85.057 77.908 ;
			RECT	85.193 77.844 85.225 77.908 ;
			RECT	85.361 77.844 85.393 77.908 ;
			RECT	85.529 77.844 85.561 77.908 ;
			RECT	85.697 77.844 85.729 77.908 ;
			RECT	85.865 77.844 85.897 77.908 ;
			RECT	86.033 77.844 86.065 77.908 ;
			RECT	86.201 77.844 86.233 77.908 ;
			RECT	86.369 77.844 86.401 77.908 ;
			RECT	86.537 77.844 86.569 77.908 ;
			RECT	86.705 77.844 86.737 77.908 ;
			RECT	86.873 77.844 86.905 77.908 ;
			RECT	87.041 77.844 87.073 77.908 ;
			RECT	87.209 77.844 87.241 77.908 ;
			RECT	87.377 77.844 87.409 77.908 ;
			RECT	87.545 77.844 87.577 77.908 ;
			RECT	87.713 77.844 87.745 77.908 ;
			RECT	87.881 77.844 87.913 77.908 ;
			RECT	88.049 77.844 88.081 77.908 ;
			RECT	88.217 77.844 88.249 77.908 ;
			RECT	88.385 77.844 88.417 77.908 ;
			RECT	88.553 77.844 88.585 77.908 ;
			RECT	88.721 77.844 88.753 77.908 ;
			RECT	88.889 77.844 88.921 77.908 ;
			RECT	89.057 77.844 89.089 77.908 ;
			RECT	89.225 77.844 89.257 77.908 ;
			RECT	89.393 77.844 89.425 77.908 ;
			RECT	89.561 77.844 89.593 77.908 ;
			RECT	89.729 77.844 89.761 77.908 ;
			RECT	89.897 77.844 89.929 77.908 ;
			RECT	90.065 77.844 90.097 77.908 ;
			RECT	90.233 77.844 90.265 77.908 ;
			RECT	90.401 77.844 90.433 77.908 ;
			RECT	90.569 77.844 90.601 77.908 ;
			RECT	90.737 77.844 90.769 77.908 ;
			RECT	90.905 77.844 90.937 77.908 ;
			RECT	91.073 77.844 91.105 77.908 ;
			RECT	91.241 77.844 91.273 77.908 ;
			RECT	91.409 77.844 91.441 77.908 ;
			RECT	91.577 77.844 91.609 77.908 ;
			RECT	91.745 77.844 91.777 77.908 ;
			RECT	91.913 77.844 91.945 77.908 ;
			RECT	92.081 77.844 92.113 77.908 ;
			RECT	92.249 77.844 92.281 77.908 ;
			RECT	92.417 77.844 92.449 77.908 ;
			RECT	92.585 77.844 92.617 77.908 ;
			RECT	92.753 77.844 92.785 77.908 ;
			RECT	92.921 77.844 92.953 77.908 ;
			RECT	93.089 77.844 93.121 77.908 ;
			RECT	93.257 77.844 93.289 77.908 ;
			RECT	93.425 77.844 93.457 77.908 ;
			RECT	93.593 77.844 93.625 77.908 ;
			RECT	93.761 77.844 93.793 77.908 ;
			RECT	93.929 77.844 93.961 77.908 ;
			RECT	94.097 77.844 94.129 77.908 ;
			RECT	94.265 77.844 94.297 77.908 ;
			RECT	94.433 77.844 94.465 77.908 ;
			RECT	94.601 77.844 94.633 77.908 ;
			RECT	94.769 77.844 94.801 77.908 ;
			RECT	94.937 77.844 94.969 77.908 ;
			RECT	95.105 77.844 95.137 77.908 ;
			RECT	95.273 77.844 95.305 77.908 ;
			RECT	95.441 77.844 95.473 77.908 ;
			RECT	95.609 77.844 95.641 77.908 ;
			RECT	95.777 77.844 95.809 77.908 ;
			RECT	95.945 77.844 95.977 77.908 ;
			RECT	96.113 77.844 96.145 77.908 ;
			RECT	96.281 77.844 96.313 77.908 ;
			RECT	96.449 77.844 96.481 77.908 ;
			RECT	96.617 77.844 96.649 77.908 ;
			RECT	96.785 77.844 96.817 77.908 ;
			RECT	96.953 77.844 96.985 77.908 ;
			RECT	97.121 77.844 97.153 77.908 ;
			RECT	97.289 77.844 97.321 77.908 ;
			RECT	97.457 77.844 97.489 77.908 ;
			RECT	97.625 77.844 97.657 77.908 ;
			RECT	97.793 77.844 97.825 77.908 ;
			RECT	97.961 77.844 97.993 77.908 ;
			RECT	98.129 77.844 98.161 77.908 ;
			RECT	98.297 77.844 98.329 77.908 ;
			RECT	98.465 77.844 98.497 77.908 ;
			RECT	98.633 77.844 98.665 77.908 ;
			RECT	98.801 77.844 98.833 77.908 ;
			RECT	98.969 77.844 99.001 77.908 ;
			RECT	99.137 77.844 99.169 77.908 ;
			RECT	99.305 77.844 99.337 77.908 ;
			RECT	99.473 77.844 99.505 77.908 ;
			RECT	99.641 77.844 99.673 77.908 ;
			RECT	99.809 77.844 99.841 77.908 ;
			RECT	99.977 77.844 100.009 77.908 ;
			RECT	100.145 77.844 100.177 77.908 ;
			RECT	100.313 77.844 100.345 77.908 ;
			RECT	100.481 77.844 100.513 77.908 ;
			RECT	100.649 77.844 100.681 77.908 ;
			RECT	100.817 77.844 100.849 77.908 ;
			RECT	100.985 77.844 101.017 77.908 ;
			RECT	101.153 77.844 101.185 77.908 ;
			RECT	101.321 77.844 101.353 77.908 ;
			RECT	101.489 77.844 101.521 77.908 ;
			RECT	101.657 77.844 101.689 77.908 ;
			RECT	101.825 77.844 101.857 77.908 ;
			RECT	101.993 77.844 102.025 77.908 ;
			RECT	102.123 77.86 102.155 77.892 ;
			RECT	102.245 77.855 102.277 77.887 ;
			RECT	102.375 77.844 102.407 77.908 ;
			RECT	103.795 77.844 103.827 77.908 ;
			RECT	103.925 77.855 103.957 77.887 ;
			RECT	104.047 77.86 104.079 77.892 ;
			RECT	104.177 77.844 104.209 77.908 ;
			RECT	104.345 77.844 104.377 77.908 ;
			RECT	104.513 77.844 104.545 77.908 ;
			RECT	104.681 77.844 104.713 77.908 ;
			RECT	104.849 77.844 104.881 77.908 ;
			RECT	105.017 77.844 105.049 77.908 ;
			RECT	105.185 77.844 105.217 77.908 ;
			RECT	105.353 77.844 105.385 77.908 ;
			RECT	105.521 77.844 105.553 77.908 ;
			RECT	105.689 77.844 105.721 77.908 ;
			RECT	105.857 77.844 105.889 77.908 ;
			RECT	106.025 77.844 106.057 77.908 ;
			RECT	106.193 77.844 106.225 77.908 ;
			RECT	106.361 77.844 106.393 77.908 ;
			RECT	106.529 77.844 106.561 77.908 ;
			RECT	106.697 77.844 106.729 77.908 ;
			RECT	106.865 77.844 106.897 77.908 ;
			RECT	107.033 77.844 107.065 77.908 ;
			RECT	107.201 77.844 107.233 77.908 ;
			RECT	107.369 77.844 107.401 77.908 ;
			RECT	107.537 77.844 107.569 77.908 ;
			RECT	107.705 77.844 107.737 77.908 ;
			RECT	107.873 77.844 107.905 77.908 ;
			RECT	108.041 77.844 108.073 77.908 ;
			RECT	108.209 77.844 108.241 77.908 ;
			RECT	108.377 77.844 108.409 77.908 ;
			RECT	108.545 77.844 108.577 77.908 ;
			RECT	108.713 77.844 108.745 77.908 ;
			RECT	108.881 77.844 108.913 77.908 ;
			RECT	109.049 77.844 109.081 77.908 ;
			RECT	109.217 77.844 109.249 77.908 ;
			RECT	109.385 77.844 109.417 77.908 ;
			RECT	109.553 77.844 109.585 77.908 ;
			RECT	109.721 77.844 109.753 77.908 ;
			RECT	109.889 77.844 109.921 77.908 ;
			RECT	110.057 77.844 110.089 77.908 ;
			RECT	110.225 77.844 110.257 77.908 ;
			RECT	110.393 77.844 110.425 77.908 ;
			RECT	110.561 77.844 110.593 77.908 ;
			RECT	110.729 77.844 110.761 77.908 ;
			RECT	110.897 77.844 110.929 77.908 ;
			RECT	111.065 77.844 111.097 77.908 ;
			RECT	111.233 77.844 111.265 77.908 ;
			RECT	111.401 77.844 111.433 77.908 ;
			RECT	111.569 77.844 111.601 77.908 ;
			RECT	111.737 77.844 111.769 77.908 ;
			RECT	111.905 77.844 111.937 77.908 ;
			RECT	112.073 77.844 112.105 77.908 ;
			RECT	112.241 77.844 112.273 77.908 ;
			RECT	112.409 77.844 112.441 77.908 ;
			RECT	112.577 77.844 112.609 77.908 ;
			RECT	112.745 77.844 112.777 77.908 ;
			RECT	112.913 77.844 112.945 77.908 ;
			RECT	113.081 77.844 113.113 77.908 ;
			RECT	113.249 77.844 113.281 77.908 ;
			RECT	113.417 77.844 113.449 77.908 ;
			RECT	113.585 77.844 113.617 77.908 ;
			RECT	113.753 77.844 113.785 77.908 ;
			RECT	113.921 77.844 113.953 77.908 ;
			RECT	114.089 77.844 114.121 77.908 ;
			RECT	114.257 77.844 114.289 77.908 ;
			RECT	114.425 77.844 114.457 77.908 ;
			RECT	114.593 77.844 114.625 77.908 ;
			RECT	114.761 77.844 114.793 77.908 ;
			RECT	114.929 77.844 114.961 77.908 ;
			RECT	115.097 77.844 115.129 77.908 ;
			RECT	115.265 77.844 115.297 77.908 ;
			RECT	115.433 77.844 115.465 77.908 ;
			RECT	115.601 77.844 115.633 77.908 ;
			RECT	115.769 77.844 115.801 77.908 ;
			RECT	115.937 77.844 115.969 77.908 ;
			RECT	116.105 77.844 116.137 77.908 ;
			RECT	116.273 77.844 116.305 77.908 ;
			RECT	116.441 77.844 116.473 77.908 ;
			RECT	116.609 77.844 116.641 77.908 ;
			RECT	116.777 77.844 116.809 77.908 ;
			RECT	116.945 77.844 116.977 77.908 ;
			RECT	117.113 77.844 117.145 77.908 ;
			RECT	117.281 77.844 117.313 77.908 ;
			RECT	117.449 77.844 117.481 77.908 ;
			RECT	117.617 77.844 117.649 77.908 ;
			RECT	117.785 77.844 117.817 77.908 ;
			RECT	117.953 77.844 117.985 77.908 ;
			RECT	118.121 77.844 118.153 77.908 ;
			RECT	118.289 77.844 118.321 77.908 ;
			RECT	118.457 77.844 118.489 77.908 ;
			RECT	118.625 77.844 118.657 77.908 ;
			RECT	118.793 77.844 118.825 77.908 ;
			RECT	118.961 77.844 118.993 77.908 ;
			RECT	119.129 77.844 119.161 77.908 ;
			RECT	119.297 77.844 119.329 77.908 ;
			RECT	119.465 77.844 119.497 77.908 ;
			RECT	119.633 77.844 119.665 77.908 ;
			RECT	119.801 77.844 119.833 77.908 ;
			RECT	119.969 77.844 120.001 77.908 ;
			RECT	120.137 77.844 120.169 77.908 ;
			RECT	120.305 77.844 120.337 77.908 ;
			RECT	120.473 77.844 120.505 77.908 ;
			RECT	120.641 77.844 120.673 77.908 ;
			RECT	120.809 77.844 120.841 77.908 ;
			RECT	120.977 77.844 121.009 77.908 ;
			RECT	121.145 77.844 121.177 77.908 ;
			RECT	121.313 77.844 121.345 77.908 ;
			RECT	121.481 77.844 121.513 77.908 ;
			RECT	121.649 77.844 121.681 77.908 ;
			RECT	121.817 77.844 121.849 77.908 ;
			RECT	121.985 77.844 122.017 77.908 ;
			RECT	122.153 77.844 122.185 77.908 ;
			RECT	122.321 77.844 122.353 77.908 ;
			RECT	122.489 77.844 122.521 77.908 ;
			RECT	122.657 77.844 122.689 77.908 ;
			RECT	122.825 77.844 122.857 77.908 ;
			RECT	122.993 77.844 123.025 77.908 ;
			RECT	123.161 77.844 123.193 77.908 ;
			RECT	123.329 77.844 123.361 77.908 ;
			RECT	123.497 77.844 123.529 77.908 ;
			RECT	123.665 77.844 123.697 77.908 ;
			RECT	123.833 77.844 123.865 77.908 ;
			RECT	124.001 77.844 124.033 77.908 ;
			RECT	124.169 77.844 124.201 77.908 ;
			RECT	124.337 77.844 124.369 77.908 ;
			RECT	124.505 77.844 124.537 77.908 ;
			RECT	124.673 77.844 124.705 77.908 ;
			RECT	124.841 77.844 124.873 77.908 ;
			RECT	125.009 77.844 125.041 77.908 ;
			RECT	125.177 77.844 125.209 77.908 ;
			RECT	125.345 77.844 125.377 77.908 ;
			RECT	125.513 77.844 125.545 77.908 ;
			RECT	125.681 77.844 125.713 77.908 ;
			RECT	125.849 77.844 125.881 77.908 ;
			RECT	126.017 77.844 126.049 77.908 ;
			RECT	126.185 77.844 126.217 77.908 ;
			RECT	126.353 77.844 126.385 77.908 ;
			RECT	126.521 77.844 126.553 77.908 ;
			RECT	126.689 77.844 126.721 77.908 ;
			RECT	126.857 77.844 126.889 77.908 ;
			RECT	127.025 77.844 127.057 77.908 ;
			RECT	127.193 77.844 127.225 77.908 ;
			RECT	127.361 77.844 127.393 77.908 ;
			RECT	127.529 77.844 127.561 77.908 ;
			RECT	127.697 77.844 127.729 77.908 ;
			RECT	127.865 77.844 127.897 77.908 ;
			RECT	128.033 77.844 128.065 77.908 ;
			RECT	128.201 77.844 128.233 77.908 ;
			RECT	128.369 77.844 128.401 77.908 ;
			RECT	128.537 77.844 128.569 77.908 ;
			RECT	128.705 77.844 128.737 77.908 ;
			RECT	128.873 77.844 128.905 77.908 ;
			RECT	129.041 77.844 129.073 77.908 ;
			RECT	129.209 77.844 129.241 77.908 ;
			RECT	129.377 77.844 129.409 77.908 ;
			RECT	129.545 77.844 129.577 77.908 ;
			RECT	129.713 77.844 129.745 77.908 ;
			RECT	129.881 77.844 129.913 77.908 ;
			RECT	130.049 77.844 130.081 77.908 ;
			RECT	130.217 77.844 130.249 77.908 ;
			RECT	130.385 77.844 130.417 77.908 ;
			RECT	130.553 77.844 130.585 77.908 ;
			RECT	130.721 77.844 130.753 77.908 ;
			RECT	130.889 77.844 130.921 77.908 ;
			RECT	131.057 77.844 131.089 77.908 ;
			RECT	131.225 77.844 131.257 77.908 ;
			RECT	131.393 77.844 131.425 77.908 ;
			RECT	131.561 77.844 131.593 77.908 ;
			RECT	131.729 77.844 131.761 77.908 ;
			RECT	131.897 77.844 131.929 77.908 ;
			RECT	132.065 77.844 132.097 77.908 ;
			RECT	132.233 77.844 132.265 77.908 ;
			RECT	132.401 77.844 132.433 77.908 ;
			RECT	132.569 77.844 132.601 77.908 ;
			RECT	132.737 77.844 132.769 77.908 ;
			RECT	132.905 77.844 132.937 77.908 ;
			RECT	133.073 77.844 133.105 77.908 ;
			RECT	133.241 77.844 133.273 77.908 ;
			RECT	133.409 77.844 133.441 77.908 ;
			RECT	133.577 77.844 133.609 77.908 ;
			RECT	133.745 77.844 133.777 77.908 ;
			RECT	133.913 77.844 133.945 77.908 ;
			RECT	134.081 77.844 134.113 77.908 ;
			RECT	134.249 77.844 134.281 77.908 ;
			RECT	134.417 77.844 134.449 77.908 ;
			RECT	134.585 77.844 134.617 77.908 ;
			RECT	134.753 77.844 134.785 77.908 ;
			RECT	134.921 77.844 134.953 77.908 ;
			RECT	135.089 77.844 135.121 77.908 ;
			RECT	135.257 77.844 135.289 77.908 ;
			RECT	135.425 77.844 135.457 77.908 ;
			RECT	135.593 77.844 135.625 77.908 ;
			RECT	135.761 77.844 135.793 77.908 ;
			RECT	135.929 77.844 135.961 77.908 ;
			RECT	136.097 77.844 136.129 77.908 ;
			RECT	136.265 77.844 136.297 77.908 ;
			RECT	136.433 77.844 136.465 77.908 ;
			RECT	136.601 77.844 136.633 77.908 ;
			RECT	136.769 77.844 136.801 77.908 ;
			RECT	136.937 77.844 136.969 77.908 ;
			RECT	137.105 77.844 137.137 77.908 ;
			RECT	137.273 77.844 137.305 77.908 ;
			RECT	137.441 77.844 137.473 77.908 ;
			RECT	137.609 77.844 137.641 77.908 ;
			RECT	137.777 77.844 137.809 77.908 ;
			RECT	137.945 77.844 137.977 77.908 ;
			RECT	138.113 77.844 138.145 77.908 ;
			RECT	138.281 77.844 138.313 77.908 ;
			RECT	138.449 77.844 138.481 77.908 ;
			RECT	138.617 77.844 138.649 77.908 ;
			RECT	138.785 77.844 138.817 77.908 ;
			RECT	138.953 77.844 138.985 77.908 ;
			RECT	139.121 77.844 139.153 77.908 ;
			RECT	139.289 77.844 139.321 77.908 ;
			RECT	139.457 77.844 139.489 77.908 ;
			RECT	139.625 77.844 139.657 77.908 ;
			RECT	139.793 77.844 139.825 77.908 ;
			RECT	139.961 77.844 139.993 77.908 ;
			RECT	140.129 77.844 140.161 77.908 ;
			RECT	140.297 77.844 140.329 77.908 ;
			RECT	140.465 77.844 140.497 77.908 ;
			RECT	140.633 77.844 140.665 77.908 ;
			RECT	140.801 77.844 140.833 77.908 ;
			RECT	140.969 77.844 141.001 77.908 ;
			RECT	141.137 77.844 141.169 77.908 ;
			RECT	141.305 77.844 141.337 77.908 ;
			RECT	141.473 77.844 141.505 77.908 ;
			RECT	141.641 77.844 141.673 77.908 ;
			RECT	141.809 77.844 141.841 77.908 ;
			RECT	141.977 77.844 142.009 77.908 ;
			RECT	142.145 77.844 142.177 77.908 ;
			RECT	142.313 77.844 142.345 77.908 ;
			RECT	142.481 77.844 142.513 77.908 ;
			RECT	142.649 77.844 142.681 77.908 ;
			RECT	142.817 77.844 142.849 77.908 ;
			RECT	142.985 77.844 143.017 77.908 ;
			RECT	143.153 77.844 143.185 77.908 ;
			RECT	143.321 77.844 143.353 77.908 ;
			RECT	143.489 77.844 143.521 77.908 ;
			RECT	143.657 77.844 143.689 77.908 ;
			RECT	143.825 77.844 143.857 77.908 ;
			RECT	143.993 77.844 144.025 77.908 ;
			RECT	144.161 77.844 144.193 77.908 ;
			RECT	144.329 77.844 144.361 77.908 ;
			RECT	144.497 77.844 144.529 77.908 ;
			RECT	144.665 77.844 144.697 77.908 ;
			RECT	144.833 77.844 144.865 77.908 ;
			RECT	145.001 77.844 145.033 77.908 ;
			RECT	145.169 77.844 145.201 77.908 ;
			RECT	145.337 77.844 145.369 77.908 ;
			RECT	145.505 77.844 145.537 77.908 ;
			RECT	145.673 77.844 145.705 77.908 ;
			RECT	145.841 77.844 145.873 77.908 ;
			RECT	146.009 77.844 146.041 77.908 ;
			RECT	146.177 77.844 146.209 77.908 ;
			RECT	146.345 77.844 146.377 77.908 ;
			RECT	146.513 77.844 146.545 77.908 ;
			RECT	146.681 77.844 146.713 77.908 ;
			RECT	146.849 77.844 146.881 77.908 ;
			RECT	147.017 77.844 147.049 77.908 ;
			RECT	147.185 77.844 147.217 77.908 ;
			RECT	147.316 77.86 147.348 77.892 ;
			RECT	147.437 77.86 147.469 77.892 ;
			RECT	147.567 77.844 147.599 77.908 ;
			RECT	149.879 77.844 149.911 77.908 ;
			RECT	151.13 77.844 151.194 77.908 ;
			RECT	151.81 77.844 151.842 77.908 ;
			RECT	152.249 77.844 152.281 77.908 ;
			RECT	153.56 77.844 153.624 77.908 ;
			RECT	156.601 77.844 156.633 77.908 ;
			RECT	156.731 77.86 156.763 77.892 ;
			RECT	156.852 77.86 156.884 77.892 ;
			RECT	156.983 77.844 157.015 77.908 ;
			RECT	157.151 77.844 157.183 77.908 ;
			RECT	157.319 77.844 157.351 77.908 ;
			RECT	157.487 77.844 157.519 77.908 ;
			RECT	157.655 77.844 157.687 77.908 ;
			RECT	157.823 77.844 157.855 77.908 ;
			RECT	157.991 77.844 158.023 77.908 ;
			RECT	158.159 77.844 158.191 77.908 ;
			RECT	158.327 77.844 158.359 77.908 ;
			RECT	158.495 77.844 158.527 77.908 ;
			RECT	158.663 77.844 158.695 77.908 ;
			RECT	158.831 77.844 158.863 77.908 ;
			RECT	158.999 77.844 159.031 77.908 ;
			RECT	159.167 77.844 159.199 77.908 ;
			RECT	159.335 77.844 159.367 77.908 ;
			RECT	159.503 77.844 159.535 77.908 ;
			RECT	159.671 77.844 159.703 77.908 ;
			RECT	159.839 77.844 159.871 77.908 ;
			RECT	160.007 77.844 160.039 77.908 ;
			RECT	160.175 77.844 160.207 77.908 ;
			RECT	160.343 77.844 160.375 77.908 ;
			RECT	160.511 77.844 160.543 77.908 ;
			RECT	160.679 77.844 160.711 77.908 ;
			RECT	160.847 77.844 160.879 77.908 ;
			RECT	161.015 77.844 161.047 77.908 ;
			RECT	161.183 77.844 161.215 77.908 ;
			RECT	161.351 77.844 161.383 77.908 ;
			RECT	161.519 77.844 161.551 77.908 ;
			RECT	161.687 77.844 161.719 77.908 ;
			RECT	161.855 77.844 161.887 77.908 ;
			RECT	162.023 77.844 162.055 77.908 ;
			RECT	162.191 77.844 162.223 77.908 ;
			RECT	162.359 77.844 162.391 77.908 ;
			RECT	162.527 77.844 162.559 77.908 ;
			RECT	162.695 77.844 162.727 77.908 ;
			RECT	162.863 77.844 162.895 77.908 ;
			RECT	163.031 77.844 163.063 77.908 ;
			RECT	163.199 77.844 163.231 77.908 ;
			RECT	163.367 77.844 163.399 77.908 ;
			RECT	163.535 77.844 163.567 77.908 ;
			RECT	163.703 77.844 163.735 77.908 ;
			RECT	163.871 77.844 163.903 77.908 ;
			RECT	164.039 77.844 164.071 77.908 ;
			RECT	164.207 77.844 164.239 77.908 ;
			RECT	164.375 77.844 164.407 77.908 ;
			RECT	164.543 77.844 164.575 77.908 ;
			RECT	164.711 77.844 164.743 77.908 ;
			RECT	164.879 77.844 164.911 77.908 ;
			RECT	165.047 77.844 165.079 77.908 ;
			RECT	165.215 77.844 165.247 77.908 ;
			RECT	165.383 77.844 165.415 77.908 ;
			RECT	165.551 77.844 165.583 77.908 ;
			RECT	165.719 77.844 165.751 77.908 ;
			RECT	165.887 77.844 165.919 77.908 ;
			RECT	166.055 77.844 166.087 77.908 ;
			RECT	166.223 77.844 166.255 77.908 ;
			RECT	166.391 77.844 166.423 77.908 ;
			RECT	166.559 77.844 166.591 77.908 ;
			RECT	166.727 77.844 166.759 77.908 ;
			RECT	166.895 77.844 166.927 77.908 ;
			RECT	167.063 77.844 167.095 77.908 ;
			RECT	167.231 77.844 167.263 77.908 ;
			RECT	167.399 77.844 167.431 77.908 ;
			RECT	167.567 77.844 167.599 77.908 ;
			RECT	167.735 77.844 167.767 77.908 ;
			RECT	167.903 77.844 167.935 77.908 ;
			RECT	168.071 77.844 168.103 77.908 ;
			RECT	168.239 77.844 168.271 77.908 ;
			RECT	168.407 77.844 168.439 77.908 ;
			RECT	168.575 77.844 168.607 77.908 ;
			RECT	168.743 77.844 168.775 77.908 ;
			RECT	168.911 77.844 168.943 77.908 ;
			RECT	169.079 77.844 169.111 77.908 ;
			RECT	169.247 77.844 169.279 77.908 ;
			RECT	169.415 77.844 169.447 77.908 ;
			RECT	169.583 77.844 169.615 77.908 ;
			RECT	169.751 77.844 169.783 77.908 ;
			RECT	169.919 77.844 169.951 77.908 ;
			RECT	170.087 77.844 170.119 77.908 ;
			RECT	170.255 77.844 170.287 77.908 ;
			RECT	170.423 77.844 170.455 77.908 ;
			RECT	170.591 77.844 170.623 77.908 ;
			RECT	170.759 77.844 170.791 77.908 ;
			RECT	170.927 77.844 170.959 77.908 ;
			RECT	171.095 77.844 171.127 77.908 ;
			RECT	171.263 77.844 171.295 77.908 ;
			RECT	171.431 77.844 171.463 77.908 ;
			RECT	171.599 77.844 171.631 77.908 ;
			RECT	171.767 77.844 171.799 77.908 ;
			RECT	171.935 77.844 171.967 77.908 ;
			RECT	172.103 77.844 172.135 77.908 ;
			RECT	172.271 77.844 172.303 77.908 ;
			RECT	172.439 77.844 172.471 77.908 ;
			RECT	172.607 77.844 172.639 77.908 ;
			RECT	172.775 77.844 172.807 77.908 ;
			RECT	172.943 77.844 172.975 77.908 ;
			RECT	173.111 77.844 173.143 77.908 ;
			RECT	173.279 77.844 173.311 77.908 ;
			RECT	173.447 77.844 173.479 77.908 ;
			RECT	173.615 77.844 173.647 77.908 ;
			RECT	173.783 77.844 173.815 77.908 ;
			RECT	173.951 77.844 173.983 77.908 ;
			RECT	174.119 77.844 174.151 77.908 ;
			RECT	174.287 77.844 174.319 77.908 ;
			RECT	174.455 77.844 174.487 77.908 ;
			RECT	174.623 77.844 174.655 77.908 ;
			RECT	174.791 77.844 174.823 77.908 ;
			RECT	174.959 77.844 174.991 77.908 ;
			RECT	175.127 77.844 175.159 77.908 ;
			RECT	175.295 77.844 175.327 77.908 ;
			RECT	175.463 77.844 175.495 77.908 ;
			RECT	175.631 77.844 175.663 77.908 ;
			RECT	175.799 77.844 175.831 77.908 ;
			RECT	175.967 77.844 175.999 77.908 ;
			RECT	176.135 77.844 176.167 77.908 ;
			RECT	176.303 77.844 176.335 77.908 ;
			RECT	176.471 77.844 176.503 77.908 ;
			RECT	176.639 77.844 176.671 77.908 ;
			RECT	176.807 77.844 176.839 77.908 ;
			RECT	176.975 77.844 177.007 77.908 ;
			RECT	177.143 77.844 177.175 77.908 ;
			RECT	177.311 77.844 177.343 77.908 ;
			RECT	177.479 77.844 177.511 77.908 ;
			RECT	177.647 77.844 177.679 77.908 ;
			RECT	177.815 77.844 177.847 77.908 ;
			RECT	177.983 77.844 178.015 77.908 ;
			RECT	178.151 77.844 178.183 77.908 ;
			RECT	178.319 77.844 178.351 77.908 ;
			RECT	178.487 77.844 178.519 77.908 ;
			RECT	178.655 77.844 178.687 77.908 ;
			RECT	178.823 77.844 178.855 77.908 ;
			RECT	178.991 77.844 179.023 77.908 ;
			RECT	179.159 77.844 179.191 77.908 ;
			RECT	179.327 77.844 179.359 77.908 ;
			RECT	179.495 77.844 179.527 77.908 ;
			RECT	179.663 77.844 179.695 77.908 ;
			RECT	179.831 77.844 179.863 77.908 ;
			RECT	179.999 77.844 180.031 77.908 ;
			RECT	180.167 77.844 180.199 77.908 ;
			RECT	180.335 77.844 180.367 77.908 ;
			RECT	180.503 77.844 180.535 77.908 ;
			RECT	180.671 77.844 180.703 77.908 ;
			RECT	180.839 77.844 180.871 77.908 ;
			RECT	181.007 77.844 181.039 77.908 ;
			RECT	181.175 77.844 181.207 77.908 ;
			RECT	181.343 77.844 181.375 77.908 ;
			RECT	181.511 77.844 181.543 77.908 ;
			RECT	181.679 77.844 181.711 77.908 ;
			RECT	181.847 77.844 181.879 77.908 ;
			RECT	182.015 77.844 182.047 77.908 ;
			RECT	182.183 77.844 182.215 77.908 ;
			RECT	182.351 77.844 182.383 77.908 ;
			RECT	182.519 77.844 182.551 77.908 ;
			RECT	182.687 77.844 182.719 77.908 ;
			RECT	182.855 77.844 182.887 77.908 ;
			RECT	183.023 77.844 183.055 77.908 ;
			RECT	183.191 77.844 183.223 77.908 ;
			RECT	183.359 77.844 183.391 77.908 ;
			RECT	183.527 77.844 183.559 77.908 ;
			RECT	183.695 77.844 183.727 77.908 ;
			RECT	183.863 77.844 183.895 77.908 ;
			RECT	184.031 77.844 184.063 77.908 ;
			RECT	184.199 77.844 184.231 77.908 ;
			RECT	184.367 77.844 184.399 77.908 ;
			RECT	184.535 77.844 184.567 77.908 ;
			RECT	184.703 77.844 184.735 77.908 ;
			RECT	184.871 77.844 184.903 77.908 ;
			RECT	185.039 77.844 185.071 77.908 ;
			RECT	185.207 77.844 185.239 77.908 ;
			RECT	185.375 77.844 185.407 77.908 ;
			RECT	185.543 77.844 185.575 77.908 ;
			RECT	185.711 77.844 185.743 77.908 ;
			RECT	185.879 77.844 185.911 77.908 ;
			RECT	186.047 77.844 186.079 77.908 ;
			RECT	186.215 77.844 186.247 77.908 ;
			RECT	186.383 77.844 186.415 77.908 ;
			RECT	186.551 77.844 186.583 77.908 ;
			RECT	186.719 77.844 186.751 77.908 ;
			RECT	186.887 77.844 186.919 77.908 ;
			RECT	187.055 77.844 187.087 77.908 ;
			RECT	187.223 77.844 187.255 77.908 ;
			RECT	187.391 77.844 187.423 77.908 ;
			RECT	187.559 77.844 187.591 77.908 ;
			RECT	187.727 77.844 187.759 77.908 ;
			RECT	187.895 77.844 187.927 77.908 ;
			RECT	188.063 77.844 188.095 77.908 ;
			RECT	188.231 77.844 188.263 77.908 ;
			RECT	188.399 77.844 188.431 77.908 ;
			RECT	188.567 77.844 188.599 77.908 ;
			RECT	188.735 77.844 188.767 77.908 ;
			RECT	188.903 77.844 188.935 77.908 ;
			RECT	189.071 77.844 189.103 77.908 ;
			RECT	189.239 77.844 189.271 77.908 ;
			RECT	189.407 77.844 189.439 77.908 ;
			RECT	189.575 77.844 189.607 77.908 ;
			RECT	189.743 77.844 189.775 77.908 ;
			RECT	189.911 77.844 189.943 77.908 ;
			RECT	190.079 77.844 190.111 77.908 ;
			RECT	190.247 77.844 190.279 77.908 ;
			RECT	190.415 77.844 190.447 77.908 ;
			RECT	190.583 77.844 190.615 77.908 ;
			RECT	190.751 77.844 190.783 77.908 ;
			RECT	190.919 77.844 190.951 77.908 ;
			RECT	191.087 77.844 191.119 77.908 ;
			RECT	191.255 77.844 191.287 77.908 ;
			RECT	191.423 77.844 191.455 77.908 ;
			RECT	191.591 77.844 191.623 77.908 ;
			RECT	191.759 77.844 191.791 77.908 ;
			RECT	191.927 77.844 191.959 77.908 ;
			RECT	192.095 77.844 192.127 77.908 ;
			RECT	192.263 77.844 192.295 77.908 ;
			RECT	192.431 77.844 192.463 77.908 ;
			RECT	192.599 77.844 192.631 77.908 ;
			RECT	192.767 77.844 192.799 77.908 ;
			RECT	192.935 77.844 192.967 77.908 ;
			RECT	193.103 77.844 193.135 77.908 ;
			RECT	193.271 77.844 193.303 77.908 ;
			RECT	193.439 77.844 193.471 77.908 ;
			RECT	193.607 77.844 193.639 77.908 ;
			RECT	193.775 77.844 193.807 77.908 ;
			RECT	193.943 77.844 193.975 77.908 ;
			RECT	194.111 77.844 194.143 77.908 ;
			RECT	194.279 77.844 194.311 77.908 ;
			RECT	194.447 77.844 194.479 77.908 ;
			RECT	194.615 77.844 194.647 77.908 ;
			RECT	194.783 77.844 194.815 77.908 ;
			RECT	194.951 77.844 194.983 77.908 ;
			RECT	195.119 77.844 195.151 77.908 ;
			RECT	195.287 77.844 195.319 77.908 ;
			RECT	195.455 77.844 195.487 77.908 ;
			RECT	195.623 77.844 195.655 77.908 ;
			RECT	195.791 77.844 195.823 77.908 ;
			RECT	195.959 77.844 195.991 77.908 ;
			RECT	196.127 77.844 196.159 77.908 ;
			RECT	196.295 77.844 196.327 77.908 ;
			RECT	196.463 77.844 196.495 77.908 ;
			RECT	196.631 77.844 196.663 77.908 ;
			RECT	196.799 77.844 196.831 77.908 ;
			RECT	196.967 77.844 196.999 77.908 ;
			RECT	197.135 77.844 197.167 77.908 ;
			RECT	197.303 77.844 197.335 77.908 ;
			RECT	197.471 77.844 197.503 77.908 ;
			RECT	197.639 77.844 197.671 77.908 ;
			RECT	197.807 77.844 197.839 77.908 ;
			RECT	197.975 77.844 198.007 77.908 ;
			RECT	198.143 77.844 198.175 77.908 ;
			RECT	198.311 77.844 198.343 77.908 ;
			RECT	198.479 77.844 198.511 77.908 ;
			RECT	198.647 77.844 198.679 77.908 ;
			RECT	198.815 77.844 198.847 77.908 ;
			RECT	198.983 77.844 199.015 77.908 ;
			RECT	199.151 77.844 199.183 77.908 ;
			RECT	199.319 77.844 199.351 77.908 ;
			RECT	199.487 77.844 199.519 77.908 ;
			RECT	199.655 77.844 199.687 77.908 ;
			RECT	199.823 77.844 199.855 77.908 ;
			RECT	199.991 77.844 200.023 77.908 ;
			RECT	200.121 77.86 200.153 77.892 ;
			RECT	200.243 77.855 200.275 77.887 ;
			RECT	200.373 77.844 200.405 77.908 ;
			RECT	200.9 77.844 200.932 77.908 ;
		END

	END VSSE

	PIN WEN[0]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 2.293 0.18 2.363 ;
			LAYER	M2 ;
			RECT	0 2.292 0.134 2.364 ;
			LAYER	M3 ;
			RECT	0 2.292 0.134 2.364 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[0]

	PIN WEN[10]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 21.493 0.18 21.563 ;
			LAYER	M2 ;
			RECT	0 21.492 0.134 21.564 ;
			LAYER	M3 ;
			RECT	0 21.492 0.134 21.564 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[10]

	PIN WEN[11]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 23.413 0.18 23.483 ;
			LAYER	M2 ;
			RECT	0 23.412 0.134 23.484 ;
			LAYER	M3 ;
			RECT	0 23.412 0.134 23.484 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[11]

	PIN WEN[12]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 25.333 0.18 25.403 ;
			LAYER	M2 ;
			RECT	0 25.332 0.134 25.404 ;
			LAYER	M3 ;
			RECT	0 25.332 0.134 25.404 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[12]

	PIN WEN[13]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 27.253 0.18 27.323 ;
			LAYER	M2 ;
			RECT	0 27.252 0.134 27.324 ;
			LAYER	M3 ;
			RECT	0 27.252 0.134 27.324 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[13]

	PIN WEN[14]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 29.173 0.18 29.243 ;
			LAYER	M2 ;
			RECT	0 29.172 0.134 29.244 ;
			LAYER	M3 ;
			RECT	0 29.172 0.134 29.244 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[14]

	PIN WEN[15]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 31.093 0.18 31.163 ;
			LAYER	M2 ;
			RECT	0 31.092 0.134 31.164 ;
			LAYER	M3 ;
			RECT	0 31.092 0.134 31.164 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[15]

	PIN WEN[16]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 51.013 0.18 51.083 ;
			LAYER	M2 ;
			RECT	0 51.012 0.134 51.084 ;
			LAYER	M3 ;
			RECT	0 51.012 0.134 51.084 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[16]

	PIN WEN[17]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 52.933 0.18 53.003 ;
			LAYER	M2 ;
			RECT	0 52.932 0.134 53.004 ;
			LAYER	M3 ;
			RECT	0 52.932 0.134 53.004 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[17]

	PIN WEN[18]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 54.853 0.18 54.923 ;
			LAYER	M2 ;
			RECT	0 54.852 0.134 54.924 ;
			LAYER	M3 ;
			RECT	0 54.852 0.134 54.924 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[18]

	PIN WEN[19]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 56.773 0.18 56.843 ;
			LAYER	M2 ;
			RECT	0 56.772 0.134 56.844 ;
			LAYER	M3 ;
			RECT	0 56.772 0.134 56.844 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[19]

	PIN WEN[1]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 4.213 0.18 4.283 ;
			LAYER	M2 ;
			RECT	0 4.212 0.134 4.284 ;
			LAYER	M3 ;
			RECT	0 4.212 0.134 4.284 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[1]

	PIN WEN[20]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 58.693 0.18 58.763 ;
			LAYER	M2 ;
			RECT	0 58.692 0.134 58.764 ;
			LAYER	M3 ;
			RECT	0 58.692 0.134 58.764 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[20]

	PIN WEN[21]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 60.613 0.18 60.683 ;
			LAYER	M2 ;
			RECT	0 60.612 0.134 60.684 ;
			LAYER	M3 ;
			RECT	0 60.612 0.134 60.684 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[21]

	PIN WEN[22]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 62.533 0.18 62.603 ;
			LAYER	M2 ;
			RECT	0 62.532 0.134 62.604 ;
			LAYER	M3 ;
			RECT	0 62.532 0.134 62.604 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[22]

	PIN WEN[23]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 64.453 0.18 64.523 ;
			LAYER	M2 ;
			RECT	0 64.452 0.134 64.524 ;
			LAYER	M3 ;
			RECT	0 64.452 0.134 64.524 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[23]

	PIN WEN[24]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 66.373 0.18 66.443 ;
			LAYER	M2 ;
			RECT	0 66.372 0.134 66.444 ;
			LAYER	M3 ;
			RECT	0 66.372 0.134 66.444 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[24]

	PIN WEN[25]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 68.293 0.18 68.363 ;
			LAYER	M2 ;
			RECT	0 68.292 0.134 68.364 ;
			LAYER	M3 ;
			RECT	0 68.292 0.134 68.364 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[25]

	PIN WEN[26]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 70.213 0.18 70.283 ;
			LAYER	M2 ;
			RECT	0 70.212 0.134 70.284 ;
			LAYER	M3 ;
			RECT	0 70.212 0.134 70.284 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[26]

	PIN WEN[27]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 72.133 0.18 72.203 ;
			LAYER	M2 ;
			RECT	0 72.132 0.134 72.204 ;
			LAYER	M3 ;
			RECT	0 72.132 0.134 72.204 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[27]

	PIN WEN[28]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 74.053 0.18 74.123 ;
			LAYER	M2 ;
			RECT	0 74.052 0.134 74.124 ;
			LAYER	M3 ;
			RECT	0 74.052 0.134 74.124 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[28]

	PIN WEN[29]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 75.973 0.18 76.043 ;
			LAYER	M2 ;
			RECT	0 75.972 0.134 76.044 ;
			LAYER	M3 ;
			RECT	0 75.972 0.134 76.044 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[29]

	PIN WEN[2]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 6.133 0.18 6.203 ;
			LAYER	M2 ;
			RECT	0 6.132 0.134 6.204 ;
			LAYER	M3 ;
			RECT	0 6.132 0.134 6.204 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[2]

	PIN WEN[30]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 77.893 0.18 77.963 ;
			LAYER	M2 ;
			RECT	0 77.892 0.134 77.964 ;
			LAYER	M3 ;
			RECT	0 77.892 0.134 77.964 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[30]

	PIN WEN[31]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 79.813 0.18 79.883 ;
			LAYER	M2 ;
			RECT	0 79.812 0.134 79.884 ;
			LAYER	M3 ;
			RECT	0 79.812 0.134 79.884 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[31]

	PIN WEN[3]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 8.053 0.18 8.123 ;
			LAYER	M2 ;
			RECT	0 8.052 0.134 8.124 ;
			LAYER	M3 ;
			RECT	0 8.052 0.134 8.124 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[3]

	PIN WEN[4]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 9.973 0.18 10.043 ;
			LAYER	M2 ;
			RECT	0 9.972 0.134 10.044 ;
			LAYER	M3 ;
			RECT	0 9.972 0.134 10.044 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[4]

	PIN WEN[5]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 11.893 0.18 11.963 ;
			LAYER	M2 ;
			RECT	0 11.892 0.134 11.964 ;
			LAYER	M3 ;
			RECT	0 11.892 0.134 11.964 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[5]

	PIN WEN[6]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 13.813 0.18 13.883 ;
			LAYER	M2 ;
			RECT	0 13.812 0.134 13.884 ;
			LAYER	M3 ;
			RECT	0 13.812 0.134 13.884 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[6]

	PIN WEN[7]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 15.733 0.18 15.803 ;
			LAYER	M2 ;
			RECT	0 15.732 0.134 15.804 ;
			LAYER	M3 ;
			RECT	0 15.732 0.134 15.804 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[7]

	PIN WEN[8]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 17.653 0.18 17.723 ;
			LAYER	M2 ;
			RECT	0 17.652 0.134 17.724 ;
			LAYER	M3 ;
			RECT	0 17.652 0.134 17.724 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[8]

	PIN WEN[9]
		USE SIGNAL ;
		DIRECTION INPUT ;
		SHAPE ABUTMENT ;
		PORT
			LAYER	C4 ;
			RECT	0 19.573 0.18 19.643 ;
			LAYER	M2 ;
			RECT	0 19.572 0.134 19.644 ;
			LAYER	M3 ;
			RECT	0 19.572 0.134 19.644 ;
		END

		ANTENNAGATEAREA 0.003072 ;
		ANTENNADIFFAREA 0.00252 ;
	END WEN[9]

	OBS
		LAYER	C4 DESIGNRULEWIDTH 0.04 ;
		RECT	0.294 0 201.485 0.168 ;
		RECT	201.485 0 201.665 0.168 ;
		RECT	0.294 1.01 201.485 1.165 ;
		RECT	201.485 1.01 201.665 1.165 ;
		RECT	0.294 1.445 201.485 2.235 ;
		RECT	201.485 1.445 201.665 2.235 ;
		RECT	0.294 2.93 201.485 3.085 ;
		RECT	201.485 2.93 201.665 3.085 ;
		RECT	0.294 3.365 201.485 4.155 ;
		RECT	201.485 3.365 201.665 4.155 ;
		RECT	0.294 4.85 201.485 5.005 ;
		RECT	201.485 4.85 201.665 5.005 ;
		RECT	0.294 5.285 201.485 6.075 ;
		RECT	201.485 5.285 201.665 6.075 ;
		RECT	0.294 6.77 201.485 6.925 ;
		RECT	201.485 6.77 201.665 6.925 ;
		RECT	0.294 7.205 201.485 7.995 ;
		RECT	201.485 7.205 201.665 7.995 ;
		RECT	0.294 8.69 201.485 8.845 ;
		RECT	201.485 8.69 201.665 8.845 ;
		RECT	0.294 9.125 201.485 9.915 ;
		RECT	201.485 9.125 201.665 9.915 ;
		RECT	0.294 10.61 201.485 10.765 ;
		RECT	201.485 10.61 201.665 10.765 ;
		RECT	0.294 11.045 201.485 11.835 ;
		RECT	201.485 11.045 201.665 11.835 ;
		RECT	0.294 12.53 201.485 12.685 ;
		RECT	201.485 12.53 201.665 12.685 ;
		RECT	0.294 12.965 201.485 13.755 ;
		RECT	201.485 12.965 201.665 13.755 ;
		RECT	0.294 14.45 201.485 14.605 ;
		RECT	201.485 14.45 201.665 14.605 ;
		RECT	0.294 14.885 201.485 15.675 ;
		RECT	201.485 14.885 201.665 15.675 ;
		RECT	0.294 16.37 201.485 16.525 ;
		RECT	201.485 16.37 201.665 16.525 ;
		RECT	0.294 16.805 201.485 17.595 ;
		RECT	201.485 16.805 201.665 17.595 ;
		RECT	0.294 18.29 201.485 18.445 ;
		RECT	201.485 18.29 201.665 18.445 ;
		RECT	0.294 18.725 201.485 19.515 ;
		RECT	201.485 18.725 201.665 19.515 ;
		RECT	0.294 20.21 201.485 20.365 ;
		RECT	201.485 20.21 201.665 20.365 ;
		RECT	0.294 20.645 201.485 21.435 ;
		RECT	201.485 20.645 201.665 21.435 ;
		RECT	0.294 22.13 201.485 22.285 ;
		RECT	201.485 22.13 201.665 22.285 ;
		RECT	0.294 22.565 201.485 23.355 ;
		RECT	201.485 22.565 201.665 23.355 ;
		RECT	0.294 24.05 201.485 24.205 ;
		RECT	201.485 24.05 201.665 24.205 ;
		RECT	0.294 24.485 201.485 25.275 ;
		RECT	201.485 24.485 201.665 25.275 ;
		RECT	0.294 25.97 201.485 26.125 ;
		RECT	201.485 25.97 201.665 26.125 ;
		RECT	0.294 26.405 201.485 27.195 ;
		RECT	201.485 26.405 201.665 27.195 ;
		RECT	0.294 27.89 201.485 28.045 ;
		RECT	201.485 27.89 201.665 28.045 ;
		RECT	0.294 28.325 201.485 29.115 ;
		RECT	201.485 28.325 201.665 29.115 ;
		RECT	0.294 29.81 201.485 29.965 ;
		RECT	201.485 29.81 201.665 29.965 ;
		RECT	0.294 30.245 201.485 31.035 ;
		RECT	201.485 30.245 201.665 31.035 ;
		RECT	0.294 31.733 201.485 31.823 ;
		RECT	201.485 31.733 201.665 31.823 ;
		RECT	0.294 32.103 201.485 32.163 ;
		RECT	201.485 32.103 201.665 32.163 ;
		RECT	0.294 32.663 201.485 32.988 ;
		RECT	201.485 32.663 201.665 32.988 ;
		RECT	0.294 33.433 201.485 33.937 ;
		RECT	201.485 33.433 201.665 33.937 ;
		RECT	0.294 34.637 201.485 34.937 ;
		RECT	201.485 34.637 201.665 34.937 ;
		RECT	0.294 35.227 201.485 35.277 ;
		RECT	201.485 35.227 201.665 35.277 ;
		RECT	0.294 35.732 201.485 35.989 ;
		RECT	201.485 35.732 201.665 35.989 ;
		RECT	0.294 36.229 201.485 36.595 ;
		RECT	201.485 36.229 201.665 36.595 ;
		RECT	0.294 37.46 201.485 37.74 ;
		RECT	201.485 37.46 201.665 37.74 ;
		RECT	0.294 38.352 201.485 38.402 ;
		RECT	201.485 38.352 201.665 38.402 ;
		RECT	0.294 38.642 201.485 38.692 ;
		RECT	201.485 38.642 201.665 38.692 ;
		RECT	0.294 39.149 201.485 39.899 ;
		RECT	201.485 39.149 201.665 39.899 ;
		RECT	0.294 40.354 201.485 40.654 ;
		RECT	201.485 40.354 201.665 40.654 ;
		RECT	0.294 40.894 201.485 41.045 ;
		RECT	201.485 40.894 201.665 41.045 ;
		RECT	0.294 41.521 201.485 41.571 ;
		RECT	201.485 41.521 201.665 41.571 ;
		RECT	0.294 41.861 201.485 42.011 ;
		RECT	201.485 41.861 201.665 42.011 ;
		RECT	0.294 42.416 201.485 43.166 ;
		RECT	201.485 42.416 201.665 43.166 ;
		RECT	0.294 43.406 201.485 43.513 ;
		RECT	201.485 43.406 201.665 43.513 ;
		RECT	0.294 44.008 201.485 44.51 ;
		RECT	201.485 44.008 201.665 44.51 ;
		RECT	0.294 44.75 201.485 44.904 ;
		RECT	201.485 44.75 201.665 44.904 ;
		RECT	0.294 45.144 201.485 45.338 ;
		RECT	201.485 45.144 201.665 45.338 ;
		RECT	0.294 46.048 201.485 46.288 ;
		RECT	201.485 46.048 201.665 46.288 ;
		RECT	0.294 46.528 201.485 46.668 ;
		RECT	201.485 46.528 201.665 46.668 ;
		RECT	0.294 47.358 201.485 47.508 ;
		RECT	201.485 47.358 201.665 47.508 ;
		RECT	0.294 48.208 201.485 48.358 ;
		RECT	201.485 48.208 201.665 48.358 ;
		RECT	0.294 48.648 201.485 48.743 ;
		RECT	201.485 48.648 201.665 48.743 ;
		RECT	0.294 49.188 201.485 49.345 ;
		RECT	201.485 49.188 201.665 49.345 ;
		RECT	0.294 50.013 201.485 50.073 ;
		RECT	201.485 50.013 201.665 50.073 ;
		RECT	0.294 50.353 201.485 50.443 ;
		RECT	201.485 50.353 201.665 50.443 ;
		RECT	0.294 51.141 201.485 51.931 ;
		RECT	201.485 51.141 201.665 51.931 ;
		RECT	0.294 52.211 201.485 52.366 ;
		RECT	201.485 52.211 201.665 52.366 ;
		RECT	0.294 53.061 201.485 53.851 ;
		RECT	201.485 53.061 201.665 53.851 ;
		RECT	0.294 54.131 201.485 54.286 ;
		RECT	201.485 54.131 201.665 54.286 ;
		RECT	0.294 54.981 201.485 55.771 ;
		RECT	201.485 54.981 201.665 55.771 ;
		RECT	0.294 56.051 201.485 56.206 ;
		RECT	201.485 56.051 201.665 56.206 ;
		RECT	0.294 56.901 201.485 57.691 ;
		RECT	201.485 56.901 201.665 57.691 ;
		RECT	0.294 57.971 201.485 58.126 ;
		RECT	201.485 57.971 201.665 58.126 ;
		RECT	0.294 58.821 201.485 59.611 ;
		RECT	201.485 58.821 201.665 59.611 ;
		RECT	0.294 59.891 201.485 60.046 ;
		RECT	201.485 59.891 201.665 60.046 ;
		RECT	0.294 60.741 201.485 61.531 ;
		RECT	201.485 60.741 201.665 61.531 ;
		RECT	0.294 61.811 201.485 61.966 ;
		RECT	201.485 61.811 201.665 61.966 ;
		RECT	0.294 62.661 201.485 63.451 ;
		RECT	201.485 62.661 201.665 63.451 ;
		RECT	0.294 63.731 201.485 63.886 ;
		RECT	201.485 63.731 201.665 63.886 ;
		RECT	0.294 64.581 201.485 65.371 ;
		RECT	201.485 64.581 201.665 65.371 ;
		RECT	0.294 65.651 201.485 65.806 ;
		RECT	201.485 65.651 201.665 65.806 ;
		RECT	0.294 66.501 201.485 67.291 ;
		RECT	201.485 66.501 201.665 67.291 ;
		RECT	0.294 67.571 201.485 67.726 ;
		RECT	201.485 67.571 201.665 67.726 ;
		RECT	0.294 68.421 201.485 69.211 ;
		RECT	201.485 68.421 201.665 69.211 ;
		RECT	0.294 69.491 201.485 69.646 ;
		RECT	201.485 69.491 201.665 69.646 ;
		RECT	0.294 70.341 201.485 71.131 ;
		RECT	201.485 70.341 201.665 71.131 ;
		RECT	0.294 71.411 201.485 71.566 ;
		RECT	201.485 71.411 201.665 71.566 ;
		RECT	0.294 72.261 201.485 73.051 ;
		RECT	201.485 72.261 201.665 73.051 ;
		RECT	0.294 73.331 201.485 73.486 ;
		RECT	201.485 73.331 201.665 73.486 ;
		RECT	0.294 74.181 201.485 74.971 ;
		RECT	201.485 74.181 201.665 74.971 ;
		RECT	0.294 75.251 201.485 75.406 ;
		RECT	201.485 75.251 201.665 75.406 ;
		RECT	0.294 76.101 201.485 76.891 ;
		RECT	201.485 76.101 201.665 76.891 ;
		RECT	0.294 77.171 201.485 77.326 ;
		RECT	201.485 77.171 201.665 77.326 ;
		RECT	0.294 78.021 201.485 78.811 ;
		RECT	201.485 78.021 201.665 78.811 ;
		RECT	0.294 79.091 201.485 79.246 ;
		RECT	201.485 79.091 201.665 79.246 ;
		RECT	0.294 79.941 201.485 80.731 ;
		RECT	201.485 79.941 201.665 80.731 ;
		RECT	0.294 81.011 201.485 81.166 ;
		RECT	201.485 81.011 201.665 81.166 ;
		RECT	0.294 82.008 201.485 82.176 ;
		RECT	201.485 82.008 201.665 82.176 ;
		RECT	0 0 0.18 0.884 ;
		RECT	0 1.084 0.18 1.367 ;
		RECT	0 1.567 0.18 2.228 ;
		RECT	0 2.428 0.18 2.804 ;
		RECT	0 3.004 0.18 3.287 ;
		RECT	0 3.487 0.18 4.148 ;
		RECT	0 4.348 0.18 4.724 ;
		RECT	0 4.924 0.18 5.207 ;
		RECT	0 5.407 0.18 6.068 ;
		RECT	0 6.268 0.18 6.644 ;
		RECT	0 6.844 0.18 7.127 ;
		RECT	0 7.327 0.18 7.988 ;
		RECT	0 8.188 0.18 8.564 ;
		RECT	0 8.764 0.18 9.047 ;
		RECT	0 9.247 0.18 9.908 ;
		RECT	0 10.108 0.18 10.484 ;
		RECT	0 10.684 0.18 10.967 ;
		RECT	0 11.167 0.18 11.828 ;
		RECT	0 12.028 0.18 12.404 ;
		RECT	0 12.604 0.18 12.887 ;
		RECT	0 13.087 0.18 13.748 ;
		RECT	0 13.948 0.18 14.324 ;
		RECT	0 14.524 0.18 14.807 ;
		RECT	0 15.007 0.18 15.668 ;
		RECT	0 15.868 0.18 16.244 ;
		RECT	0 16.444 0.18 16.727 ;
		RECT	0 16.927 0.18 17.588 ;
		RECT	0 17.788 0.18 18.164 ;
		RECT	0 18.364 0.18 18.647 ;
		RECT	0 18.847 0.18 19.508 ;
		RECT	0 19.708 0.18 20.084 ;
		RECT	0 20.284 0.18 20.567 ;
		RECT	0 20.767 0.18 21.428 ;
		RECT	0 21.628 0.18 22.004 ;
		RECT	0 22.204 0.18 22.487 ;
		RECT	0 22.687 0.18 23.348 ;
		RECT	0 23.548 0.18 23.924 ;
		RECT	0 24.124 0.18 24.407 ;
		RECT	0 24.607 0.18 25.268 ;
		RECT	0 25.468 0.18 25.844 ;
		RECT	0 26.044 0.18 26.327 ;
		RECT	0 26.527 0.18 27.188 ;
		RECT	0 27.388 0.18 27.764 ;
		RECT	0 27.964 0.18 28.247 ;
		RECT	0 28.447 0.18 29.108 ;
		RECT	0 29.308 0.18 29.684 ;
		RECT	0 29.884 0.18 30.167 ;
		RECT	0 30.367 0.18 31.028 ;
		RECT	0 31.228 0.18 33.908 ;
		RECT	0 34.444 0.18 34.532 ;
		RECT	0 34.732 0.18 35.06 ;
		RECT	0 35.404 0.18 35.54 ;
		RECT	0 35.884 0.18 37.268 ;
		RECT	0 37.66 0.18 37.94 ;
		RECT	0 38.14 0.18 39.188 ;
		RECT	0 39.58 0.18 39.86 ;
		RECT	0 40.06 0.18 40.484 ;
		RECT	0 40.684 0.18 40.964 ;
		RECT	0 41.164 0.18 41.492 ;
		RECT	0 41.692 0.18 41.972 ;
		RECT	0 42.364 0.18 43.652 ;
		RECT	0 43.852 0.18 44.132 ;
		RECT	0 44.332 0.18 44.996 ;
		RECT	0 45.196 0.18 47.54 ;
		RECT	0 47.74 0.18 50.948 ;
		RECT	0 51.148 0.18 51.809 ;
		RECT	0 52.009 0.18 52.292 ;
		RECT	0 52.492 0.18 52.868 ;
		RECT	0 53.068 0.18 53.729 ;
		RECT	0 53.929 0.18 54.212 ;
		RECT	0 54.412 0.18 54.788 ;
		RECT	0 54.988 0.18 55.649 ;
		RECT	0 55.849 0.18 56.132 ;
		RECT	0 56.332 0.18 56.708 ;
		RECT	0 56.908 0.18 57.569 ;
		RECT	0 57.769 0.18 58.052 ;
		RECT	0 58.252 0.18 58.628 ;
		RECT	0 58.828 0.18 59.489 ;
		RECT	0 59.689 0.18 59.972 ;
		RECT	0 60.172 0.18 60.548 ;
		RECT	0 60.748 0.18 61.409 ;
		RECT	0 61.609 0.18 61.892 ;
		RECT	0 62.092 0.18 62.468 ;
		RECT	0 62.668 0.18 63.329 ;
		RECT	0 63.529 0.18 63.812 ;
		RECT	0 64.012 0.18 64.388 ;
		RECT	0 64.588 0.18 65.249 ;
		RECT	0 65.449 0.18 65.732 ;
		RECT	0 65.932 0.18 66.308 ;
		RECT	0 66.508 0.18 67.169 ;
		RECT	0 67.369 0.18 67.652 ;
		RECT	0 67.852 0.18 68.228 ;
		RECT	0 68.428 0.18 69.089 ;
		RECT	0 69.289 0.18 69.572 ;
		RECT	0 69.772 0.18 70.148 ;
		RECT	0 70.348 0.18 71.009 ;
		RECT	0 71.209 0.18 71.492 ;
		RECT	0 71.692 0.18 72.068 ;
		RECT	0 72.268 0.18 72.929 ;
		RECT	0 73.129 0.18 73.412 ;
		RECT	0 73.612 0.18 73.988 ;
		RECT	0 74.188 0.18 74.849 ;
		RECT	0 75.049 0.18 75.332 ;
		RECT	0 75.532 0.18 75.908 ;
		RECT	0 76.108 0.18 76.769 ;
		RECT	0 76.969 0.18 77.252 ;
		RECT	0 77.452 0.18 77.828 ;
		RECT	0 78.028 0.18 78.689 ;
		RECT	0 78.889 0.18 79.172 ;
		RECT	0 79.372 0.18 79.748 ;
		RECT	0 79.948 0.18 80.609 ;
		RECT	0 80.809 0.18 81.092 ;
		RECT	0.18 0 0.294 82.176 ;
		RECT	0 81.292 0.18 82.176 ;
		LAYER	J3 DESIGNRULEWIDTH 0 ;
		RECT	0.674 31.752 0.706 31.784 ;
		RECT	0.885 32.117 0.917 32.149 ;
		RECT	0.047 32.168 0.111 32.2 ;
		RECT	0.047 32.36 0.111 32.392 ;
		RECT	0.047 32.504 0.111 32.536 ;
		RECT	0.755 32.691 0.787 32.755 ;
		RECT	0.601 32.892 0.633 32.924 ;
		RECT	0.047 33.173 0.111 33.205 ;
		RECT	0.047 33.32 0.111 33.352 ;
		RECT	0.047 33.512 0.111 33.544 ;
		RECT	0.639 33.601 0.671 33.633 ;
		RECT	0.047 33.656 0.111 33.688 ;
		RECT	0.729 33.696 0.761 33.728 ;
		RECT	0.556 33.796 0.588 33.828 ;
		RECT	0.047 33.848 0.111 33.88 ;
		RECT	0.47 33.896 0.502 33.928 ;
		RECT	0.047 33.992 0.111 34.024 ;
		RECT	0.047 34.136 0.111 34.168 ;
		RECT	0.047 34.328 0.111 34.36 ;
		RECT	0.047 34.472 0.111 34.504 ;
		RECT	0.047 34.616 0.111 34.648 ;
		RECT	1.234 34.641 1.266 34.673 ;
		RECT	1.164 34.721 1.196 34.753 ;
		RECT	0.047 34.76 0.111 34.792 ;
		RECT	0.642 34.801 0.674 34.833 ;
		RECT	0.812 34.896 0.844 34.928 ;
		RECT	0.047 35 0.111 35.032 ;
		RECT	0.047 35.144 0.111 35.176 ;
		RECT	0.047 35.288 0.111 35.32 ;
		RECT	0.047 35.48 0.111 35.512 ;
		RECT	0.047 35.624 0.111 35.656 ;
		RECT	0.047 35.768 0.111 35.8 ;
		RECT	0.857 35.948 0.889 35.98 ;
		RECT	0.047 35.96 0.111 35.992 ;
		RECT	0.047 36.104 0.111 36.136 ;
		RECT	0.642 36.238 0.674 36.27 ;
		RECT	0.047 36.248 0.111 36.28 ;
		RECT	0.729 36.338 0.761 36.37 ;
		RECT	0.047 36.44 0.111 36.472 ;
		RECT	0.645 36.454 0.677 36.486 ;
		RECT	0.856 36.554 0.888 36.586 ;
		RECT	0.047 36.592 0.111 36.624 ;
		RECT	0.047 36.776 0.111 36.808 ;
		RECT	0.047 36.92 0.111 36.952 ;
		RECT	0.047 37.064 0.111 37.096 ;
		RECT	0.047 37.208 0.111 37.24 ;
		RECT	0.047 37.352 0.111 37.384 ;
		RECT	0.71 37.474 0.742 37.506 ;
		RECT	0.047 37.544 0.111 37.576 ;
		RECT	0.385 37.589 0.417 37.621 ;
		RECT	0.047 37.688 0.111 37.72 ;
		RECT	0.646 37.689 0.678 37.721 ;
		RECT	0.047 37.88 0.111 37.912 ;
		RECT	0.047 38.024 0.111 38.056 ;
		RECT	0.047 38.189 0.111 38.221 ;
		RECT	0.781 38.361 0.813 38.393 ;
		RECT	0.047 38.392 0.111 38.424 ;
		RECT	0.047 38.618 0.111 38.65 ;
		RECT	0.642 38.651 0.674 38.683 ;
		RECT	0.047 38.792 0.111 38.824 ;
		RECT	0.047 38.936 0.111 38.968 ;
		RECT	0.047 39.128 0.111 39.16 ;
		RECT	0.047 39.272 0.111 39.304 ;
		RECT	0.047 39.464 0.111 39.496 ;
		RECT	0.047 39.608 0.111 39.64 ;
		RECT	0.047 39.944 0.111 39.976 ;
		RECT	0.047 40.098 0.111 40.13 ;
		RECT	0.047 40.242 0.111 40.274 ;
		RECT	0.642 40.363 0.674 40.395 ;
		RECT	0.047 40.424 0.111 40.456 ;
		RECT	0.781 40.458 0.813 40.49 ;
		RECT	0.711 40.538 0.743 40.57 ;
		RECT	0.047 40.568 0.111 40.6 ;
		RECT	0.642 40.618 0.674 40.65 ;
		RECT	0.047 40.712 0.111 40.744 ;
		RECT	0.856 40.903 0.888 40.935 ;
		RECT	0.047 40.904 0.111 40.936 ;
		RECT	0.783 41.004 0.815 41.036 ;
		RECT	0.047 41.048 0.111 41.08 ;
		RECT	0.047 41.24 0.111 41.272 ;
		RECT	0.047 41.384 0.111 41.416 ;
		RECT	0.781 41.53 0.813 41.562 ;
		RECT	0.047 41.576 0.111 41.608 ;
		RECT	0.047 41.76 0.111 41.792 ;
		RECT	0.556 41.87 0.588 41.902 ;
		RECT	0.047 41.91 0.111 41.942 ;
		RECT	0.711 41.97 0.743 42.002 ;
		RECT	0.047 42.056 0.111 42.088 ;
		RECT	0.047 42.248 0.111 42.28 ;
		RECT	0.047 42.488 0.111 42.52 ;
		RECT	0.47 42.525 0.502 42.557 ;
		RECT	0.047 42.68 0.111 42.712 ;
		RECT	0.047 42.92 0.111 42.952 ;
		RECT	0.047 43.112 0.111 43.144 ;
		RECT	0.047 43.268 0.111 43.3 ;
		RECT	0.047 43.416 0.111 43.448 ;
		RECT	0.047 43.566 0.111 43.598 ;
		RECT	0.047 43.736 0.111 43.768 ;
		RECT	0.047 43.88 0.111 43.912 ;
		RECT	0.047 44.072 0.111 44.104 ;
		RECT	0.634 44.199 0.666 44.231 ;
		RECT	0.047 44.216 0.111 44.248 ;
		RECT	0.703 44.294 0.735 44.326 ;
		RECT	0.781 44.374 0.813 44.406 ;
		RECT	0.047 44.408 0.111 44.44 ;
		RECT	0.385 44.469 0.417 44.501 ;
		RECT	0.047 44.552 0.111 44.584 ;
		RECT	0.047 44.744 0.111 44.776 ;
		RECT	0.372 44.759 0.404 44.791 ;
		RECT	0.047 44.888 0.111 44.92 ;
		RECT	0.047 45.08 0.111 45.112 ;
		RECT	0.47 45.197 0.502 45.229 ;
		RECT	0.047 45.311 0.111 45.343 ;
		RECT	0.047 45.495 0.111 45.527 ;
		RECT	0.047 45.752 0.111 45.784 ;
		RECT	0.047 45.896 0.111 45.928 ;
		RECT	0.729 46.057 0.761 46.089 ;
		RECT	0.047 46.088 0.111 46.12 ;
		RECT	0.654 46.157 0.686 46.189 ;
		RECT	0.047 46.28 0.111 46.312 ;
		RECT	0.047 46.472 0.111 46.504 ;
		RECT	0.627 46.632 0.659 46.664 ;
		RECT	0.047 46.664 0.111 46.696 ;
		RECT	0.047 46.856 0.111 46.888 ;
		RECT	0.047 47 0.111 47.032 ;
		RECT	0.047 47.144 0.111 47.176 ;
		RECT	0.047 47.288 0.111 47.32 ;
		RECT	0.812 47.367 0.844 47.399 ;
		RECT	0.729 47.467 0.761 47.499 ;
		RECT	0.047 47.48 0.111 47.512 ;
		RECT	0.047 47.624 0.111 47.656 ;
		RECT	0.047 47.881 0.111 47.913 ;
		RECT	0.047 48.034 0.111 48.066 ;
		RECT	0.047 48.192 0.111 48.224 ;
		RECT	0.642 48.217 0.674 48.249 ;
		RECT	0.738 48.317 0.77 48.349 ;
		RECT	0.047 48.343 0.111 48.375 ;
		RECT	0.047 48.584 0.111 48.616 ;
		RECT	0.047 48.824 0.111 48.856 ;
		RECT	0.047 49.064 0.111 49.096 ;
		RECT	0.047 49.256 0.111 49.288 ;
		RECT	0.678 49.264 0.71 49.328 ;
		RECT	0.047 49.515 0.111 49.547 ;
		RECT	0.047 49.784 0.111 49.816 ;
		RECT	0.047 49.928 0.111 49.96 ;
		RECT	0.914 50.027 0.946 50.059 ;
		RECT	0.047 50.072 0.111 50.104 ;
		RECT	0.678 50.392 0.71 50.424 ;
		RECT	0.047 2.744 0.111 2.776 ;
		RECT	0.047 2.888 0.111 2.92 ;
		RECT	0.047 3.371 0.111 3.403 ;
		RECT	0.756 3.613 0.788 3.677 ;
		RECT	0.047 4.015 0.111 4.047 ;
		RECT	0.047 4.232 0.111 4.264 ;
		RECT	0.047 4.424 0.111 4.456 ;
		RECT	0.047 20.024 0.111 20.056 ;
		RECT	0.047 20.168 0.111 20.2 ;
		RECT	0.047 20.651 0.111 20.683 ;
		RECT	0.756 20.893 0.788 20.957 ;
		RECT	0.047 21.295 0.111 21.327 ;
		RECT	0.047 21.512 0.111 21.544 ;
		RECT	0.047 21.704 0.111 21.736 ;
		RECT	0.047 21.944 0.111 21.976 ;
		RECT	0.047 22.088 0.111 22.12 ;
		RECT	0.047 22.571 0.111 22.603 ;
		RECT	0.756 22.813 0.788 22.877 ;
		RECT	0.047 23.215 0.111 23.247 ;
		RECT	0.047 23.432 0.111 23.464 ;
		RECT	0.047 23.624 0.111 23.656 ;
		RECT	0.047 23.864 0.111 23.896 ;
		RECT	0.047 24.008 0.111 24.04 ;
		RECT	0.047 24.491 0.111 24.523 ;
		RECT	0.756 24.733 0.788 24.797 ;
		RECT	0.047 25.135 0.111 25.167 ;
		RECT	0.047 25.352 0.111 25.384 ;
		RECT	0.047 25.544 0.111 25.576 ;
		RECT	0.047 25.784 0.111 25.816 ;
		RECT	0.047 25.928 0.111 25.96 ;
		RECT	0.047 26.411 0.111 26.443 ;
		RECT	0.756 26.653 0.788 26.717 ;
		RECT	0.047 27.055 0.111 27.087 ;
		RECT	0.047 27.272 0.111 27.304 ;
		RECT	0.047 27.464 0.111 27.496 ;
		RECT	0.047 27.704 0.111 27.736 ;
		RECT	0.047 27.848 0.111 27.88 ;
		RECT	0.047 28.331 0.111 28.363 ;
		RECT	0.756 28.573 0.788 28.637 ;
		RECT	0.047 28.975 0.111 29.007 ;
		RECT	0.047 29.192 0.111 29.224 ;
		RECT	0.047 29.384 0.111 29.416 ;
		RECT	0.047 4.664 0.111 4.696 ;
		RECT	0.047 4.808 0.111 4.84 ;
		RECT	0.047 5.291 0.111 5.323 ;
		RECT	0.756 5.533 0.788 5.597 ;
		RECT	0.047 5.935 0.111 5.967 ;
		RECT	0.047 6.152 0.111 6.184 ;
		RECT	0.047 6.344 0.111 6.376 ;
		RECT	0.047 6.584 0.111 6.616 ;
		RECT	0.047 6.728 0.111 6.76 ;
		RECT	0.047 7.211 0.111 7.243 ;
		RECT	0.756 7.453 0.788 7.517 ;
		RECT	0.047 7.855 0.111 7.887 ;
		RECT	0.047 8.072 0.111 8.104 ;
		RECT	0.047 8.264 0.111 8.296 ;
		RECT	0.047 8.504 0.111 8.536 ;
		RECT	0.047 8.648 0.111 8.68 ;
		RECT	0.047 9.131 0.111 9.163 ;
		RECT	0.756 9.373 0.788 9.437 ;
		RECT	0.047 9.775 0.111 9.807 ;
		RECT	0.047 9.992 0.111 10.024 ;
		RECT	0.047 10.184 0.111 10.216 ;
		RECT	0.047 10.424 0.111 10.456 ;
		RECT	0.047 10.568 0.111 10.6 ;
		RECT	0.047 11.051 0.111 11.083 ;
		RECT	0.756 11.293 0.788 11.357 ;
		RECT	0.047 11.695 0.111 11.727 ;
		RECT	0.047 11.912 0.111 11.944 ;
		RECT	0.047 12.104 0.111 12.136 ;
		RECT	0.047 12.344 0.111 12.376 ;
		RECT	0.047 12.488 0.111 12.52 ;
		RECT	0.047 12.971 0.111 13.003 ;
		RECT	0.756 13.213 0.788 13.277 ;
		RECT	0.047 13.615 0.111 13.647 ;
		RECT	0.047 13.832 0.111 13.864 ;
		RECT	0.047 14.024 0.111 14.056 ;
		RECT	0.047 14.264 0.111 14.296 ;
		RECT	0.047 14.408 0.111 14.44 ;
		RECT	0.047 14.891 0.111 14.923 ;
		RECT	0.756 15.133 0.788 15.197 ;
		RECT	0.047 15.535 0.111 15.567 ;
		RECT	0.047 15.752 0.111 15.784 ;
		RECT	0.047 15.944 0.111 15.976 ;
		RECT	0.047 16.184 0.111 16.216 ;
		RECT	0.047 16.328 0.111 16.36 ;
		RECT	0.047 16.811 0.111 16.843 ;
		RECT	0.756 17.053 0.788 17.117 ;
		RECT	0.047 17.455 0.111 17.487 ;
		RECT	0.047 17.672 0.111 17.704 ;
		RECT	0.047 17.864 0.111 17.896 ;
		RECT	0.047 18.104 0.111 18.136 ;
		RECT	0.047 18.248 0.111 18.28 ;
		RECT	0.047 18.731 0.111 18.763 ;
		RECT	0.756 18.973 0.788 19.037 ;
		RECT	0.047 19.375 0.111 19.407 ;
		RECT	0.047 19.592 0.111 19.624 ;
		RECT	0.047 19.784 0.111 19.816 ;
		RECT	0.047 0.824 0.111 0.856 ;
		RECT	0.047 0.968 0.111 1 ;
		RECT	0.047 1.451 0.111 1.483 ;
		RECT	0.756 1.693 0.788 1.757 ;
		RECT	0.047 2.095 0.111 2.127 ;
		RECT	0.047 2.312 0.111 2.344 ;
		RECT	0.047 2.504 0.111 2.536 ;
		RECT	0.047 29.624 0.111 29.656 ;
		RECT	0.047 29.768 0.111 29.8 ;
		RECT	0.047 30.251 0.111 30.283 ;
		RECT	0.756 30.493 0.788 30.557 ;
		RECT	0.047 30.895 0.111 30.927 ;
		RECT	0.047 31.112 0.111 31.144 ;
		RECT	0.047 31.304 0.111 31.336 ;
		RECT	0.047 0.248 0.111 0.28 ;
		RECT	0.047 0.44 0.111 0.472 ;
		RECT	0.047 54.44 0.111 54.472 ;
		RECT	0.047 54.296 0.111 54.328 ;
		RECT	0.047 53.813 0.111 53.845 ;
		RECT	0.756 53.539 0.788 53.603 ;
		RECT	0.047 53.169 0.111 53.201 ;
		RECT	0.047 52.952 0.111 52.984 ;
		RECT	0.047 52.76 0.111 52.792 ;
		RECT	0.047 71.72 0.111 71.752 ;
		RECT	0.047 71.576 0.111 71.608 ;
		RECT	0.047 71.093 0.111 71.125 ;
		RECT	0.756 70.819 0.788 70.883 ;
		RECT	0.047 70.449 0.111 70.481 ;
		RECT	0.047 70.232 0.111 70.264 ;
		RECT	0.047 70.04 0.111 70.072 ;
		RECT	0.047 73.64 0.111 73.672 ;
		RECT	0.047 73.496 0.111 73.528 ;
		RECT	0.047 73.013 0.111 73.045 ;
		RECT	0.756 72.739 0.788 72.803 ;
		RECT	0.047 72.369 0.111 72.401 ;
		RECT	0.047 72.152 0.111 72.184 ;
		RECT	0.047 71.96 0.111 71.992 ;
		RECT	0.047 75.56 0.111 75.592 ;
		RECT	0.047 75.416 0.111 75.448 ;
		RECT	0.047 74.933 0.111 74.965 ;
		RECT	0.756 74.659 0.788 74.723 ;
		RECT	0.047 74.289 0.111 74.321 ;
		RECT	0.047 74.072 0.111 74.104 ;
		RECT	0.047 73.88 0.111 73.912 ;
		RECT	0.047 77.48 0.111 77.512 ;
		RECT	0.047 77.336 0.111 77.368 ;
		RECT	0.047 76.853 0.111 76.885 ;
		RECT	0.756 76.579 0.788 76.643 ;
		RECT	0.047 76.209 0.111 76.241 ;
		RECT	0.047 75.992 0.111 76.024 ;
		RECT	0.047 75.8 0.111 75.832 ;
		RECT	0.047 79.4 0.111 79.432 ;
		RECT	0.047 79.256 0.111 79.288 ;
		RECT	0.047 78.773 0.111 78.805 ;
		RECT	0.756 78.499 0.788 78.563 ;
		RECT	0.047 78.129 0.111 78.161 ;
		RECT	0.047 77.912 0.111 77.944 ;
		RECT	0.047 77.72 0.111 77.752 ;
		RECT	0.047 56.36 0.111 56.392 ;
		RECT	0.047 56.216 0.111 56.248 ;
		RECT	0.047 55.733 0.111 55.765 ;
		RECT	0.756 55.459 0.788 55.523 ;
		RECT	0.047 55.089 0.111 55.121 ;
		RECT	0.047 54.872 0.111 54.904 ;
		RECT	0.047 54.68 0.111 54.712 ;
		RECT	0.047 58.28 0.111 58.312 ;
		RECT	0.047 58.136 0.111 58.168 ;
		RECT	0.047 57.653 0.111 57.685 ;
		RECT	0.756 57.379 0.788 57.443 ;
		RECT	0.047 57.009 0.111 57.041 ;
		RECT	0.047 56.792 0.111 56.824 ;
		RECT	0.047 56.6 0.111 56.632 ;
		RECT	0.047 60.2 0.111 60.232 ;
		RECT	0.047 60.056 0.111 60.088 ;
		RECT	0.047 59.573 0.111 59.605 ;
		RECT	0.756 59.299 0.788 59.363 ;
		RECT	0.047 58.929 0.111 58.961 ;
		RECT	0.047 58.712 0.111 58.744 ;
		RECT	0.047 58.52 0.111 58.552 ;
		RECT	0.047 62.12 0.111 62.152 ;
		RECT	0.047 61.976 0.111 62.008 ;
		RECT	0.047 61.493 0.111 61.525 ;
		RECT	0.756 61.219 0.788 61.283 ;
		RECT	0.047 60.849 0.111 60.881 ;
		RECT	0.047 60.632 0.111 60.664 ;
		RECT	0.047 60.44 0.111 60.472 ;
		RECT	0.047 64.04 0.111 64.072 ;
		RECT	0.047 63.896 0.111 63.928 ;
		RECT	0.047 63.413 0.111 63.445 ;
		RECT	0.756 63.139 0.788 63.203 ;
		RECT	0.047 62.769 0.111 62.801 ;
		RECT	0.047 62.552 0.111 62.584 ;
		RECT	0.047 62.36 0.111 62.392 ;
		RECT	0.047 65.96 0.111 65.992 ;
		RECT	0.047 65.816 0.111 65.848 ;
		RECT	0.047 65.333 0.111 65.365 ;
		RECT	0.756 65.059 0.788 65.123 ;
		RECT	0.047 64.689 0.111 64.721 ;
		RECT	0.047 64.472 0.111 64.504 ;
		RECT	0.047 64.28 0.111 64.312 ;
		RECT	0.047 67.88 0.111 67.912 ;
		RECT	0.047 67.736 0.111 67.768 ;
		RECT	0.047 67.253 0.111 67.285 ;
		RECT	0.756 66.979 0.788 67.043 ;
		RECT	0.047 66.609 0.111 66.641 ;
		RECT	0.047 66.392 0.111 66.424 ;
		RECT	0.047 66.2 0.111 66.232 ;
		RECT	0.047 69.8 0.111 69.832 ;
		RECT	0.047 69.656 0.111 69.688 ;
		RECT	0.047 69.173 0.111 69.205 ;
		RECT	0.756 68.899 0.788 68.963 ;
		RECT	0.047 68.529 0.111 68.561 ;
		RECT	0.047 68.312 0.111 68.344 ;
		RECT	0.047 68.12 0.111 68.152 ;
		RECT	0.047 52.52 0.111 52.552 ;
		RECT	0.047 52.376 0.111 52.408 ;
		RECT	0.047 51.893 0.111 51.925 ;
		RECT	0.756 51.619 0.788 51.683 ;
		RECT	0.047 51.249 0.111 51.281 ;
		RECT	0.047 51.032 0.111 51.064 ;
		RECT	0.047 50.84 0.111 50.872 ;
		RECT	0.047 81.32 0.111 81.352 ;
		RECT	0.047 81.176 0.111 81.208 ;
		RECT	0.047 80.693 0.111 80.725 ;
		RECT	0.756 80.419 0.788 80.483 ;
		RECT	0.047 80.049 0.111 80.081 ;
		RECT	0.047 79.832 0.111 79.864 ;
		RECT	0.047 79.64 0.111 79.672 ;
		RECT	0.047 81.896 0.111 81.928 ;
		RECT	0.047 81.704 0.111 81.736 ;
		RECT	2.339 32.691 2.371 32.755 ;
		RECT	3.755 32.691 3.787 32.755 ;
		RECT	3.049 32.876 3.081 32.94 ;
		RECT	1.517 32.89 1.549 32.922 ;
		RECT	1.645 33.696 1.709 33.728 ;
		RECT	2.124 33.696 2.156 33.728 ;
		RECT	3.438 33.696 3.47 33.728 ;
		RECT	4.195 33.696 4.227 33.728 ;
		RECT	4.944 33.696 5.008 33.728 ;
		RECT	2.954 33.796 2.986 33.828 ;
		RECT	4.035 33.796 4.067 33.828 ;
		RECT	4.623 34.801 4.655 34.833 ;
		RECT	4.805 34.801 4.837 34.833 ;
		RECT	3.356 34.896 3.388 34.928 ;
		RECT	4.19 34.896 4.222 34.928 ;
		RECT	4.056 35.236 4.088 35.268 ;
		RECT	3.181 35.741 3.213 35.773 ;
		RECT	3.181 35.948 3.213 35.98 ;
		RECT	4.558 35.948 4.59 35.98 ;
		RECT	3.355 36.238 3.387 36.27 ;
		RECT	4.129 36.238 4.161 36.27 ;
		RECT	2.197 36.338 2.229 36.37 ;
		RECT	5.051 36.338 5.083 36.37 ;
		RECT	3.181 37.474 3.213 37.506 ;
		RECT	4.425 37.474 4.457 37.506 ;
		RECT	4.74 37.474 4.772 37.506 ;
		RECT	3.719 37.589 3.751 37.621 ;
		RECT	5.068 37.589 5.1 37.621 ;
		RECT	3.181 37.689 3.213 37.721 ;
		RECT	4.425 37.689 4.457 37.721 ;
		RECT	3.355 38.361 3.387 38.393 ;
		RECT	4.12 38.361 4.152 38.393 ;
		RECT	3.19 38.651 3.222 38.683 ;
		RECT	4.419 38.651 4.451 38.683 ;
		RECT	2.197 39.202 2.229 39.266 ;
		RECT	2.339 39.202 2.371 39.266 ;
		RECT	3.289 39.202 3.353 39.266 ;
		RECT	4.354 39.202 4.386 39.266 ;
		RECT	2.197 39.42 2.229 39.484 ;
		RECT	2.339 39.42 2.371 39.484 ;
		RECT	3.289 39.42 3.353 39.484 ;
		RECT	4.139 39.42 4.171 39.484 ;
		RECT	4.354 39.42 4.386 39.484 ;
		RECT	2.197 39.672 2.229 39.736 ;
		RECT	2.339 39.672 2.371 39.736 ;
		RECT	3.289 39.672 3.353 39.736 ;
		RECT	4.139 39.672 4.171 39.736 ;
		RECT	4.354 39.672 4.386 39.736 ;
		RECT	1.661 39.858 1.693 39.89 ;
		RECT	3.438 39.858 3.47 39.89 ;
		RECT	4.52 39.858 4.584 39.89 ;
		RECT	3.181 40.363 3.213 40.395 ;
		RECT	4.196 40.363 4.228 40.395 ;
		RECT	4.623 40.458 4.655 40.49 ;
		RECT	4.805 40.458 4.837 40.49 ;
		RECT	4.056 40.538 4.088 40.57 ;
		RECT	4.282 40.538 4.314 40.57 ;
		RECT	4.485 40.618 4.517 40.65 ;
		RECT	4.675 40.618 4.707 40.65 ;
		RECT	3.181 40.903 3.213 40.935 ;
		RECT	4.281 40.903 4.313 40.935 ;
		RECT	3.247 41.004 3.279 41.036 ;
		RECT	4.122 41.004 4.154 41.036 ;
		RECT	2.127 41.53 2.159 41.562 ;
		RECT	4.056 41.97 4.088 42.002 ;
		RECT	4.428 41.97 4.46 42.002 ;
		RECT	4.982 42.525 5.014 42.557 ;
		RECT	2.345 42.835 2.377 42.899 ;
		RECT	2.197 42.851 2.229 42.883 ;
		RECT	4.354 42.851 4.386 42.883 ;
		RECT	2.345 43.069 2.377 43.133 ;
		RECT	2.197 43.085 2.229 43.117 ;
		RECT	4.354 43.085 4.386 43.117 ;
		RECT	1.661 43.433 1.693 43.497 ;
		RECT	3.451 43.433 3.483 43.497 ;
		RECT	4.61 43.433 4.642 43.497 ;
		RECT	4.805 43.433 4.837 43.497 ;
		RECT	2.339 44.026 2.371 44.09 ;
		RECT	4.354 44.026 4.386 44.09 ;
		RECT	3.18 44.199 3.212 44.231 ;
		RECT	4.061 44.199 4.093 44.231 ;
		RECT	3.246 44.469 3.278 44.501 ;
		RECT	4.277 44.469 4.309 44.501 ;
		RECT	3.18 44.759 3.212 44.791 ;
		RECT	4.21 44.759 4.242 44.791 ;
		RECT	3.075 46.057 3.107 46.089 ;
		RECT	4.061 46.057 4.093 46.089 ;
		RECT	1.981 46.157 2.013 46.189 ;
		RECT	4.49 46.157 4.522 46.189 ;
		RECT	2.323 46.248 2.387 46.28 ;
		RECT	4.351 46.248 4.383 46.28 ;
		RECT	2.045 47.367 2.077 47.399 ;
		RECT	2.323 47.367 2.387 47.399 ;
		RECT	4.354 47.367 4.386 47.399 ;
		RECT	4.895 47.367 4.927 47.399 ;
		RECT	1.965 49.28 1.997 49.312 ;
		RECT	3.699 49.28 3.731 49.312 ;
		RECT	4.8 49.28 4.832 49.312 ;
		RECT	3.081 2.939 3.113 2.971 ;
		RECT	2.029 3.479 2.093 3.511 ;
		RECT	3.585 3.613 3.617 3.677 ;
		RECT	4.72 3.613 4.752 3.677 ;
		RECT	2.323 3.629 2.387 3.661 ;
		RECT	3.723 3.779 3.755 3.811 ;
		RECT	3.167 3.884 3.199 3.916 ;
		RECT	3.333 3.994 3.365 4.026 ;
		RECT	3.792 4.099 3.824 4.131 ;
		RECT	3.081 20.219 3.113 20.251 ;
		RECT	2.029 20.759 2.093 20.791 ;
		RECT	3.585 20.893 3.617 20.957 ;
		RECT	4.72 20.893 4.752 20.957 ;
		RECT	2.323 20.909 2.387 20.941 ;
		RECT	3.723 21.059 3.755 21.091 ;
		RECT	3.167 21.164 3.199 21.196 ;
		RECT	3.333 21.274 3.365 21.306 ;
		RECT	3.792 21.379 3.824 21.411 ;
		RECT	3.081 22.139 3.113 22.171 ;
		RECT	2.029 22.679 2.093 22.711 ;
		RECT	3.585 22.813 3.617 22.877 ;
		RECT	4.72 22.813 4.752 22.877 ;
		RECT	2.323 22.829 2.387 22.861 ;
		RECT	3.723 22.979 3.755 23.011 ;
		RECT	3.167 23.084 3.199 23.116 ;
		RECT	3.333 23.194 3.365 23.226 ;
		RECT	3.792 23.299 3.824 23.331 ;
		RECT	3.081 24.059 3.113 24.091 ;
		RECT	2.029 24.599 2.093 24.631 ;
		RECT	3.585 24.733 3.617 24.797 ;
		RECT	4.72 24.733 4.752 24.797 ;
		RECT	2.323 24.749 2.387 24.781 ;
		RECT	3.723 24.899 3.755 24.931 ;
		RECT	3.167 25.004 3.199 25.036 ;
		RECT	3.333 25.114 3.365 25.146 ;
		RECT	3.792 25.219 3.824 25.251 ;
		RECT	3.081 25.979 3.113 26.011 ;
		RECT	2.029 26.519 2.093 26.551 ;
		RECT	3.585 26.653 3.617 26.717 ;
		RECT	4.72 26.653 4.752 26.717 ;
		RECT	2.323 26.669 2.387 26.701 ;
		RECT	3.723 26.819 3.755 26.851 ;
		RECT	3.167 26.924 3.199 26.956 ;
		RECT	3.333 27.034 3.365 27.066 ;
		RECT	3.792 27.139 3.824 27.171 ;
		RECT	3.081 27.899 3.113 27.931 ;
		RECT	2.029 28.439 2.093 28.471 ;
		RECT	3.585 28.573 3.617 28.637 ;
		RECT	4.72 28.573 4.752 28.637 ;
		RECT	2.323 28.589 2.387 28.621 ;
		RECT	3.723 28.739 3.755 28.771 ;
		RECT	3.167 28.844 3.199 28.876 ;
		RECT	3.333 28.954 3.365 28.986 ;
		RECT	3.792 29.059 3.824 29.091 ;
		RECT	3.081 4.859 3.113 4.891 ;
		RECT	2.029 5.399 2.093 5.431 ;
		RECT	3.585 5.533 3.617 5.597 ;
		RECT	4.72 5.533 4.752 5.597 ;
		RECT	2.323 5.549 2.387 5.581 ;
		RECT	3.723 5.699 3.755 5.731 ;
		RECT	3.167 5.804 3.199 5.836 ;
		RECT	3.333 5.914 3.365 5.946 ;
		RECT	3.792 6.019 3.824 6.051 ;
		RECT	3.081 6.779 3.113 6.811 ;
		RECT	2.029 7.319 2.093 7.351 ;
		RECT	3.585 7.453 3.617 7.517 ;
		RECT	4.72 7.453 4.752 7.517 ;
		RECT	2.323 7.469 2.387 7.501 ;
		RECT	3.723 7.619 3.755 7.651 ;
		RECT	3.167 7.724 3.199 7.756 ;
		RECT	3.333 7.834 3.365 7.866 ;
		RECT	3.792 7.939 3.824 7.971 ;
		RECT	3.081 8.699 3.113 8.731 ;
		RECT	2.029 9.239 2.093 9.271 ;
		RECT	3.585 9.373 3.617 9.437 ;
		RECT	4.72 9.373 4.752 9.437 ;
		RECT	2.323 9.389 2.387 9.421 ;
		RECT	3.723 9.539 3.755 9.571 ;
		RECT	3.167 9.644 3.199 9.676 ;
		RECT	3.333 9.754 3.365 9.786 ;
		RECT	3.792 9.859 3.824 9.891 ;
		RECT	3.081 10.619 3.113 10.651 ;
		RECT	2.029 11.159 2.093 11.191 ;
		RECT	3.585 11.293 3.617 11.357 ;
		RECT	4.72 11.293 4.752 11.357 ;
		RECT	2.323 11.309 2.387 11.341 ;
		RECT	3.723 11.459 3.755 11.491 ;
		RECT	3.167 11.564 3.199 11.596 ;
		RECT	3.333 11.674 3.365 11.706 ;
		RECT	3.792 11.779 3.824 11.811 ;
		RECT	3.081 12.539 3.113 12.571 ;
		RECT	2.029 13.079 2.093 13.111 ;
		RECT	3.585 13.213 3.617 13.277 ;
		RECT	4.72 13.213 4.752 13.277 ;
		RECT	2.323 13.229 2.387 13.261 ;
		RECT	3.723 13.379 3.755 13.411 ;
		RECT	3.167 13.484 3.199 13.516 ;
		RECT	3.333 13.594 3.365 13.626 ;
		RECT	3.792 13.699 3.824 13.731 ;
		RECT	3.081 14.459 3.113 14.491 ;
		RECT	2.029 14.999 2.093 15.031 ;
		RECT	3.585 15.133 3.617 15.197 ;
		RECT	4.72 15.133 4.752 15.197 ;
		RECT	2.323 15.149 2.387 15.181 ;
		RECT	3.723 15.299 3.755 15.331 ;
		RECT	3.167 15.404 3.199 15.436 ;
		RECT	3.333 15.514 3.365 15.546 ;
		RECT	3.792 15.619 3.824 15.651 ;
		RECT	3.081 16.379 3.113 16.411 ;
		RECT	2.029 16.919 2.093 16.951 ;
		RECT	3.585 17.053 3.617 17.117 ;
		RECT	4.72 17.053 4.752 17.117 ;
		RECT	2.323 17.069 2.387 17.101 ;
		RECT	3.723 17.219 3.755 17.251 ;
		RECT	3.167 17.324 3.199 17.356 ;
		RECT	3.333 17.434 3.365 17.466 ;
		RECT	3.792 17.539 3.824 17.571 ;
		RECT	3.081 18.299 3.113 18.331 ;
		RECT	2.029 18.839 2.093 18.871 ;
		RECT	3.585 18.973 3.617 19.037 ;
		RECT	4.72 18.973 4.752 19.037 ;
		RECT	2.323 18.989 2.387 19.021 ;
		RECT	3.723 19.139 3.755 19.171 ;
		RECT	3.167 19.244 3.199 19.276 ;
		RECT	3.333 19.354 3.365 19.386 ;
		RECT	3.792 19.459 3.824 19.491 ;
		RECT	3.081 1.019 3.113 1.051 ;
		RECT	2.029 1.559 2.093 1.591 ;
		RECT	3.585 1.693 3.617 1.757 ;
		RECT	4.72 1.693 4.752 1.757 ;
		RECT	2.323 1.709 2.387 1.741 ;
		RECT	3.723 1.859 3.755 1.891 ;
		RECT	3.167 1.964 3.199 1.996 ;
		RECT	3.333 2.074 3.365 2.106 ;
		RECT	3.792 2.179 3.824 2.211 ;
		RECT	3.081 29.819 3.113 29.851 ;
		RECT	2.029 30.359 2.093 30.391 ;
		RECT	3.585 30.493 3.617 30.557 ;
		RECT	4.72 30.493 4.752 30.557 ;
		RECT	2.323 30.509 2.387 30.541 ;
		RECT	3.723 30.659 3.755 30.691 ;
		RECT	3.167 30.764 3.199 30.796 ;
		RECT	3.333 30.874 3.365 30.906 ;
		RECT	3.792 30.979 3.824 31.011 ;
		RECT	5.064 45.197 5.096 45.229 ;
		RECT	3.922 51.485 3.954 51.517 ;
		RECT	3.922 51.165 3.954 51.197 ;
		RECT	3.922 1.859 3.954 1.891 ;
		RECT	3.922 2.179 3.954 2.211 ;
		RECT	3.922 21.059 3.954 21.091 ;
		RECT	3.922 21.379 3.954 21.411 ;
		RECT	3.922 70.685 3.954 70.717 ;
		RECT	3.922 70.365 3.954 70.397 ;
		RECT	3.922 22.979 3.954 23.011 ;
		RECT	3.922 23.299 3.954 23.331 ;
		RECT	3.922 72.605 3.954 72.637 ;
		RECT	3.922 72.285 3.954 72.317 ;
		RECT	3.922 24.899 3.954 24.931 ;
		RECT	3.922 25.219 3.954 25.251 ;
		RECT	3.922 74.525 3.954 74.557 ;
		RECT	3.922 74.205 3.954 74.237 ;
		RECT	3.922 26.819 3.954 26.851 ;
		RECT	3.922 27.139 3.954 27.171 ;
		RECT	3.922 76.445 3.954 76.477 ;
		RECT	3.922 76.125 3.954 76.157 ;
		RECT	3.922 28.739 3.954 28.771 ;
		RECT	3.922 29.059 3.954 29.091 ;
		RECT	3.922 78.365 3.954 78.397 ;
		RECT	3.922 78.045 3.954 78.077 ;
		RECT	3.922 30.659 3.954 30.691 ;
		RECT	3.922 30.979 3.954 31.011 ;
		RECT	3.922 80.285 3.954 80.317 ;
		RECT	3.922 79.965 3.954 79.997 ;
		RECT	3.922 53.405 3.954 53.437 ;
		RECT	3.922 53.085 3.954 53.117 ;
		RECT	3.922 3.779 3.954 3.811 ;
		RECT	3.922 4.099 3.954 4.131 ;
		RECT	3.922 55.325 3.954 55.357 ;
		RECT	3.922 55.005 3.954 55.037 ;
		RECT	3.922 5.699 3.954 5.731 ;
		RECT	3.922 6.019 3.954 6.051 ;
		RECT	3.922 57.245 3.954 57.277 ;
		RECT	3.922 56.925 3.954 56.957 ;
		RECT	3.922 7.619 3.954 7.651 ;
		RECT	3.922 7.939 3.954 7.971 ;
		RECT	3.922 59.165 3.954 59.197 ;
		RECT	3.922 58.845 3.954 58.877 ;
		RECT	3.922 9.539 3.954 9.571 ;
		RECT	3.922 9.859 3.954 9.891 ;
		RECT	3.922 61.085 3.954 61.117 ;
		RECT	3.922 60.765 3.954 60.797 ;
		RECT	3.922 11.459 3.954 11.491 ;
		RECT	3.922 11.779 3.954 11.811 ;
		RECT	3.922 63.005 3.954 63.037 ;
		RECT	3.922 62.685 3.954 62.717 ;
		RECT	3.922 13.379 3.954 13.411 ;
		RECT	3.922 13.699 3.954 13.731 ;
		RECT	3.922 64.925 3.954 64.957 ;
		RECT	3.922 64.605 3.954 64.637 ;
		RECT	3.922 15.299 3.954 15.331 ;
		RECT	3.922 15.619 3.954 15.651 ;
		RECT	3.922 17.219 3.954 17.251 ;
		RECT	3.922 17.539 3.954 17.571 ;
		RECT	3.922 66.845 3.954 66.877 ;
		RECT	3.922 66.525 3.954 66.557 ;
		RECT	3.922 19.139 3.954 19.171 ;
		RECT	3.922 19.459 3.954 19.491 ;
		RECT	3.922 68.765 3.954 68.797 ;
		RECT	3.922 68.445 3.954 68.477 ;
		RECT	3.382 41.87 3.414 41.902 ;
		RECT	3.081 54.245 3.113 54.277 ;
		RECT	2.029 53.705 2.093 53.737 ;
		RECT	3.585 53.539 3.617 53.603 ;
		RECT	4.72 53.539 4.752 53.603 ;
		RECT	2.323 53.555 2.387 53.587 ;
		RECT	3.723 53.405 3.755 53.437 ;
		RECT	3.167 53.3 3.199 53.332 ;
		RECT	3.333 53.19 3.365 53.222 ;
		RECT	3.792 53.085 3.824 53.117 ;
		RECT	3.081 71.525 3.113 71.557 ;
		RECT	2.029 70.985 2.093 71.017 ;
		RECT	3.585 70.819 3.617 70.883 ;
		RECT	4.72 70.819 4.752 70.883 ;
		RECT	2.323 70.835 2.387 70.867 ;
		RECT	3.723 70.685 3.755 70.717 ;
		RECT	3.167 70.58 3.199 70.612 ;
		RECT	3.333 70.47 3.365 70.502 ;
		RECT	3.792 70.365 3.824 70.397 ;
		RECT	3.081 73.445 3.113 73.477 ;
		RECT	2.029 72.905 2.093 72.937 ;
		RECT	3.585 72.739 3.617 72.803 ;
		RECT	4.72 72.739 4.752 72.803 ;
		RECT	2.323 72.755 2.387 72.787 ;
		RECT	3.723 72.605 3.755 72.637 ;
		RECT	3.167 72.5 3.199 72.532 ;
		RECT	3.333 72.39 3.365 72.422 ;
		RECT	3.792 72.285 3.824 72.317 ;
		RECT	3.081 75.365 3.113 75.397 ;
		RECT	2.029 74.825 2.093 74.857 ;
		RECT	3.585 74.659 3.617 74.723 ;
		RECT	4.72 74.659 4.752 74.723 ;
		RECT	2.323 74.675 2.387 74.707 ;
		RECT	3.723 74.525 3.755 74.557 ;
		RECT	3.167 74.42 3.199 74.452 ;
		RECT	3.333 74.31 3.365 74.342 ;
		RECT	3.792 74.205 3.824 74.237 ;
		RECT	3.081 77.285 3.113 77.317 ;
		RECT	2.029 76.745 2.093 76.777 ;
		RECT	3.585 76.579 3.617 76.643 ;
		RECT	4.72 76.579 4.752 76.643 ;
		RECT	2.323 76.595 2.387 76.627 ;
		RECT	3.723 76.445 3.755 76.477 ;
		RECT	3.167 76.34 3.199 76.372 ;
		RECT	3.333 76.23 3.365 76.262 ;
		RECT	3.792 76.125 3.824 76.157 ;
		RECT	3.081 79.205 3.113 79.237 ;
		RECT	2.029 78.665 2.093 78.697 ;
		RECT	3.585 78.499 3.617 78.563 ;
		RECT	4.72 78.499 4.752 78.563 ;
		RECT	2.323 78.515 2.387 78.547 ;
		RECT	3.723 78.365 3.755 78.397 ;
		RECT	3.167 78.26 3.199 78.292 ;
		RECT	3.333 78.15 3.365 78.182 ;
		RECT	3.792 78.045 3.824 78.077 ;
		RECT	3.081 56.165 3.113 56.197 ;
		RECT	2.029 55.625 2.093 55.657 ;
		RECT	3.585 55.459 3.617 55.523 ;
		RECT	4.72 55.459 4.752 55.523 ;
		RECT	2.323 55.475 2.387 55.507 ;
		RECT	3.723 55.325 3.755 55.357 ;
		RECT	3.167 55.22 3.199 55.252 ;
		RECT	3.333 55.11 3.365 55.142 ;
		RECT	3.792 55.005 3.824 55.037 ;
		RECT	3.081 58.085 3.113 58.117 ;
		RECT	2.029 57.545 2.093 57.577 ;
		RECT	3.585 57.379 3.617 57.443 ;
		RECT	4.72 57.379 4.752 57.443 ;
		RECT	2.323 57.395 2.387 57.427 ;
		RECT	3.723 57.245 3.755 57.277 ;
		RECT	3.167 57.14 3.199 57.172 ;
		RECT	3.333 57.03 3.365 57.062 ;
		RECT	3.792 56.925 3.824 56.957 ;
		RECT	3.081 60.005 3.113 60.037 ;
		RECT	2.029 59.465 2.093 59.497 ;
		RECT	3.585 59.299 3.617 59.363 ;
		RECT	4.72 59.299 4.752 59.363 ;
		RECT	2.323 59.315 2.387 59.347 ;
		RECT	3.723 59.165 3.755 59.197 ;
		RECT	3.167 59.06 3.199 59.092 ;
		RECT	3.333 58.95 3.365 58.982 ;
		RECT	3.792 58.845 3.824 58.877 ;
		RECT	3.081 61.925 3.113 61.957 ;
		RECT	2.029 61.385 2.093 61.417 ;
		RECT	3.585 61.219 3.617 61.283 ;
		RECT	4.72 61.219 4.752 61.283 ;
		RECT	2.323 61.235 2.387 61.267 ;
		RECT	3.723 61.085 3.755 61.117 ;
		RECT	3.167 60.98 3.199 61.012 ;
		RECT	3.333 60.87 3.365 60.902 ;
		RECT	3.792 60.765 3.824 60.797 ;
		RECT	3.081 63.845 3.113 63.877 ;
		RECT	2.029 63.305 2.093 63.337 ;
		RECT	3.585 63.139 3.617 63.203 ;
		RECT	4.72 63.139 4.752 63.203 ;
		RECT	2.323 63.155 2.387 63.187 ;
		RECT	3.723 63.005 3.755 63.037 ;
		RECT	3.167 62.9 3.199 62.932 ;
		RECT	3.333 62.79 3.365 62.822 ;
		RECT	3.792 62.685 3.824 62.717 ;
		RECT	3.081 65.765 3.113 65.797 ;
		RECT	2.029 65.225 2.093 65.257 ;
		RECT	3.585 65.059 3.617 65.123 ;
		RECT	4.72 65.059 4.752 65.123 ;
		RECT	2.323 65.075 2.387 65.107 ;
		RECT	3.723 64.925 3.755 64.957 ;
		RECT	3.167 64.82 3.199 64.852 ;
		RECT	3.333 64.71 3.365 64.742 ;
		RECT	3.792 64.605 3.824 64.637 ;
		RECT	3.081 67.685 3.113 67.717 ;
		RECT	2.029 67.145 2.093 67.177 ;
		RECT	3.585 66.979 3.617 67.043 ;
		RECT	4.72 66.979 4.752 67.043 ;
		RECT	2.323 66.995 2.387 67.027 ;
		RECT	3.723 66.845 3.755 66.877 ;
		RECT	3.167 66.74 3.199 66.772 ;
		RECT	3.333 66.63 3.365 66.662 ;
		RECT	3.792 66.525 3.824 66.557 ;
		RECT	3.081 69.605 3.113 69.637 ;
		RECT	2.029 69.065 2.093 69.097 ;
		RECT	3.585 68.899 3.617 68.963 ;
		RECT	4.72 68.899 4.752 68.963 ;
		RECT	2.323 68.915 2.387 68.947 ;
		RECT	3.723 68.765 3.755 68.797 ;
		RECT	3.167 68.66 3.199 68.692 ;
		RECT	3.333 68.55 3.365 68.582 ;
		RECT	3.792 68.445 3.824 68.477 ;
		RECT	3.081 52.325 3.113 52.357 ;
		RECT	2.029 51.785 2.093 51.817 ;
		RECT	3.585 51.619 3.617 51.683 ;
		RECT	4.72 51.619 4.752 51.683 ;
		RECT	2.323 51.635 2.387 51.667 ;
		RECT	3.723 51.485 3.755 51.517 ;
		RECT	3.167 51.38 3.199 51.412 ;
		RECT	3.333 51.27 3.365 51.302 ;
		RECT	3.792 51.165 3.824 51.197 ;
		RECT	3.081 81.125 3.113 81.157 ;
		RECT	2.029 80.585 2.093 80.617 ;
		RECT	3.585 80.419 3.617 80.483 ;
		RECT	4.72 80.419 4.752 80.483 ;
		RECT	2.323 80.435 2.387 80.467 ;
		RECT	3.723 80.285 3.755 80.317 ;
		RECT	3.167 80.18 3.199 80.212 ;
		RECT	3.333 80.07 3.365 80.102 ;
		RECT	3.792 79.965 3.824 79.997 ;
		RECT	4.944 51.485 5.008 51.517 ;
		RECT	4.944 51.165 5.008 51.197 ;
		RECT	4.944 1.859 5.008 1.891 ;
		RECT	4.944 2.179 5.008 2.211 ;
		RECT	4.944 21.059 5.008 21.091 ;
		RECT	4.944 21.379 5.008 21.411 ;
		RECT	4.944 70.685 5.008 70.717 ;
		RECT	4.944 70.365 5.008 70.397 ;
		RECT	4.944 22.979 5.008 23.011 ;
		RECT	4.944 23.299 5.008 23.331 ;
		RECT	4.944 72.605 5.008 72.637 ;
		RECT	4.944 72.285 5.008 72.317 ;
		RECT	4.944 24.899 5.008 24.931 ;
		RECT	4.944 25.219 5.008 25.251 ;
		RECT	4.944 74.525 5.008 74.557 ;
		RECT	4.944 74.205 5.008 74.237 ;
		RECT	4.944 26.819 5.008 26.851 ;
		RECT	4.944 27.139 5.008 27.171 ;
		RECT	4.944 76.445 5.008 76.477 ;
		RECT	4.944 76.125 5.008 76.157 ;
		RECT	4.944 28.739 5.008 28.771 ;
		RECT	4.944 29.059 5.008 29.091 ;
		RECT	4.944 78.365 5.008 78.397 ;
		RECT	4.944 78.045 5.008 78.077 ;
		RECT	4.944 30.659 5.008 30.691 ;
		RECT	4.944 30.979 5.008 31.011 ;
		RECT	4.944 80.285 5.008 80.317 ;
		RECT	4.944 79.965 5.008 79.997 ;
		RECT	4.944 53.405 5.008 53.437 ;
		RECT	4.944 53.085 5.008 53.117 ;
		RECT	4.944 3.779 5.008 3.811 ;
		RECT	4.944 4.099 5.008 4.131 ;
		RECT	4.944 55.325 5.008 55.357 ;
		RECT	4.944 55.005 5.008 55.037 ;
		RECT	4.944 5.699 5.008 5.731 ;
		RECT	4.944 6.019 5.008 6.051 ;
		RECT	4.944 57.245 5.008 57.277 ;
		RECT	4.944 56.925 5.008 56.957 ;
		RECT	4.944 7.619 5.008 7.651 ;
		RECT	4.944 7.939 5.008 7.971 ;
		RECT	4.944 59.165 5.008 59.197 ;
		RECT	4.944 58.845 5.008 58.877 ;
		RECT	4.944 9.539 5.008 9.571 ;
		RECT	4.944 9.859 5.008 9.891 ;
		RECT	4.944 61.085 5.008 61.117 ;
		RECT	4.944 60.765 5.008 60.797 ;
		RECT	4.944 11.459 5.008 11.491 ;
		RECT	4.944 11.779 5.008 11.811 ;
		RECT	4.944 63.005 5.008 63.037 ;
		RECT	4.944 62.685 5.008 62.717 ;
		RECT	4.944 13.379 5.008 13.411 ;
		RECT	4.944 13.699 5.008 13.731 ;
		RECT	4.944 64.925 5.008 64.957 ;
		RECT	4.944 64.605 5.008 64.637 ;
		RECT	4.944 15.299 5.008 15.331 ;
		RECT	4.944 15.619 5.008 15.651 ;
		RECT	4.944 17.219 5.008 17.251 ;
		RECT	4.944 17.539 5.008 17.571 ;
		RECT	4.944 66.845 5.008 66.877 ;
		RECT	4.944 66.525 5.008 66.557 ;
		RECT	4.944 19.139 5.008 19.171 ;
		RECT	4.944 19.459 5.008 19.491 ;
		RECT	4.944 68.765 5.008 68.797 ;
		RECT	4.944 68.445 5.008 68.477 ;
		RECT	1.645 1.709 1.709 1.741 ;
		RECT	3.438 1.693 3.47 1.757 ;
		RECT	4.195 1.693 4.227 1.757 ;
		RECT	4.944 1.709 5.008 1.741 ;
		RECT	1.645 51.635 1.709 51.667 ;
		RECT	3.438 51.619 3.47 51.683 ;
		RECT	4.195 51.619 4.227 51.683 ;
		RECT	4.944 51.635 5.008 51.667 ;
		RECT	1.645 32.691 1.709 32.755 ;
		RECT	3.438 32.691 3.47 32.755 ;
		RECT	4.195 32.691 4.227 32.755 ;
		RECT	4.944 32.691 5.008 32.755 ;
		RECT	2.323 33.696 2.387 33.728 ;
		RECT	4.536 39.202 4.568 39.266 ;
		RECT	4.536 39.42 4.568 39.484 ;
		RECT	4.536 39.672 4.568 39.736 ;
		RECT	1.645 42.835 1.709 42.899 ;
		RECT	3.451 42.835 3.483 42.899 ;
		RECT	4.805 42.835 4.837 42.899 ;
		RECT	1.645 43.069 1.709 43.133 ;
		RECT	3.451 43.069 3.483 43.133 ;
		RECT	4.61 43.069 4.642 43.133 ;
		RECT	4.805 43.069 4.837 43.133 ;
		RECT	1.645 44.042 1.709 44.074 ;
		RECT	3.451 44.026 3.483 44.09 ;
		RECT	4.805 44.026 4.837 44.09 ;
		RECT	3.451 46.248 3.483 46.28 ;
		RECT	1.645 20.909 1.709 20.941 ;
		RECT	3.438 20.893 3.47 20.957 ;
		RECT	4.195 20.893 4.227 20.957 ;
		RECT	4.944 20.909 5.008 20.941 ;
		RECT	1.645 70.835 1.709 70.867 ;
		RECT	3.438 70.819 3.47 70.883 ;
		RECT	4.195 70.819 4.227 70.883 ;
		RECT	4.944 70.835 5.008 70.867 ;
		RECT	1.645 22.829 1.709 22.861 ;
		RECT	3.438 22.813 3.47 22.877 ;
		RECT	4.195 22.813 4.227 22.877 ;
		RECT	4.944 22.829 5.008 22.861 ;
		RECT	1.645 72.755 1.709 72.787 ;
		RECT	3.438 72.739 3.47 72.803 ;
		RECT	4.195 72.739 4.227 72.803 ;
		RECT	4.944 72.755 5.008 72.787 ;
		RECT	1.645 24.749 1.709 24.781 ;
		RECT	3.438 24.733 3.47 24.797 ;
		RECT	4.195 24.733 4.227 24.797 ;
		RECT	4.944 24.749 5.008 24.781 ;
		RECT	1.645 74.675 1.709 74.707 ;
		RECT	3.438 74.659 3.47 74.723 ;
		RECT	4.195 74.659 4.227 74.723 ;
		RECT	4.944 74.675 5.008 74.707 ;
		RECT	1.645 26.669 1.709 26.701 ;
		RECT	3.438 26.653 3.47 26.717 ;
		RECT	4.195 26.653 4.227 26.717 ;
		RECT	4.944 26.669 5.008 26.701 ;
		RECT	1.645 76.595 1.709 76.627 ;
		RECT	3.438 76.579 3.47 76.643 ;
		RECT	4.195 76.579 4.227 76.643 ;
		RECT	4.944 76.595 5.008 76.627 ;
		RECT	1.645 28.589 1.709 28.621 ;
		RECT	3.438 28.573 3.47 28.637 ;
		RECT	4.195 28.573 4.227 28.637 ;
		RECT	4.944 28.589 5.008 28.621 ;
		RECT	1.645 78.515 1.709 78.547 ;
		RECT	3.438 78.499 3.47 78.563 ;
		RECT	4.195 78.499 4.227 78.563 ;
		RECT	4.944 78.515 5.008 78.547 ;
		RECT	1.645 30.509 1.709 30.541 ;
		RECT	3.438 30.493 3.47 30.557 ;
		RECT	4.195 30.493 4.227 30.557 ;
		RECT	4.944 30.509 5.008 30.541 ;
		RECT	1.645 80.435 1.709 80.467 ;
		RECT	3.438 80.419 3.47 80.483 ;
		RECT	4.195 80.419 4.227 80.483 ;
		RECT	4.944 80.435 5.008 80.467 ;
		RECT	1.645 3.629 1.709 3.661 ;
		RECT	3.438 3.613 3.47 3.677 ;
		RECT	4.195 3.613 4.227 3.677 ;
		RECT	4.944 3.629 5.008 3.661 ;
		RECT	1.645 53.555 1.709 53.587 ;
		RECT	3.438 53.539 3.47 53.603 ;
		RECT	4.195 53.539 4.227 53.603 ;
		RECT	4.944 53.555 5.008 53.587 ;
		RECT	1.645 5.549 1.709 5.581 ;
		RECT	3.438 5.533 3.47 5.597 ;
		RECT	4.195 5.533 4.227 5.597 ;
		RECT	4.944 5.549 5.008 5.581 ;
		RECT	1.645 55.475 1.709 55.507 ;
		RECT	3.438 55.459 3.47 55.523 ;
		RECT	4.195 55.459 4.227 55.523 ;
		RECT	4.944 55.475 5.008 55.507 ;
		RECT	1.645 7.469 1.709 7.501 ;
		RECT	3.438 7.453 3.47 7.517 ;
		RECT	4.195 7.453 4.227 7.517 ;
		RECT	4.944 7.469 5.008 7.501 ;
		RECT	1.645 57.395 1.709 57.427 ;
		RECT	3.438 57.379 3.47 57.443 ;
		RECT	4.195 57.379 4.227 57.443 ;
		RECT	4.944 57.395 5.008 57.427 ;
		RECT	1.645 9.389 1.709 9.421 ;
		RECT	3.438 9.373 3.47 9.437 ;
		RECT	4.195 9.373 4.227 9.437 ;
		RECT	4.944 9.389 5.008 9.421 ;
		RECT	1.645 59.315 1.709 59.347 ;
		RECT	3.438 59.299 3.47 59.363 ;
		RECT	4.195 59.299 4.227 59.363 ;
		RECT	4.944 59.315 5.008 59.347 ;
		RECT	1.645 11.309 1.709 11.341 ;
		RECT	3.438 11.293 3.47 11.357 ;
		RECT	4.195 11.293 4.227 11.357 ;
		RECT	4.944 11.309 5.008 11.341 ;
		RECT	1.645 61.235 1.709 61.267 ;
		RECT	3.438 61.219 3.47 61.283 ;
		RECT	4.195 61.219 4.227 61.283 ;
		RECT	4.944 61.235 5.008 61.267 ;
		RECT	1.645 13.229 1.709 13.261 ;
		RECT	3.438 13.213 3.47 13.277 ;
		RECT	4.195 13.213 4.227 13.277 ;
		RECT	4.944 13.229 5.008 13.261 ;
		RECT	1.645 63.155 1.709 63.187 ;
		RECT	3.438 63.139 3.47 63.203 ;
		RECT	4.195 63.139 4.227 63.203 ;
		RECT	4.944 63.155 5.008 63.187 ;
		RECT	1.645 15.149 1.709 15.181 ;
		RECT	3.438 15.133 3.47 15.197 ;
		RECT	4.195 15.133 4.227 15.197 ;
		RECT	4.944 15.149 5.008 15.181 ;
		RECT	1.645 65.075 1.709 65.107 ;
		RECT	3.438 65.059 3.47 65.123 ;
		RECT	4.195 65.059 4.227 65.123 ;
		RECT	4.944 65.075 5.008 65.107 ;
		RECT	1.645 17.069 1.709 17.101 ;
		RECT	3.438 17.053 3.47 17.117 ;
		RECT	4.195 17.053 4.227 17.117 ;
		RECT	4.944 17.069 5.008 17.101 ;
		RECT	1.645 66.995 1.709 67.027 ;
		RECT	3.438 66.979 3.47 67.043 ;
		RECT	4.195 66.979 4.227 67.043 ;
		RECT	4.944 66.995 5.008 67.027 ;
		RECT	1.645 18.989 1.709 19.021 ;
		RECT	3.438 18.973 3.47 19.037 ;
		RECT	4.195 18.973 4.227 19.037 ;
		RECT	4.944 18.989 5.008 19.021 ;
		RECT	1.645 68.915 1.709 68.947 ;
		RECT	3.438 68.899 3.47 68.963 ;
		RECT	4.195 68.899 4.227 68.963 ;
		RECT	4.944 68.915 5.008 68.947 ;
		RECT	102.995 44.026 103.027 44.09 ;
		RECT	103.175 44.026 103.207 44.09 ;
		RECT	102.995 1.693 103.027 1.757 ;
		RECT	103.175 1.693 103.207 1.757 ;
		RECT	102.995 3.613 103.027 3.677 ;
		RECT	103.175 3.613 103.207 3.677 ;
		RECT	102.995 20.893 103.027 20.957 ;
		RECT	103.175 20.893 103.207 20.957 ;
		RECT	102.995 22.813 103.027 22.877 ;
		RECT	103.175 22.813 103.207 22.877 ;
		RECT	102.995 24.733 103.027 24.797 ;
		RECT	103.175 24.733 103.207 24.797 ;
		RECT	102.995 26.653 103.027 26.717 ;
		RECT	103.175 26.653 103.207 26.717 ;
		RECT	102.995 28.573 103.027 28.637 ;
		RECT	103.175 28.573 103.207 28.637 ;
		RECT	102.995 30.493 103.027 30.557 ;
		RECT	103.175 30.493 103.207 30.557 ;
		RECT	102.995 5.533 103.027 5.597 ;
		RECT	103.175 5.533 103.207 5.597 ;
		RECT	102.995 7.453 103.027 7.517 ;
		RECT	103.175 7.453 103.207 7.517 ;
		RECT	102.995 9.373 103.027 9.437 ;
		RECT	103.175 9.373 103.207 9.437 ;
		RECT	102.995 11.293 103.027 11.357 ;
		RECT	103.175 11.293 103.207 11.357 ;
		RECT	102.995 13.213 103.027 13.277 ;
		RECT	103.175 13.213 103.207 13.277 ;
		RECT	102.995 15.133 103.027 15.197 ;
		RECT	103.175 15.133 103.207 15.197 ;
		RECT	102.995 17.053 103.027 17.117 ;
		RECT	103.175 17.053 103.207 17.117 ;
		RECT	102.995 18.973 103.027 19.037 ;
		RECT	103.175 18.973 103.207 19.037 ;
		RECT	102.995 51.619 103.027 51.683 ;
		RECT	103.175 51.619 103.207 51.683 ;
		RECT	102.995 53.539 103.027 53.603 ;
		RECT	103.175 53.539 103.207 53.603 ;
		RECT	102.995 70.819 103.027 70.883 ;
		RECT	103.175 70.819 103.207 70.883 ;
		RECT	102.995 72.739 103.027 72.803 ;
		RECT	103.175 72.739 103.207 72.803 ;
		RECT	102.995 74.659 103.027 74.723 ;
		RECT	103.175 74.659 103.207 74.723 ;
		RECT	102.995 76.579 103.027 76.643 ;
		RECT	103.175 76.579 103.207 76.643 ;
		RECT	102.995 78.499 103.027 78.563 ;
		RECT	103.175 78.499 103.207 78.563 ;
		RECT	102.995 80.419 103.027 80.483 ;
		RECT	103.175 80.419 103.207 80.483 ;
		RECT	102.995 55.459 103.027 55.523 ;
		RECT	103.175 55.459 103.207 55.523 ;
		RECT	102.995 57.379 103.027 57.443 ;
		RECT	103.175 57.379 103.207 57.443 ;
		RECT	102.995 59.299 103.027 59.363 ;
		RECT	103.175 59.299 103.207 59.363 ;
		RECT	102.995 61.219 103.027 61.283 ;
		RECT	103.175 61.219 103.207 61.283 ;
		RECT	102.995 63.139 103.027 63.203 ;
		RECT	103.175 63.139 103.207 63.203 ;
		RECT	102.995 65.059 103.027 65.123 ;
		RECT	103.175 65.059 103.207 65.123 ;
		RECT	102.995 66.979 103.027 67.043 ;
		RECT	103.175 66.979 103.207 67.043 ;
		RECT	102.995 68.899 103.027 68.963 ;
		RECT	103.175 68.899 103.207 68.963 ;
		RECT	52.003 33.796 52.035 33.828 ;
		RECT	52.124 32.691 52.156 32.755 ;
		RECT	52.578 32.691 52.61 32.755 ;
		RECT	52.968 32.691 53.032 32.755 ;
		RECT	54.251 32.691 54.283 32.755 ;
		RECT	55.562 32.691 55.626 32.755 ;
		RECT	55.803 32.691 55.835 32.755 ;
		RECT	54.959 32.876 54.991 32.94 ;
		RECT	50.33 33.437 50.362 33.469 ;
		RECT	57.931 33.437 57.963 33.469 ;
		RECT	52.078 33.701 52.11 33.733 ;
		RECT	54.963 33.701 54.995 33.733 ;
		RECT	54.279 34.641 54.311 34.673 ;
		RECT	55.458 34.721 55.49 34.753 ;
		RECT	53.245 34.801 53.277 34.833 ;
		RECT	52.454 34.896 52.486 34.928 ;
		RECT	50.588 35.948 50.62 35.98 ;
		RECT	52.291 36.454 52.323 36.486 ;
		RECT	54.359 36.454 54.391 36.486 ;
		RECT	57.838 36.454 57.87 36.486 ;
		RECT	53.105 37.589 53.137 37.621 ;
		RECT	51.886 37.689 51.918 37.721 ;
		RECT	52.15 38.361 52.182 38.393 ;
		RECT	53.104 38.651 53.136 38.683 ;
		RECT	51.92 39.191 51.952 39.255 ;
		RECT	50.417 39.192 50.481 39.256 ;
		RECT	51.274 39.192 51.306 39.256 ;
		RECT	53.91 39.192 53.942 39.256 ;
		RECT	54.363 39.192 54.427 39.256 ;
		RECT	54.812 39.192 54.844 39.256 ;
		RECT	55.208 39.192 55.272 39.256 ;
		RECT	55.562 39.192 55.626 39.256 ;
		RECT	55.969 39.192 56.033 39.256 ;
		RECT	57.363 39.192 57.395 39.256 ;
		RECT	56.144 39.193 56.176 39.257 ;
		RECT	55.035 39.399 55.067 39.431 ;
		RECT	52.968 39.672 53.032 39.736 ;
		RECT	55.528 39.672 55.592 39.736 ;
		RECT	56.664 39.672 56.696 39.736 ;
		RECT	57.509 39.672 57.573 39.736 ;
		RECT	54.137 39.853 54.169 39.885 ;
		RECT	57.51 39.853 57.542 39.885 ;
		RECT	52.15 40.363 52.182 40.395 ;
		RECT	50.33 40.458 50.362 40.49 ;
		RECT	52.221 40.538 52.253 40.57 ;
		RECT	55.876 40.618 55.908 40.65 ;
		RECT	52.15 40.903 52.182 40.935 ;
		RECT	54.065 41.53 54.097 41.562 ;
		RECT	55.81 41.53 55.842 41.562 ;
		RECT	52.078 41.87 52.11 41.902 ;
		RECT	54.065 41.87 54.097 41.902 ;
		RECT	53.104 41.97 53.136 42.002 ;
		RECT	50.662 42.425 50.694 42.457 ;
		RECT	52.291 42.425 52.323 42.457 ;
		RECT	52.454 42.425 52.486 42.457 ;
		RECT	54.359 42.425 54.391 42.457 ;
		RECT	55.81 42.425 55.842 42.457 ;
		RECT	52.221 42.52 52.253 42.552 ;
		RECT	57.253 42.52 57.285 42.552 ;
		RECT	50.658 42.659 50.69 42.723 ;
		RECT	52.968 42.675 53.032 42.707 ;
		RECT	54.251 42.675 54.283 42.707 ;
		RECT	55.562 42.675 55.626 42.707 ;
		RECT	50.658 42.864 50.69 42.928 ;
		RECT	52.968 42.864 53.032 42.928 ;
		RECT	54.251 42.864 54.283 42.928 ;
		RECT	55.562 42.864 55.626 42.928 ;
		RECT	50.658 43.069 50.69 43.133 ;
		RECT	54.251 43.069 54.283 43.133 ;
		RECT	52.968 43.085 53.032 43.117 ;
		RECT	55.562 43.085 55.626 43.117 ;
		RECT	52.454 43.467 52.486 43.499 ;
		RECT	52.026 44.026 52.058 44.09 ;
		RECT	54.251 44.026 54.283 44.09 ;
		RECT	55.842 44.026 55.874 44.09 ;
		RECT	52.968 44.042 53.032 44.074 ;
		RECT	55.562 44.042 55.626 44.074 ;
		RECT	52.13 44.199 52.162 44.231 ;
		RECT	53.104 44.469 53.136 44.501 ;
		RECT	53.104 44.759 53.136 44.791 ;
		RECT	50.658 45.197 50.69 45.229 ;
		RECT	53.245 45.197 53.277 45.229 ;
		RECT	53.094 46.057 53.126 46.089 ;
		RECT	53.095 46.632 53.127 46.664 ;
		RECT	50.557 47.367 50.589 47.399 ;
		RECT	52.277 47.467 52.309 47.499 ;
		RECT	54.359 47.467 54.391 47.499 ;
		RECT	52.454 48.217 52.486 48.249 ;
		RECT	50.332 48.317 50.364 48.349 ;
		RECT	52.047 49.263 52.079 49.327 ;
		RECT	54.735 50.027 54.767 50.059 ;
		RECT	53.997 34.896 54.029 34.928 ;
		RECT	58.031 45.197 58.063 45.229 ;
		RECT	52.15 37.474 52.182 37.506 ;
		RECT	55.462 47.367 55.494 47.399 ;
		RECT	53.104 41.004 53.136 41.036 ;
		RECT	55.528 35.741 55.56 35.773 ;
		RECT	52.15 39.192 52.182 39.256 ;
		RECT	52.454 39.192 52.486 39.256 ;
		RECT	52.968 39.192 53.032 39.256 ;
		RECT	56.664 39.192 56.696 39.256 ;
		RECT	50.417 39.672 50.481 39.736 ;
		RECT	51.274 39.672 51.306 39.736 ;
		RECT	51.92 39.672 51.952 39.736 ;
		RECT	53.894 39.672 53.926 39.736 ;
		RECT	54.363 39.672 54.427 39.736 ;
		RECT	54.804 39.672 54.836 39.736 ;
		RECT	55.969 39.672 56.033 39.736 ;
		RECT	56.144 39.672 56.176 39.736 ;
		RECT	57.363 39.672 57.395 39.736 ;
		RECT	51.92 42.659 51.952 42.723 ;
		RECT	53.91 42.659 53.942 42.723 ;
		RECT	54.812 42.659 54.844 42.723 ;
		RECT	55.969 42.675 56.033 42.707 ;
		RECT	51.92 42.864 51.952 42.928 ;
		RECT	53.91 42.864 53.942 42.928 ;
		RECT	54.812 42.864 54.844 42.928 ;
		RECT	55.969 42.864 56.033 42.928 ;
		RECT	51.92 43.069 51.952 43.133 ;
		RECT	53.91 43.069 53.942 43.133 ;
		RECT	54.812 43.069 54.844 43.133 ;
		RECT	55.969 43.085 56.033 43.117 ;
		RECT	54.657 44.026 54.689 44.09 ;
		RECT	54.809 44.026 54.841 44.09 ;
		RECT	55.208 44.042 55.272 44.074 ;
		RECT	51.967 2.939 51.999 2.971 ;
		RECT	53.91 3.044 53.942 3.076 ;
		RECT	50.379 3.374 50.443 3.406 ;
		RECT	51.274 3.374 51.306 3.406 ;
		RECT	51.794 3.374 51.826 3.406 ;
		RECT	53.707 3.374 53.739 3.406 ;
		RECT	55.216 3.374 55.28 3.406 ;
		RECT	56.144 3.374 56.176 3.406 ;
		RECT	56.664 3.374 56.696 3.406 ;
		RECT	57.531 3.374 57.595 3.406 ;
		RECT	52.036 3.479 52.068 3.511 ;
		RECT	55.57 3.613 55.602 3.677 ;
		RECT	52.124 3.629 52.156 3.661 ;
		RECT	52.577 3.629 52.609 3.661 ;
		RECT	53.148 3.629 53.18 3.661 ;
		RECT	54.246 3.629 54.278 3.661 ;
		RECT	55.807 3.629 55.839 3.661 ;
		RECT	51.967 20.219 51.999 20.251 ;
		RECT	53.91 20.324 53.942 20.356 ;
		RECT	50.379 20.654 50.443 20.686 ;
		RECT	51.274 20.654 51.306 20.686 ;
		RECT	51.794 20.654 51.826 20.686 ;
		RECT	53.707 20.654 53.739 20.686 ;
		RECT	55.216 20.654 55.28 20.686 ;
		RECT	56.144 20.654 56.176 20.686 ;
		RECT	56.664 20.654 56.696 20.686 ;
		RECT	57.531 20.654 57.595 20.686 ;
		RECT	52.036 20.759 52.068 20.791 ;
		RECT	55.57 20.893 55.602 20.957 ;
		RECT	52.124 20.909 52.156 20.941 ;
		RECT	52.577 20.909 52.609 20.941 ;
		RECT	53.148 20.909 53.18 20.941 ;
		RECT	54.246 20.909 54.278 20.941 ;
		RECT	55.807 20.909 55.839 20.941 ;
		RECT	51.967 22.139 51.999 22.171 ;
		RECT	53.91 22.244 53.942 22.276 ;
		RECT	50.379 22.574 50.443 22.606 ;
		RECT	51.274 22.574 51.306 22.606 ;
		RECT	51.794 22.574 51.826 22.606 ;
		RECT	53.707 22.574 53.739 22.606 ;
		RECT	55.216 22.574 55.28 22.606 ;
		RECT	56.144 22.574 56.176 22.606 ;
		RECT	56.664 22.574 56.696 22.606 ;
		RECT	57.531 22.574 57.595 22.606 ;
		RECT	52.036 22.679 52.068 22.711 ;
		RECT	55.57 22.813 55.602 22.877 ;
		RECT	52.124 22.829 52.156 22.861 ;
		RECT	52.577 22.829 52.609 22.861 ;
		RECT	53.148 22.829 53.18 22.861 ;
		RECT	54.246 22.829 54.278 22.861 ;
		RECT	55.807 22.829 55.839 22.861 ;
		RECT	51.967 24.059 51.999 24.091 ;
		RECT	53.91 24.164 53.942 24.196 ;
		RECT	50.379 24.494 50.443 24.526 ;
		RECT	51.274 24.494 51.306 24.526 ;
		RECT	51.794 24.494 51.826 24.526 ;
		RECT	53.707 24.494 53.739 24.526 ;
		RECT	55.216 24.494 55.28 24.526 ;
		RECT	56.144 24.494 56.176 24.526 ;
		RECT	56.664 24.494 56.696 24.526 ;
		RECT	57.531 24.494 57.595 24.526 ;
		RECT	52.036 24.599 52.068 24.631 ;
		RECT	55.57 24.733 55.602 24.797 ;
		RECT	52.124 24.749 52.156 24.781 ;
		RECT	52.577 24.749 52.609 24.781 ;
		RECT	53.148 24.749 53.18 24.781 ;
		RECT	54.246 24.749 54.278 24.781 ;
		RECT	55.807 24.749 55.839 24.781 ;
		RECT	51.967 25.979 51.999 26.011 ;
		RECT	53.91 26.084 53.942 26.116 ;
		RECT	50.379 26.414 50.443 26.446 ;
		RECT	51.274 26.414 51.306 26.446 ;
		RECT	51.794 26.414 51.826 26.446 ;
		RECT	53.707 26.414 53.739 26.446 ;
		RECT	55.216 26.414 55.28 26.446 ;
		RECT	56.144 26.414 56.176 26.446 ;
		RECT	56.664 26.414 56.696 26.446 ;
		RECT	57.531 26.414 57.595 26.446 ;
		RECT	52.036 26.519 52.068 26.551 ;
		RECT	55.57 26.653 55.602 26.717 ;
		RECT	52.124 26.669 52.156 26.701 ;
		RECT	52.577 26.669 52.609 26.701 ;
		RECT	53.148 26.669 53.18 26.701 ;
		RECT	54.246 26.669 54.278 26.701 ;
		RECT	55.807 26.669 55.839 26.701 ;
		RECT	51.967 27.899 51.999 27.931 ;
		RECT	53.91 28.004 53.942 28.036 ;
		RECT	50.379 28.334 50.443 28.366 ;
		RECT	51.274 28.334 51.306 28.366 ;
		RECT	51.794 28.334 51.826 28.366 ;
		RECT	53.707 28.334 53.739 28.366 ;
		RECT	55.216 28.334 55.28 28.366 ;
		RECT	56.144 28.334 56.176 28.366 ;
		RECT	56.664 28.334 56.696 28.366 ;
		RECT	57.531 28.334 57.595 28.366 ;
		RECT	52.036 28.439 52.068 28.471 ;
		RECT	55.57 28.573 55.602 28.637 ;
		RECT	52.124 28.589 52.156 28.621 ;
		RECT	52.577 28.589 52.609 28.621 ;
		RECT	53.148 28.589 53.18 28.621 ;
		RECT	54.246 28.589 54.278 28.621 ;
		RECT	55.807 28.589 55.839 28.621 ;
		RECT	51.967 4.859 51.999 4.891 ;
		RECT	53.91 4.964 53.942 4.996 ;
		RECT	50.379 5.294 50.443 5.326 ;
		RECT	51.274 5.294 51.306 5.326 ;
		RECT	51.794 5.294 51.826 5.326 ;
		RECT	53.707 5.294 53.739 5.326 ;
		RECT	55.216 5.294 55.28 5.326 ;
		RECT	56.144 5.294 56.176 5.326 ;
		RECT	56.664 5.294 56.696 5.326 ;
		RECT	57.531 5.294 57.595 5.326 ;
		RECT	52.036 5.399 52.068 5.431 ;
		RECT	55.57 5.533 55.602 5.597 ;
		RECT	52.124 5.549 52.156 5.581 ;
		RECT	52.577 5.549 52.609 5.581 ;
		RECT	53.148 5.549 53.18 5.581 ;
		RECT	54.246 5.549 54.278 5.581 ;
		RECT	55.807 5.549 55.839 5.581 ;
		RECT	51.967 6.779 51.999 6.811 ;
		RECT	53.91 6.884 53.942 6.916 ;
		RECT	50.379 7.214 50.443 7.246 ;
		RECT	51.274 7.214 51.306 7.246 ;
		RECT	51.794 7.214 51.826 7.246 ;
		RECT	53.707 7.214 53.739 7.246 ;
		RECT	55.216 7.214 55.28 7.246 ;
		RECT	56.144 7.214 56.176 7.246 ;
		RECT	56.664 7.214 56.696 7.246 ;
		RECT	57.531 7.214 57.595 7.246 ;
		RECT	52.036 7.319 52.068 7.351 ;
		RECT	55.57 7.453 55.602 7.517 ;
		RECT	52.124 7.469 52.156 7.501 ;
		RECT	52.577 7.469 52.609 7.501 ;
		RECT	53.148 7.469 53.18 7.501 ;
		RECT	54.246 7.469 54.278 7.501 ;
		RECT	55.807 7.469 55.839 7.501 ;
		RECT	51.967 8.699 51.999 8.731 ;
		RECT	53.91 8.804 53.942 8.836 ;
		RECT	50.379 9.134 50.443 9.166 ;
		RECT	51.274 9.134 51.306 9.166 ;
		RECT	51.794 9.134 51.826 9.166 ;
		RECT	53.707 9.134 53.739 9.166 ;
		RECT	55.216 9.134 55.28 9.166 ;
		RECT	56.144 9.134 56.176 9.166 ;
		RECT	56.664 9.134 56.696 9.166 ;
		RECT	57.531 9.134 57.595 9.166 ;
		RECT	52.036 9.239 52.068 9.271 ;
		RECT	55.57 9.373 55.602 9.437 ;
		RECT	52.124 9.389 52.156 9.421 ;
		RECT	52.577 9.389 52.609 9.421 ;
		RECT	53.148 9.389 53.18 9.421 ;
		RECT	54.246 9.389 54.278 9.421 ;
		RECT	55.807 9.389 55.839 9.421 ;
		RECT	51.967 10.619 51.999 10.651 ;
		RECT	53.91 10.724 53.942 10.756 ;
		RECT	50.379 11.054 50.443 11.086 ;
		RECT	51.274 11.054 51.306 11.086 ;
		RECT	51.794 11.054 51.826 11.086 ;
		RECT	53.707 11.054 53.739 11.086 ;
		RECT	55.216 11.054 55.28 11.086 ;
		RECT	56.144 11.054 56.176 11.086 ;
		RECT	56.664 11.054 56.696 11.086 ;
		RECT	57.531 11.054 57.595 11.086 ;
		RECT	52.036 11.159 52.068 11.191 ;
		RECT	55.57 11.293 55.602 11.357 ;
		RECT	52.124 11.309 52.156 11.341 ;
		RECT	52.577 11.309 52.609 11.341 ;
		RECT	53.148 11.309 53.18 11.341 ;
		RECT	54.246 11.309 54.278 11.341 ;
		RECT	55.807 11.309 55.839 11.341 ;
		RECT	51.967 12.539 51.999 12.571 ;
		RECT	53.91 12.644 53.942 12.676 ;
		RECT	50.379 12.974 50.443 13.006 ;
		RECT	51.274 12.974 51.306 13.006 ;
		RECT	51.794 12.974 51.826 13.006 ;
		RECT	53.707 12.974 53.739 13.006 ;
		RECT	55.216 12.974 55.28 13.006 ;
		RECT	56.144 12.974 56.176 13.006 ;
		RECT	56.664 12.974 56.696 13.006 ;
		RECT	57.531 12.974 57.595 13.006 ;
		RECT	52.036 13.079 52.068 13.111 ;
		RECT	55.57 13.213 55.602 13.277 ;
		RECT	52.124 13.229 52.156 13.261 ;
		RECT	52.577 13.229 52.609 13.261 ;
		RECT	53.148 13.229 53.18 13.261 ;
		RECT	54.246 13.229 54.278 13.261 ;
		RECT	55.807 13.229 55.839 13.261 ;
		RECT	51.967 14.459 51.999 14.491 ;
		RECT	53.91 14.564 53.942 14.596 ;
		RECT	50.379 14.894 50.443 14.926 ;
		RECT	51.274 14.894 51.306 14.926 ;
		RECT	51.794 14.894 51.826 14.926 ;
		RECT	53.707 14.894 53.739 14.926 ;
		RECT	55.216 14.894 55.28 14.926 ;
		RECT	56.144 14.894 56.176 14.926 ;
		RECT	56.664 14.894 56.696 14.926 ;
		RECT	57.531 14.894 57.595 14.926 ;
		RECT	52.036 14.999 52.068 15.031 ;
		RECT	55.57 15.133 55.602 15.197 ;
		RECT	52.124 15.149 52.156 15.181 ;
		RECT	52.577 15.149 52.609 15.181 ;
		RECT	53.148 15.149 53.18 15.181 ;
		RECT	54.246 15.149 54.278 15.181 ;
		RECT	55.807 15.149 55.839 15.181 ;
		RECT	51.967 16.379 51.999 16.411 ;
		RECT	53.91 16.484 53.942 16.516 ;
		RECT	50.379 16.814 50.443 16.846 ;
		RECT	51.274 16.814 51.306 16.846 ;
		RECT	51.794 16.814 51.826 16.846 ;
		RECT	53.707 16.814 53.739 16.846 ;
		RECT	55.216 16.814 55.28 16.846 ;
		RECT	56.144 16.814 56.176 16.846 ;
		RECT	56.664 16.814 56.696 16.846 ;
		RECT	57.531 16.814 57.595 16.846 ;
		RECT	52.036 16.919 52.068 16.951 ;
		RECT	55.57 17.053 55.602 17.117 ;
		RECT	52.124 17.069 52.156 17.101 ;
		RECT	52.577 17.069 52.609 17.101 ;
		RECT	53.148 17.069 53.18 17.101 ;
		RECT	54.246 17.069 54.278 17.101 ;
		RECT	55.807 17.069 55.839 17.101 ;
		RECT	51.967 18.299 51.999 18.331 ;
		RECT	53.91 18.404 53.942 18.436 ;
		RECT	50.379 18.734 50.443 18.766 ;
		RECT	51.274 18.734 51.306 18.766 ;
		RECT	51.794 18.734 51.826 18.766 ;
		RECT	53.707 18.734 53.739 18.766 ;
		RECT	55.216 18.734 55.28 18.766 ;
		RECT	56.144 18.734 56.176 18.766 ;
		RECT	56.664 18.734 56.696 18.766 ;
		RECT	57.531 18.734 57.595 18.766 ;
		RECT	52.036 18.839 52.068 18.871 ;
		RECT	55.57 18.973 55.602 19.037 ;
		RECT	52.124 18.989 52.156 19.021 ;
		RECT	52.577 18.989 52.609 19.021 ;
		RECT	53.148 18.989 53.18 19.021 ;
		RECT	54.246 18.989 54.278 19.021 ;
		RECT	55.807 18.989 55.839 19.021 ;
		RECT	51.967 1.019 51.999 1.051 ;
		RECT	53.91 1.124 53.942 1.156 ;
		RECT	50.379 1.454 50.443 1.486 ;
		RECT	51.274 1.454 51.306 1.486 ;
		RECT	51.794 1.454 51.826 1.486 ;
		RECT	53.707 1.454 53.739 1.486 ;
		RECT	55.216 1.454 55.28 1.486 ;
		RECT	56.144 1.454 56.176 1.486 ;
		RECT	56.664 1.454 56.696 1.486 ;
		RECT	57.531 1.454 57.595 1.486 ;
		RECT	52.036 1.559 52.068 1.591 ;
		RECT	55.57 1.693 55.602 1.757 ;
		RECT	52.124 1.709 52.156 1.741 ;
		RECT	52.577 1.709 52.609 1.741 ;
		RECT	53.148 1.709 53.18 1.741 ;
		RECT	54.246 1.709 54.278 1.741 ;
		RECT	55.807 1.709 55.839 1.741 ;
		RECT	51.967 29.819 51.999 29.851 ;
		RECT	53.91 29.924 53.942 29.956 ;
		RECT	50.379 30.254 50.443 30.286 ;
		RECT	51.274 30.254 51.306 30.286 ;
		RECT	51.794 30.254 51.826 30.286 ;
		RECT	53.707 30.254 53.739 30.286 ;
		RECT	55.216 30.254 55.28 30.286 ;
		RECT	56.144 30.254 56.176 30.286 ;
		RECT	56.664 30.254 56.696 30.286 ;
		RECT	57.531 30.254 57.595 30.286 ;
		RECT	52.036 30.359 52.068 30.391 ;
		RECT	55.57 30.493 55.602 30.557 ;
		RECT	52.124 30.509 52.156 30.541 ;
		RECT	52.577 30.509 52.609 30.541 ;
		RECT	53.148 30.509 53.18 30.541 ;
		RECT	54.246 30.509 54.278 30.541 ;
		RECT	55.807 30.509 55.839 30.541 ;
		RECT	52.459 2.074 52.491 2.106 ;
		RECT	52.459 3.994 52.491 4.026 ;
		RECT	52.459 5.914 52.491 5.946 ;
		RECT	52.459 7.834 52.491 7.866 ;
		RECT	52.459 9.754 52.491 9.786 ;
		RECT	52.459 11.674 52.491 11.706 ;
		RECT	52.459 13.594 52.491 13.626 ;
		RECT	52.459 15.514 52.491 15.546 ;
		RECT	52.459 17.434 52.491 17.466 ;
		RECT	52.459 19.354 52.491 19.386 ;
		RECT	52.459 21.274 52.491 21.306 ;
		RECT	52.459 23.194 52.491 23.226 ;
		RECT	52.459 25.114 52.491 25.146 ;
		RECT	52.459 27.034 52.491 27.066 ;
		RECT	52.459 28.954 52.491 28.986 ;
		RECT	52.459 30.874 52.491 30.906 ;
		RECT	53.91 1.693 53.942 1.757 ;
		RECT	53.91 20.893 53.942 20.957 ;
		RECT	53.91 22.813 53.942 22.877 ;
		RECT	53.91 24.733 53.942 24.797 ;
		RECT	53.91 26.653 53.942 26.717 ;
		RECT	53.91 28.573 53.942 28.637 ;
		RECT	53.91 30.493 53.942 30.557 ;
		RECT	53.91 3.613 53.942 3.677 ;
		RECT	53.91 5.533 53.942 5.597 ;
		RECT	53.91 7.453 53.942 7.517 ;
		RECT	53.91 9.373 53.942 9.437 ;
		RECT	53.91 11.293 53.942 11.357 ;
		RECT	53.91 13.213 53.942 13.277 ;
		RECT	53.91 15.133 53.942 15.197 ;
		RECT	53.91 17.053 53.942 17.117 ;
		RECT	53.91 18.973 53.942 19.037 ;
		RECT	51.967 54.245 51.999 54.277 ;
		RECT	53.91 54.14 53.942 54.172 ;
		RECT	50.379 53.81 50.443 53.842 ;
		RECT	51.274 53.81 51.306 53.842 ;
		RECT	51.794 53.81 51.826 53.842 ;
		RECT	53.707 53.81 53.739 53.842 ;
		RECT	55.216 53.81 55.28 53.842 ;
		RECT	56.144 53.81 56.176 53.842 ;
		RECT	56.664 53.81 56.696 53.842 ;
		RECT	57.531 53.81 57.595 53.842 ;
		RECT	52.036 53.705 52.068 53.737 ;
		RECT	55.57 53.539 55.602 53.603 ;
		RECT	52.124 53.555 52.156 53.587 ;
		RECT	52.577 53.555 52.609 53.587 ;
		RECT	53.148 53.555 53.18 53.587 ;
		RECT	54.246 53.555 54.278 53.587 ;
		RECT	55.807 53.555 55.839 53.587 ;
		RECT	51.967 71.525 51.999 71.557 ;
		RECT	53.91 71.42 53.942 71.452 ;
		RECT	50.379 71.09 50.443 71.122 ;
		RECT	51.274 71.09 51.306 71.122 ;
		RECT	51.794 71.09 51.826 71.122 ;
		RECT	53.707 71.09 53.739 71.122 ;
		RECT	55.216 71.09 55.28 71.122 ;
		RECT	56.144 71.09 56.176 71.122 ;
		RECT	56.664 71.09 56.696 71.122 ;
		RECT	57.531 71.09 57.595 71.122 ;
		RECT	52.036 70.985 52.068 71.017 ;
		RECT	55.57 70.819 55.602 70.883 ;
		RECT	52.124 70.835 52.156 70.867 ;
		RECT	52.577 70.835 52.609 70.867 ;
		RECT	53.148 70.835 53.18 70.867 ;
		RECT	54.246 70.835 54.278 70.867 ;
		RECT	55.807 70.835 55.839 70.867 ;
		RECT	51.967 73.445 51.999 73.477 ;
		RECT	53.91 73.34 53.942 73.372 ;
		RECT	50.379 73.01 50.443 73.042 ;
		RECT	51.274 73.01 51.306 73.042 ;
		RECT	51.794 73.01 51.826 73.042 ;
		RECT	53.707 73.01 53.739 73.042 ;
		RECT	55.216 73.01 55.28 73.042 ;
		RECT	56.144 73.01 56.176 73.042 ;
		RECT	56.664 73.01 56.696 73.042 ;
		RECT	57.531 73.01 57.595 73.042 ;
		RECT	52.036 72.905 52.068 72.937 ;
		RECT	55.57 72.739 55.602 72.803 ;
		RECT	52.124 72.755 52.156 72.787 ;
		RECT	52.577 72.755 52.609 72.787 ;
		RECT	53.148 72.755 53.18 72.787 ;
		RECT	54.246 72.755 54.278 72.787 ;
		RECT	55.807 72.755 55.839 72.787 ;
		RECT	51.967 75.365 51.999 75.397 ;
		RECT	53.91 75.26 53.942 75.292 ;
		RECT	50.379 74.93 50.443 74.962 ;
		RECT	51.274 74.93 51.306 74.962 ;
		RECT	51.794 74.93 51.826 74.962 ;
		RECT	53.707 74.93 53.739 74.962 ;
		RECT	55.216 74.93 55.28 74.962 ;
		RECT	56.144 74.93 56.176 74.962 ;
		RECT	56.664 74.93 56.696 74.962 ;
		RECT	57.531 74.93 57.595 74.962 ;
		RECT	52.036 74.825 52.068 74.857 ;
		RECT	55.57 74.659 55.602 74.723 ;
		RECT	52.124 74.675 52.156 74.707 ;
		RECT	52.577 74.675 52.609 74.707 ;
		RECT	53.148 74.675 53.18 74.707 ;
		RECT	54.246 74.675 54.278 74.707 ;
		RECT	55.807 74.675 55.839 74.707 ;
		RECT	51.967 77.285 51.999 77.317 ;
		RECT	53.91 77.18 53.942 77.212 ;
		RECT	50.379 76.85 50.443 76.882 ;
		RECT	51.274 76.85 51.306 76.882 ;
		RECT	51.794 76.85 51.826 76.882 ;
		RECT	53.707 76.85 53.739 76.882 ;
		RECT	55.216 76.85 55.28 76.882 ;
		RECT	56.144 76.85 56.176 76.882 ;
		RECT	56.664 76.85 56.696 76.882 ;
		RECT	57.531 76.85 57.595 76.882 ;
		RECT	52.036 76.745 52.068 76.777 ;
		RECT	55.57 76.579 55.602 76.643 ;
		RECT	52.124 76.595 52.156 76.627 ;
		RECT	52.577 76.595 52.609 76.627 ;
		RECT	53.148 76.595 53.18 76.627 ;
		RECT	54.246 76.595 54.278 76.627 ;
		RECT	55.807 76.595 55.839 76.627 ;
		RECT	51.967 79.205 51.999 79.237 ;
		RECT	53.91 79.1 53.942 79.132 ;
		RECT	50.379 78.77 50.443 78.802 ;
		RECT	51.274 78.77 51.306 78.802 ;
		RECT	51.794 78.77 51.826 78.802 ;
		RECT	53.707 78.77 53.739 78.802 ;
		RECT	55.216 78.77 55.28 78.802 ;
		RECT	56.144 78.77 56.176 78.802 ;
		RECT	56.664 78.77 56.696 78.802 ;
		RECT	57.531 78.77 57.595 78.802 ;
		RECT	52.036 78.665 52.068 78.697 ;
		RECT	55.57 78.499 55.602 78.563 ;
		RECT	52.124 78.515 52.156 78.547 ;
		RECT	52.577 78.515 52.609 78.547 ;
		RECT	53.148 78.515 53.18 78.547 ;
		RECT	54.246 78.515 54.278 78.547 ;
		RECT	55.807 78.515 55.839 78.547 ;
		RECT	51.967 56.165 51.999 56.197 ;
		RECT	53.91 56.06 53.942 56.092 ;
		RECT	50.379 55.73 50.443 55.762 ;
		RECT	51.274 55.73 51.306 55.762 ;
		RECT	51.794 55.73 51.826 55.762 ;
		RECT	53.707 55.73 53.739 55.762 ;
		RECT	55.216 55.73 55.28 55.762 ;
		RECT	56.144 55.73 56.176 55.762 ;
		RECT	56.664 55.73 56.696 55.762 ;
		RECT	57.531 55.73 57.595 55.762 ;
		RECT	52.036 55.625 52.068 55.657 ;
		RECT	55.57 55.459 55.602 55.523 ;
		RECT	52.124 55.475 52.156 55.507 ;
		RECT	52.577 55.475 52.609 55.507 ;
		RECT	53.148 55.475 53.18 55.507 ;
		RECT	54.246 55.475 54.278 55.507 ;
		RECT	55.807 55.475 55.839 55.507 ;
		RECT	51.967 58.085 51.999 58.117 ;
		RECT	53.91 57.98 53.942 58.012 ;
		RECT	50.379 57.65 50.443 57.682 ;
		RECT	51.274 57.65 51.306 57.682 ;
		RECT	51.794 57.65 51.826 57.682 ;
		RECT	53.707 57.65 53.739 57.682 ;
		RECT	55.216 57.65 55.28 57.682 ;
		RECT	56.144 57.65 56.176 57.682 ;
		RECT	56.664 57.65 56.696 57.682 ;
		RECT	57.531 57.65 57.595 57.682 ;
		RECT	52.036 57.545 52.068 57.577 ;
		RECT	55.57 57.379 55.602 57.443 ;
		RECT	52.124 57.395 52.156 57.427 ;
		RECT	52.577 57.395 52.609 57.427 ;
		RECT	53.148 57.395 53.18 57.427 ;
		RECT	54.246 57.395 54.278 57.427 ;
		RECT	55.807 57.395 55.839 57.427 ;
		RECT	51.967 60.005 51.999 60.037 ;
		RECT	53.91 59.9 53.942 59.932 ;
		RECT	50.379 59.57 50.443 59.602 ;
		RECT	51.274 59.57 51.306 59.602 ;
		RECT	51.794 59.57 51.826 59.602 ;
		RECT	53.707 59.57 53.739 59.602 ;
		RECT	55.216 59.57 55.28 59.602 ;
		RECT	56.144 59.57 56.176 59.602 ;
		RECT	56.664 59.57 56.696 59.602 ;
		RECT	57.531 59.57 57.595 59.602 ;
		RECT	52.036 59.465 52.068 59.497 ;
		RECT	55.57 59.299 55.602 59.363 ;
		RECT	52.124 59.315 52.156 59.347 ;
		RECT	52.577 59.315 52.609 59.347 ;
		RECT	53.148 59.315 53.18 59.347 ;
		RECT	54.246 59.315 54.278 59.347 ;
		RECT	55.807 59.315 55.839 59.347 ;
		RECT	51.967 61.925 51.999 61.957 ;
		RECT	53.91 61.82 53.942 61.852 ;
		RECT	50.379 61.49 50.443 61.522 ;
		RECT	51.274 61.49 51.306 61.522 ;
		RECT	51.794 61.49 51.826 61.522 ;
		RECT	53.707 61.49 53.739 61.522 ;
		RECT	55.216 61.49 55.28 61.522 ;
		RECT	56.144 61.49 56.176 61.522 ;
		RECT	56.664 61.49 56.696 61.522 ;
		RECT	57.531 61.49 57.595 61.522 ;
		RECT	52.036 61.385 52.068 61.417 ;
		RECT	55.57 61.219 55.602 61.283 ;
		RECT	52.124 61.235 52.156 61.267 ;
		RECT	52.577 61.235 52.609 61.267 ;
		RECT	53.148 61.235 53.18 61.267 ;
		RECT	54.246 61.235 54.278 61.267 ;
		RECT	55.807 61.235 55.839 61.267 ;
		RECT	51.967 63.845 51.999 63.877 ;
		RECT	53.91 63.74 53.942 63.772 ;
		RECT	50.379 63.41 50.443 63.442 ;
		RECT	51.274 63.41 51.306 63.442 ;
		RECT	51.794 63.41 51.826 63.442 ;
		RECT	53.707 63.41 53.739 63.442 ;
		RECT	55.216 63.41 55.28 63.442 ;
		RECT	56.144 63.41 56.176 63.442 ;
		RECT	56.664 63.41 56.696 63.442 ;
		RECT	57.531 63.41 57.595 63.442 ;
		RECT	52.036 63.305 52.068 63.337 ;
		RECT	55.57 63.139 55.602 63.203 ;
		RECT	52.124 63.155 52.156 63.187 ;
		RECT	52.577 63.155 52.609 63.187 ;
		RECT	53.148 63.155 53.18 63.187 ;
		RECT	54.246 63.155 54.278 63.187 ;
		RECT	55.807 63.155 55.839 63.187 ;
		RECT	51.967 65.765 51.999 65.797 ;
		RECT	53.91 65.66 53.942 65.692 ;
		RECT	50.379 65.33 50.443 65.362 ;
		RECT	51.274 65.33 51.306 65.362 ;
		RECT	51.794 65.33 51.826 65.362 ;
		RECT	53.707 65.33 53.739 65.362 ;
		RECT	55.216 65.33 55.28 65.362 ;
		RECT	56.144 65.33 56.176 65.362 ;
		RECT	56.664 65.33 56.696 65.362 ;
		RECT	57.531 65.33 57.595 65.362 ;
		RECT	52.036 65.225 52.068 65.257 ;
		RECT	55.57 65.059 55.602 65.123 ;
		RECT	52.124 65.075 52.156 65.107 ;
		RECT	52.577 65.075 52.609 65.107 ;
		RECT	53.148 65.075 53.18 65.107 ;
		RECT	54.246 65.075 54.278 65.107 ;
		RECT	55.807 65.075 55.839 65.107 ;
		RECT	51.967 67.685 51.999 67.717 ;
		RECT	53.91 67.58 53.942 67.612 ;
		RECT	50.379 67.25 50.443 67.282 ;
		RECT	51.274 67.25 51.306 67.282 ;
		RECT	51.794 67.25 51.826 67.282 ;
		RECT	53.707 67.25 53.739 67.282 ;
		RECT	55.216 67.25 55.28 67.282 ;
		RECT	56.144 67.25 56.176 67.282 ;
		RECT	56.664 67.25 56.696 67.282 ;
		RECT	57.531 67.25 57.595 67.282 ;
		RECT	52.036 67.145 52.068 67.177 ;
		RECT	55.57 66.979 55.602 67.043 ;
		RECT	52.124 66.995 52.156 67.027 ;
		RECT	52.577 66.995 52.609 67.027 ;
		RECT	53.148 66.995 53.18 67.027 ;
		RECT	54.246 66.995 54.278 67.027 ;
		RECT	55.807 66.995 55.839 67.027 ;
		RECT	51.967 69.605 51.999 69.637 ;
		RECT	53.91 69.5 53.942 69.532 ;
		RECT	50.379 69.17 50.443 69.202 ;
		RECT	51.274 69.17 51.306 69.202 ;
		RECT	51.794 69.17 51.826 69.202 ;
		RECT	53.707 69.17 53.739 69.202 ;
		RECT	55.216 69.17 55.28 69.202 ;
		RECT	56.144 69.17 56.176 69.202 ;
		RECT	56.664 69.17 56.696 69.202 ;
		RECT	57.531 69.17 57.595 69.202 ;
		RECT	52.036 69.065 52.068 69.097 ;
		RECT	55.57 68.899 55.602 68.963 ;
		RECT	52.124 68.915 52.156 68.947 ;
		RECT	52.577 68.915 52.609 68.947 ;
		RECT	53.148 68.915 53.18 68.947 ;
		RECT	54.246 68.915 54.278 68.947 ;
		RECT	55.807 68.915 55.839 68.947 ;
		RECT	51.967 52.325 51.999 52.357 ;
		RECT	53.91 52.22 53.942 52.252 ;
		RECT	50.379 51.89 50.443 51.922 ;
		RECT	51.274 51.89 51.306 51.922 ;
		RECT	51.794 51.89 51.826 51.922 ;
		RECT	53.707 51.89 53.739 51.922 ;
		RECT	55.216 51.89 55.28 51.922 ;
		RECT	56.144 51.89 56.176 51.922 ;
		RECT	56.664 51.89 56.696 51.922 ;
		RECT	57.531 51.89 57.595 51.922 ;
		RECT	52.036 51.785 52.068 51.817 ;
		RECT	55.57 51.619 55.602 51.683 ;
		RECT	52.124 51.635 52.156 51.667 ;
		RECT	52.577 51.635 52.609 51.667 ;
		RECT	53.148 51.635 53.18 51.667 ;
		RECT	54.246 51.635 54.278 51.667 ;
		RECT	55.807 51.635 55.839 51.667 ;
		RECT	51.967 81.125 51.999 81.157 ;
		RECT	53.91 81.02 53.942 81.052 ;
		RECT	50.379 80.69 50.443 80.722 ;
		RECT	51.274 80.69 51.306 80.722 ;
		RECT	51.794 80.69 51.826 80.722 ;
		RECT	53.707 80.69 53.739 80.722 ;
		RECT	55.216 80.69 55.28 80.722 ;
		RECT	56.144 80.69 56.176 80.722 ;
		RECT	56.664 80.69 56.696 80.722 ;
		RECT	57.531 80.69 57.595 80.722 ;
		RECT	52.036 80.585 52.068 80.617 ;
		RECT	55.57 80.419 55.602 80.483 ;
		RECT	52.124 80.435 52.156 80.467 ;
		RECT	52.577 80.435 52.609 80.467 ;
		RECT	53.148 80.435 53.18 80.467 ;
		RECT	54.246 80.435 54.278 80.467 ;
		RECT	55.807 80.435 55.839 80.467 ;
		RECT	52.459 51.27 52.491 51.302 ;
		RECT	52.459 53.19 52.491 53.222 ;
		RECT	52.459 55.11 52.491 55.142 ;
		RECT	52.459 57.03 52.491 57.062 ;
		RECT	52.459 58.95 52.491 58.982 ;
		RECT	52.459 60.87 52.491 60.902 ;
		RECT	52.459 62.79 52.491 62.822 ;
		RECT	52.459 64.71 52.491 64.742 ;
		RECT	52.459 66.63 52.491 66.662 ;
		RECT	52.459 68.55 52.491 68.582 ;
		RECT	52.459 70.47 52.491 70.502 ;
		RECT	52.459 72.39 52.491 72.422 ;
		RECT	52.459 74.31 52.491 74.342 ;
		RECT	52.459 76.23 52.491 76.262 ;
		RECT	52.459 78.15 52.491 78.182 ;
		RECT	52.459 80.07 52.491 80.102 ;
		RECT	53.91 51.619 53.942 51.683 ;
		RECT	53.91 70.819 53.942 70.883 ;
		RECT	53.91 72.739 53.942 72.803 ;
		RECT	53.91 74.659 53.942 74.723 ;
		RECT	53.91 76.579 53.942 76.643 ;
		RECT	53.91 78.499 53.942 78.563 ;
		RECT	53.91 80.419 53.942 80.483 ;
		RECT	53.91 53.539 53.942 53.603 ;
		RECT	53.91 55.459 53.942 55.523 ;
		RECT	53.91 57.379 53.942 57.443 ;
		RECT	53.91 59.299 53.942 59.363 ;
		RECT	53.91 61.219 53.942 61.283 ;
		RECT	53.91 63.139 53.942 63.203 ;
		RECT	53.91 65.059 53.942 65.123 ;
		RECT	53.91 66.979 53.942 67.043 ;
		RECT	53.91 68.899 53.942 68.963 ;
		RECT	5.514 31.762 5.578 31.794 ;
		RECT	5.514 50.382 5.578 50.414 ;
		RECT	27.557 39.858 27.589 39.89 ;
		RECT	24.197 39.358 24.229 39.39 ;
		RECT	23.861 39.358 23.893 39.39 ;
		RECT	23.525 39.258 23.557 39.29 ;
		RECT	23.189 39.258 23.221 39.29 ;
		RECT	22.853 39.158 22.885 39.19 ;
		RECT	22.517 39.158 22.549 39.19 ;
		RECT	22.181 39.858 22.213 39.89 ;
		RECT	21.845 39.858 21.877 39.89 ;
		RECT	21.509 39.758 21.541 39.79 ;
		RECT	21.173 39.758 21.205 39.79 ;
		RECT	27.221 39.858 27.253 39.89 ;
		RECT	20.837 39.658 20.869 39.69 ;
		RECT	20.501 39.658 20.533 39.69 ;
		RECT	20.165 39.558 20.197 39.59 ;
		RECT	19.829 39.558 19.861 39.59 ;
		RECT	19.493 39.458 19.525 39.49 ;
		RECT	19.157 39.458 19.189 39.49 ;
		RECT	18.821 39.358 18.853 39.39 ;
		RECT	18.485 39.358 18.517 39.39 ;
		RECT	18.149 39.258 18.181 39.29 ;
		RECT	17.813 39.258 17.845 39.29 ;
		RECT	26.885 39.758 26.917 39.79 ;
		RECT	17.477 39.158 17.509 39.19 ;
		RECT	17.141 39.158 17.173 39.19 ;
		RECT	16.805 39.858 16.837 39.89 ;
		RECT	16.469 39.858 16.501 39.89 ;
		RECT	16.133 39.758 16.165 39.79 ;
		RECT	15.797 39.758 15.829 39.79 ;
		RECT	15.461 39.658 15.493 39.69 ;
		RECT	15.125 39.658 15.157 39.69 ;
		RECT	14.789 39.558 14.821 39.59 ;
		RECT	14.453 39.558 14.485 39.59 ;
		RECT	26.549 39.758 26.581 39.79 ;
		RECT	14.117 39.458 14.149 39.49 ;
		RECT	13.781 39.458 13.813 39.49 ;
		RECT	13.445 39.358 13.477 39.39 ;
		RECT	13.109 39.358 13.141 39.39 ;
		RECT	12.773 39.258 12.805 39.29 ;
		RECT	12.437 39.258 12.469 39.29 ;
		RECT	12.101 39.158 12.133 39.19 ;
		RECT	11.765 39.158 11.797 39.19 ;
		RECT	11.429 39.858 11.461 39.89 ;
		RECT	11.093 39.858 11.125 39.89 ;
		RECT	26.213 39.658 26.245 39.69 ;
		RECT	10.757 39.758 10.789 39.79 ;
		RECT	10.421 39.758 10.453 39.79 ;
		RECT	10.085 39.658 10.117 39.69 ;
		RECT	9.749 39.658 9.781 39.69 ;
		RECT	9.413 39.558 9.445 39.59 ;
		RECT	9.077 39.558 9.109 39.59 ;
		RECT	8.741 39.458 8.773 39.49 ;
		RECT	8.405 39.458 8.437 39.49 ;
		RECT	8.069 39.358 8.101 39.39 ;
		RECT	7.733 39.358 7.765 39.39 ;
		RECT	25.877 39.658 25.909 39.69 ;
		RECT	7.397 39.258 7.429 39.29 ;
		RECT	7.061 39.258 7.093 39.29 ;
		RECT	6.725 39.158 6.757 39.19 ;
		RECT	6.389 39.158 6.421 39.19 ;
		RECT	25.541 39.558 25.573 39.59 ;
		RECT	25.205 39.558 25.237 39.59 ;
		RECT	24.869 39.458 24.901 39.49 ;
		RECT	24.533 39.458 24.565 39.49 ;
		RECT	27.557 42.825 27.589 42.857 ;
		RECT	24.197 42.825 24.229 42.857 ;
		RECT	23.861 42.825 23.893 42.857 ;
		RECT	23.525 42.825 23.557 42.857 ;
		RECT	23.189 42.825 23.221 42.857 ;
		RECT	22.853 42.825 22.885 42.857 ;
		RECT	22.517 42.825 22.549 42.857 ;
		RECT	22.181 42.925 22.213 42.957 ;
		RECT	21.845 42.925 21.877 42.957 ;
		RECT	21.509 42.925 21.541 42.957 ;
		RECT	21.173 42.925 21.205 42.957 ;
		RECT	27.221 42.825 27.253 42.857 ;
		RECT	20.837 42.925 20.869 42.957 ;
		RECT	20.501 42.925 20.533 42.957 ;
		RECT	20.165 42.925 20.197 42.957 ;
		RECT	19.829 42.925 19.861 42.957 ;
		RECT	19.493 42.925 19.525 42.957 ;
		RECT	19.157 42.925 19.189 42.957 ;
		RECT	18.821 42.925 18.853 42.957 ;
		RECT	18.485 42.925 18.517 42.957 ;
		RECT	18.149 42.925 18.181 42.957 ;
		RECT	17.813 42.925 17.845 42.957 ;
		RECT	26.885 42.825 26.917 42.857 ;
		RECT	17.477 42.925 17.509 42.957 ;
		RECT	17.141 42.925 17.173 42.957 ;
		RECT	16.805 43.025 16.837 43.057 ;
		RECT	16.469 43.025 16.501 43.057 ;
		RECT	16.133 43.025 16.165 43.057 ;
		RECT	15.797 43.025 15.829 43.057 ;
		RECT	15.461 43.025 15.493 43.057 ;
		RECT	15.125 43.025 15.157 43.057 ;
		RECT	14.789 43.025 14.821 43.057 ;
		RECT	14.453 43.025 14.485 43.057 ;
		RECT	26.549 42.825 26.581 42.857 ;
		RECT	14.117 43.025 14.149 43.057 ;
		RECT	13.781 43.025 13.813 43.057 ;
		RECT	13.445 43.025 13.477 43.057 ;
		RECT	13.109 43.025 13.141 43.057 ;
		RECT	12.773 43.025 12.805 43.057 ;
		RECT	12.437 43.025 12.469 43.057 ;
		RECT	12.101 43.025 12.133 43.057 ;
		RECT	11.765 43.025 11.797 43.057 ;
		RECT	11.429 43.125 11.461 43.157 ;
		RECT	11.093 43.125 11.125 43.157 ;
		RECT	26.213 42.825 26.245 42.857 ;
		RECT	10.757 43.125 10.789 43.157 ;
		RECT	10.421 43.125 10.453 43.157 ;
		RECT	10.085 43.125 10.117 43.157 ;
		RECT	9.749 43.125 9.781 43.157 ;
		RECT	9.413 43.125 9.445 43.157 ;
		RECT	9.077 43.125 9.109 43.157 ;
		RECT	8.741 43.125 8.773 43.157 ;
		RECT	8.405 43.125 8.437 43.157 ;
		RECT	8.069 43.125 8.101 43.157 ;
		RECT	7.733 43.125 7.765 43.157 ;
		RECT	25.877 42.825 25.909 42.857 ;
		RECT	7.397 43.125 7.429 43.157 ;
		RECT	7.061 43.125 7.093 43.157 ;
		RECT	6.725 43.125 6.757 43.157 ;
		RECT	6.389 43.125 6.421 43.157 ;
		RECT	25.541 42.825 25.573 42.857 ;
		RECT	25.205 42.825 25.237 42.857 ;
		RECT	24.869 42.825 24.901 42.857 ;
		RECT	24.533 42.825 24.565 42.857 ;
		RECT	27.515 32.691 27.547 32.755 ;
		RECT	49.711 39.672 49.743 39.736 ;
		RECT	49.675 44.026 49.707 44.09 ;
		RECT	24.155 32.691 24.187 32.755 ;
		RECT	23.819 32.691 23.851 32.755 ;
		RECT	23.483 32.691 23.515 32.755 ;
		RECT	23.147 32.691 23.179 32.755 ;
		RECT	22.811 32.691 22.843 32.755 ;
		RECT	22.475 32.691 22.507 32.755 ;
		RECT	22.139 32.691 22.171 32.755 ;
		RECT	21.803 32.691 21.835 32.755 ;
		RECT	21.467 32.691 21.499 32.755 ;
		RECT	21.131 32.691 21.163 32.755 ;
		RECT	27.179 32.691 27.211 32.755 ;
		RECT	20.795 32.691 20.827 32.755 ;
		RECT	20.459 32.691 20.491 32.755 ;
		RECT	20.123 32.691 20.155 32.755 ;
		RECT	19.787 32.691 19.819 32.755 ;
		RECT	19.451 32.691 19.483 32.755 ;
		RECT	19.115 32.691 19.147 32.755 ;
		RECT	18.779 32.691 18.811 32.755 ;
		RECT	18.443 32.691 18.475 32.755 ;
		RECT	18.107 32.691 18.139 32.755 ;
		RECT	17.771 32.691 17.803 32.755 ;
		RECT	26.843 32.691 26.875 32.755 ;
		RECT	17.435 32.691 17.467 32.755 ;
		RECT	17.099 32.691 17.131 32.755 ;
		RECT	16.763 32.691 16.795 32.755 ;
		RECT	16.427 32.691 16.459 32.755 ;
		RECT	16.091 32.691 16.123 32.755 ;
		RECT	15.755 32.691 15.787 32.755 ;
		RECT	15.419 32.691 15.451 32.755 ;
		RECT	15.083 32.691 15.115 32.755 ;
		RECT	14.747 32.691 14.779 32.755 ;
		RECT	14.411 32.691 14.443 32.755 ;
		RECT	26.507 32.691 26.539 32.755 ;
		RECT	14.075 32.691 14.107 32.755 ;
		RECT	13.739 32.691 13.771 32.755 ;
		RECT	13.403 32.691 13.435 32.755 ;
		RECT	13.067 32.691 13.099 32.755 ;
		RECT	12.731 32.691 12.763 32.755 ;
		RECT	12.395 32.691 12.427 32.755 ;
		RECT	12.059 32.691 12.091 32.755 ;
		RECT	11.723 32.691 11.755 32.755 ;
		RECT	11.387 32.691 11.419 32.755 ;
		RECT	11.051 32.691 11.083 32.755 ;
		RECT	26.171 32.691 26.203 32.755 ;
		RECT	10.715 32.691 10.747 32.755 ;
		RECT	10.379 32.691 10.411 32.755 ;
		RECT	10.043 32.691 10.075 32.755 ;
		RECT	9.707 32.691 9.739 32.755 ;
		RECT	9.371 32.691 9.403 32.755 ;
		RECT	9.035 32.691 9.067 32.755 ;
		RECT	8.699 32.691 8.731 32.755 ;
		RECT	8.363 32.691 8.395 32.755 ;
		RECT	8.027 32.691 8.059 32.755 ;
		RECT	7.691 32.691 7.723 32.755 ;
		RECT	25.835 32.691 25.867 32.755 ;
		RECT	7.355 32.691 7.387 32.755 ;
		RECT	7.019 32.691 7.051 32.755 ;
		RECT	6.683 32.691 6.715 32.755 ;
		RECT	6.347 32.691 6.379 32.755 ;
		RECT	25.499 32.691 25.531 32.755 ;
		RECT	25.163 32.691 25.195 32.755 ;
		RECT	24.827 32.691 24.859 32.755 ;
		RECT	24.491 32.691 24.523 32.755 ;
		RECT	43.68 43.125 43.712 43.157 ;
		RECT	42.672 43.125 42.704 43.157 ;
		RECT	41.328 43.125 41.36 43.157 ;
		RECT	40.32 43.125 40.352 43.157 ;
		RECT	38.64 43.125 38.672 43.157 ;
		RECT	38.304 43.125 38.336 43.157 ;
		RECT	36.96 43.125 36.992 43.157 ;
		RECT	35.952 43.125 35.984 43.157 ;
		RECT	49.056 44.026 49.088 44.09 ;
		RECT	45.36 44.026 45.392 44.09 ;
		RECT	31.92 44.026 31.952 44.09 ;
		RECT	30.576 44.026 30.608 44.09 ;
		RECT	28.56 44.026 28.592 44.09 ;
		RECT	5.793 44.026 5.825 44.09 ;
		RECT	49.311 32.691 49.375 32.755 ;
		RECT	49.704 39.399 49.736 39.431 ;
		RECT	49.531 41.87 49.563 41.902 ;
		RECT	49.641 42.425 49.673 42.457 ;
		RECT	49.921 43.431 49.953 43.495 ;
		RECT	49.327 44.026 49.359 44.09 ;
		RECT	27.557 44.026 27.589 44.09 ;
		RECT	27.221 44.026 27.253 44.09 ;
		RECT	24.197 44.026 24.229 44.09 ;
		RECT	23.861 44.026 23.893 44.09 ;
		RECT	23.525 44.026 23.557 44.09 ;
		RECT	23.189 44.026 23.221 44.09 ;
		RECT	22.853 44.026 22.885 44.09 ;
		RECT	22.517 44.026 22.549 44.09 ;
		RECT	22.181 44.026 22.213 44.09 ;
		RECT	21.845 44.026 21.877 44.09 ;
		RECT	21.509 44.026 21.541 44.09 ;
		RECT	21.173 44.026 21.205 44.09 ;
		RECT	26.885 44.026 26.917 44.09 ;
		RECT	20.837 44.026 20.869 44.09 ;
		RECT	20.501 44.026 20.533 44.09 ;
		RECT	20.165 44.026 20.197 44.09 ;
		RECT	19.829 44.026 19.861 44.09 ;
		RECT	19.493 44.026 19.525 44.09 ;
		RECT	19.157 44.026 19.189 44.09 ;
		RECT	18.821 44.026 18.853 44.09 ;
		RECT	18.485 44.026 18.517 44.09 ;
		RECT	18.149 44.026 18.181 44.09 ;
		RECT	17.813 44.026 17.845 44.09 ;
		RECT	26.549 44.026 26.581 44.09 ;
		RECT	17.477 44.026 17.509 44.09 ;
		RECT	17.141 44.026 17.173 44.09 ;
		RECT	16.805 44.026 16.837 44.09 ;
		RECT	16.469 44.026 16.501 44.09 ;
		RECT	16.133 44.026 16.165 44.09 ;
		RECT	15.797 44.026 15.829 44.09 ;
		RECT	15.461 44.026 15.493 44.09 ;
		RECT	15.125 44.026 15.157 44.09 ;
		RECT	14.789 44.026 14.821 44.09 ;
		RECT	14.453 44.026 14.485 44.09 ;
		RECT	26.213 44.026 26.245 44.09 ;
		RECT	14.117 44.026 14.149 44.09 ;
		RECT	13.781 44.026 13.813 44.09 ;
		RECT	13.445 44.026 13.477 44.09 ;
		RECT	13.109 44.026 13.141 44.09 ;
		RECT	12.773 44.026 12.805 44.09 ;
		RECT	12.437 44.026 12.469 44.09 ;
		RECT	12.101 44.026 12.133 44.09 ;
		RECT	11.765 44.026 11.797 44.09 ;
		RECT	11.429 44.026 11.461 44.09 ;
		RECT	11.093 44.026 11.125 44.09 ;
		RECT	25.877 44.026 25.909 44.09 ;
		RECT	10.757 44.026 10.789 44.09 ;
		RECT	10.421 44.026 10.453 44.09 ;
		RECT	10.085 44.026 10.117 44.09 ;
		RECT	9.749 44.026 9.781 44.09 ;
		RECT	9.413 44.026 9.445 44.09 ;
		RECT	9.077 44.026 9.109 44.09 ;
		RECT	8.741 44.026 8.773 44.09 ;
		RECT	8.405 44.026 8.437 44.09 ;
		RECT	8.069 44.026 8.101 44.09 ;
		RECT	7.733 44.026 7.765 44.09 ;
		RECT	25.541 44.026 25.573 44.09 ;
		RECT	7.397 44.026 7.429 44.09 ;
		RECT	7.061 44.026 7.093 44.09 ;
		RECT	6.725 44.026 6.757 44.09 ;
		RECT	25.205 44.026 25.237 44.09 ;
		RECT	24.869 44.026 24.901 44.09 ;
		RECT	24.533 44.026 24.565 44.09 ;
		RECT	48.767 33.488 48.799 33.552 ;
		RECT	28.271 33.488 28.303 33.552 ;
		RECT	49.103 33.65 49.135 33.714 ;
		RECT	27.935 33.65 27.967 33.714 ;
		RECT	48.095 33.896 48.127 33.928 ;
		RECT	48.767 34.641 48.799 34.673 ;
		RECT	28.271 34.641 28.303 34.673 ;
		RECT	49.103 34.721 49.135 34.753 ;
		RECT	27.935 34.721 27.967 34.753 ;
		RECT	44.352 39.158 44.384 39.19 ;
		RECT	38.976 39.158 39.008 39.19 ;
		RECT	35.616 39.158 35.648 39.19 ;
		RECT	33.6 39.158 33.632 39.19 ;
		RECT	28.224 39.158 28.256 39.19 ;
		RECT	49.091 39.187 49.123 39.251 ;
		RECT	48.52 39.187 48.584 39.251 ;
		RECT	48.384 39.187 48.416 39.251 ;
		RECT	47.04 39.187 47.072 39.251 ;
		RECT	46.368 39.187 46.4 39.251 ;
		RECT	45.024 39.258 45.056 39.29 ;
		RECT	39.312 39.258 39.344 39.29 ;
		RECT	36.288 39.258 36.32 39.29 ;
		RECT	33.936 39.258 33.968 39.29 ;
		RECT	28.896 39.258 28.928 39.29 ;
		RECT	45.696 39.358 45.728 39.39 ;
		RECT	36.624 39.358 36.656 39.39 ;
		RECT	34.944 39.358 34.976 39.39 ;
		RECT	29.568 39.358 29.6 39.39 ;
		RECT	49.091 39.413 49.123 39.477 ;
		RECT	48.52 39.413 48.584 39.477 ;
		RECT	48.384 39.413 48.416 39.477 ;
		RECT	46.368 39.458 46.4 39.49 ;
		RECT	36.96 39.458 36.992 39.49 ;
		RECT	35.616 39.458 35.648 39.49 ;
		RECT	30.24 39.458 30.272 39.49 ;
		RECT	47.04 39.558 47.072 39.59 ;
		RECT	41.664 39.558 41.696 39.59 ;
		RECT	39.984 39.558 40.016 39.59 ;
		RECT	36.288 39.558 36.32 39.59 ;
		RECT	30.912 39.558 30.944 39.59 ;
		RECT	47.376 39.658 47.408 39.69 ;
		RECT	42 39.658 42.032 39.69 ;
		RECT	40.32 39.658 40.352 39.69 ;
		RECT	36.96 39.658 36.992 39.69 ;
		RECT	31.584 39.658 31.616 39.69 ;
		RECT	48.384 39.758 48.416 39.79 ;
		RECT	43.008 39.758 43.04 39.79 ;
		RECT	40.656 39.758 40.688 39.79 ;
		RECT	37.632 39.758 37.664 39.79 ;
		RECT	32.256 39.758 32.288 39.79 ;
		RECT	49.091 39.858 49.123 39.89 ;
		RECT	43.68 39.858 43.712 39.89 ;
		RECT	40.992 39.858 41.024 39.89 ;
		RECT	37.968 39.858 38 39.89 ;
		RECT	32.928 39.858 32.96 39.89 ;
		RECT	48.384 41.87 48.416 41.902 ;
		RECT	47.04 42.425 47.072 42.457 ;
		RECT	41.664 42.425 41.696 42.457 ;
		RECT	48.52 42.454 48.584 42.518 ;
		RECT	40.656 42.525 40.688 42.557 ;
		RECT	39.984 42.625 40.016 42.657 ;
		RECT	35.28 42.625 35.312 42.657 ;
		RECT	43.68 42.649 43.712 42.713 ;
		RECT	42.672 42.649 42.704 42.713 ;
		RECT	41.328 42.649 41.36 42.713 ;
		RECT	48.52 42.659 48.584 42.723 ;
		RECT	47.04 42.659 47.072 42.723 ;
		RECT	46.032 42.659 46.064 42.723 ;
		RECT	39.312 42.725 39.344 42.757 ;
		RECT	32.592 42.725 32.624 42.757 ;
		RECT	37.964 42.825 37.996 42.857 ;
		RECT	43.68 42.854 43.712 42.918 ;
		RECT	42.672 42.854 42.704 42.918 ;
		RECT	41.328 42.854 41.36 42.918 ;
		RECT	40.32 42.854 40.352 42.918 ;
		RECT	38.64 42.859 38.672 42.923 ;
		RECT	38.304 42.859 38.336 42.923 ;
		RECT	48.52 42.864 48.584 42.928 ;
		RECT	47.04 42.864 47.072 42.928 ;
		RECT	46.032 42.864 46.064 42.928 ;
		RECT	37.628 42.925 37.66 42.957 ;
		RECT	45.024 43.025 45.056 43.057 ;
		RECT	44.352 43.025 44.384 43.057 ;
		RECT	43.344 43.025 43.376 43.057 ;
		RECT	43.008 43.025 43.04 43.057 ;
		RECT	42.336 43.025 42.368 43.057 ;
		RECT	42 43.025 42.032 43.057 ;
		RECT	40.992 43.025 41.024 43.057 ;
		RECT	39.648 43.025 39.68 43.057 ;
		RECT	38.976 43.025 39.008 43.057 ;
		RECT	36.624 43.025 36.656 43.057 ;
		RECT	36.284 43.025 36.316 43.057 ;
		RECT	48.536 43.069 48.568 43.133 ;
		RECT	47.04 43.069 47.072 43.133 ;
		RECT	46.032 43.069 46.064 43.133 ;
		RECT	45.36 43.125 45.392 43.157 ;
		RECT	44.688 43.125 44.72 43.157 ;
		RECT	44.016 43.125 44.048 43.157 ;
		RECT	37.296 43.125 37.328 43.157 ;
		RECT	35.616 43.125 35.648 43.157 ;
		RECT	35.276 43.125 35.308 43.157 ;
		RECT	48.536 44.026 48.568 44.09 ;
		RECT	47.04 44.026 47.072 44.09 ;
		RECT	46.032 44.026 46.064 44.09 ;
		RECT	43.68 44.026 43.712 44.09 ;
		RECT	42.672 44.026 42.704 44.09 ;
		RECT	41.328 44.026 41.36 44.09 ;
		RECT	40.32 44.026 40.352 44.09 ;
		RECT	39.648 44.026 39.68 44.09 ;
		RECT	38.64 44.026 38.672 44.09 ;
		RECT	38.304 44.026 38.336 44.09 ;
		RECT	37.296 44.026 37.328 44.09 ;
		RECT	36.96 44.026 36.992 44.09 ;
		RECT	35.952 44.026 35.984 44.09 ;
		RECT	35.616 44.026 35.648 44.09 ;
		RECT	34.608 44.026 34.64 44.09 ;
		RECT	34.272 44.026 34.304 44.09 ;
		RECT	32.592 44.026 32.624 44.09 ;
		RECT	31.584 44.026 31.616 44.09 ;
		RECT	30.912 44.026 30.944 44.09 ;
		RECT	30.24 44.026 30.272 44.09 ;
		RECT	29.904 44.026 29.936 44.09 ;
		RECT	29.568 44.026 29.6 44.09 ;
		RECT	29.232 44.026 29.264 44.09 ;
		RECT	27.888 44.026 27.92 44.09 ;
		RECT	5.789 43.431 5.821 43.495 ;
		RECT	6.389 44.026 6.421 44.09 ;
		RECT	102.626 31.762 102.69 31.794 ;
		RECT	102.626 50.382 102.69 50.414 ;
		RECT	80.615 39.858 80.647 39.89 ;
		RECT	83.975 39.358 84.007 39.39 ;
		RECT	84.311 39.358 84.343 39.39 ;
		RECT	84.647 39.258 84.679 39.29 ;
		RECT	84.983 39.258 85.015 39.29 ;
		RECT	85.319 39.158 85.351 39.19 ;
		RECT	85.655 39.158 85.687 39.19 ;
		RECT	85.991 39.858 86.023 39.89 ;
		RECT	86.327 39.858 86.359 39.89 ;
		RECT	86.663 39.758 86.695 39.79 ;
		RECT	86.999 39.758 87.031 39.79 ;
		RECT	80.951 39.858 80.983 39.89 ;
		RECT	87.335 39.658 87.367 39.69 ;
		RECT	87.671 39.658 87.703 39.69 ;
		RECT	88.007 39.558 88.039 39.59 ;
		RECT	88.343 39.558 88.375 39.59 ;
		RECT	88.679 39.458 88.711 39.49 ;
		RECT	89.015 39.458 89.047 39.49 ;
		RECT	89.351 39.358 89.383 39.39 ;
		RECT	89.687 39.358 89.719 39.39 ;
		RECT	90.023 39.258 90.055 39.29 ;
		RECT	90.359 39.258 90.391 39.29 ;
		RECT	81.287 39.758 81.319 39.79 ;
		RECT	90.695 39.158 90.727 39.19 ;
		RECT	91.031 39.158 91.063 39.19 ;
		RECT	91.367 39.858 91.399 39.89 ;
		RECT	91.703 39.858 91.735 39.89 ;
		RECT	92.039 39.758 92.071 39.79 ;
		RECT	92.375 39.758 92.407 39.79 ;
		RECT	92.711 39.658 92.743 39.69 ;
		RECT	93.047 39.658 93.079 39.69 ;
		RECT	93.383 39.558 93.415 39.59 ;
		RECT	93.719 39.558 93.751 39.59 ;
		RECT	81.623 39.758 81.655 39.79 ;
		RECT	94.055 39.458 94.087 39.49 ;
		RECT	94.391 39.458 94.423 39.49 ;
		RECT	94.727 39.358 94.759 39.39 ;
		RECT	95.063 39.358 95.095 39.39 ;
		RECT	95.399 39.258 95.431 39.29 ;
		RECT	95.735 39.258 95.767 39.29 ;
		RECT	96.071 39.158 96.103 39.19 ;
		RECT	96.407 39.158 96.439 39.19 ;
		RECT	96.743 39.858 96.775 39.89 ;
		RECT	97.079 39.858 97.111 39.89 ;
		RECT	81.959 39.658 81.991 39.69 ;
		RECT	97.415 39.758 97.447 39.79 ;
		RECT	97.751 39.758 97.783 39.79 ;
		RECT	98.087 39.658 98.119 39.69 ;
		RECT	98.423 39.658 98.455 39.69 ;
		RECT	98.759 39.558 98.791 39.59 ;
		RECT	99.095 39.558 99.127 39.59 ;
		RECT	99.431 39.458 99.463 39.49 ;
		RECT	99.767 39.458 99.799 39.49 ;
		RECT	100.103 39.358 100.135 39.39 ;
		RECT	100.439 39.358 100.471 39.39 ;
		RECT	82.295 39.658 82.327 39.69 ;
		RECT	100.775 39.258 100.807 39.29 ;
		RECT	101.111 39.258 101.143 39.29 ;
		RECT	101.447 39.158 101.479 39.19 ;
		RECT	101.783 39.158 101.815 39.19 ;
		RECT	82.631 39.558 82.663 39.59 ;
		RECT	82.967 39.558 82.999 39.59 ;
		RECT	83.303 39.458 83.335 39.49 ;
		RECT	83.639 39.458 83.671 39.49 ;
		RECT	80.615 42.825 80.647 42.857 ;
		RECT	83.975 42.825 84.007 42.857 ;
		RECT	84.311 42.825 84.343 42.857 ;
		RECT	84.647 42.825 84.679 42.857 ;
		RECT	84.983 42.825 85.015 42.857 ;
		RECT	85.319 42.825 85.351 42.857 ;
		RECT	85.655 42.825 85.687 42.857 ;
		RECT	85.991 42.925 86.023 42.957 ;
		RECT	86.327 42.925 86.359 42.957 ;
		RECT	86.663 42.925 86.695 42.957 ;
		RECT	86.999 42.925 87.031 42.957 ;
		RECT	80.951 42.825 80.983 42.857 ;
		RECT	87.335 42.925 87.367 42.957 ;
		RECT	87.671 42.925 87.703 42.957 ;
		RECT	88.007 42.925 88.039 42.957 ;
		RECT	88.343 42.925 88.375 42.957 ;
		RECT	88.679 42.925 88.711 42.957 ;
		RECT	89.015 42.925 89.047 42.957 ;
		RECT	89.351 42.925 89.383 42.957 ;
		RECT	89.687 42.925 89.719 42.957 ;
		RECT	90.023 42.925 90.055 42.957 ;
		RECT	90.359 42.925 90.391 42.957 ;
		RECT	81.287 42.825 81.319 42.857 ;
		RECT	90.695 42.925 90.727 42.957 ;
		RECT	91.031 42.925 91.063 42.957 ;
		RECT	91.367 43.025 91.399 43.057 ;
		RECT	91.703 43.025 91.735 43.057 ;
		RECT	92.039 43.025 92.071 43.057 ;
		RECT	92.375 43.025 92.407 43.057 ;
		RECT	92.711 43.025 92.743 43.057 ;
		RECT	93.047 43.025 93.079 43.057 ;
		RECT	93.383 43.025 93.415 43.057 ;
		RECT	93.719 43.025 93.751 43.057 ;
		RECT	81.623 42.825 81.655 42.857 ;
		RECT	94.055 43.025 94.087 43.057 ;
		RECT	94.391 43.025 94.423 43.057 ;
		RECT	94.727 43.025 94.759 43.057 ;
		RECT	95.063 43.025 95.095 43.057 ;
		RECT	95.399 43.025 95.431 43.057 ;
		RECT	95.735 43.025 95.767 43.057 ;
		RECT	96.071 43.025 96.103 43.057 ;
		RECT	96.407 43.025 96.439 43.057 ;
		RECT	96.743 43.125 96.775 43.157 ;
		RECT	97.079 43.125 97.111 43.157 ;
		RECT	81.959 42.825 81.991 42.857 ;
		RECT	97.415 43.125 97.447 43.157 ;
		RECT	97.751 43.125 97.783 43.157 ;
		RECT	98.087 43.125 98.119 43.157 ;
		RECT	98.423 43.125 98.455 43.157 ;
		RECT	98.759 43.125 98.791 43.157 ;
		RECT	99.095 43.125 99.127 43.157 ;
		RECT	99.431 43.125 99.463 43.157 ;
		RECT	99.767 43.125 99.799 43.157 ;
		RECT	100.103 43.125 100.135 43.157 ;
		RECT	100.439 43.125 100.471 43.157 ;
		RECT	82.295 42.825 82.327 42.857 ;
		RECT	100.775 43.125 100.807 43.157 ;
		RECT	101.111 43.125 101.143 43.157 ;
		RECT	101.447 43.125 101.479 43.157 ;
		RECT	101.783 43.125 101.815 43.157 ;
		RECT	82.631 42.825 82.663 42.857 ;
		RECT	82.967 42.825 82.999 42.857 ;
		RECT	83.303 42.825 83.335 42.857 ;
		RECT	83.639 42.825 83.671 42.857 ;
		RECT	80.657 32.691 80.689 32.755 ;
		RECT	58.461 39.672 58.493 39.736 ;
		RECT	58.497 44.026 58.529 44.09 ;
		RECT	84.017 32.691 84.049 32.755 ;
		RECT	84.353 32.691 84.385 32.755 ;
		RECT	84.689 32.691 84.721 32.755 ;
		RECT	85.025 32.691 85.057 32.755 ;
		RECT	85.361 32.691 85.393 32.755 ;
		RECT	85.697 32.691 85.729 32.755 ;
		RECT	86.033 32.691 86.065 32.755 ;
		RECT	86.369 32.691 86.401 32.755 ;
		RECT	86.705 32.691 86.737 32.755 ;
		RECT	87.041 32.691 87.073 32.755 ;
		RECT	80.993 32.691 81.025 32.755 ;
		RECT	87.377 32.691 87.409 32.755 ;
		RECT	87.713 32.691 87.745 32.755 ;
		RECT	88.049 32.691 88.081 32.755 ;
		RECT	88.385 32.691 88.417 32.755 ;
		RECT	88.721 32.691 88.753 32.755 ;
		RECT	89.057 32.691 89.089 32.755 ;
		RECT	89.393 32.691 89.425 32.755 ;
		RECT	89.729 32.691 89.761 32.755 ;
		RECT	90.065 32.691 90.097 32.755 ;
		RECT	90.401 32.691 90.433 32.755 ;
		RECT	81.329 32.691 81.361 32.755 ;
		RECT	90.737 32.691 90.769 32.755 ;
		RECT	91.073 32.691 91.105 32.755 ;
		RECT	91.409 32.691 91.441 32.755 ;
		RECT	91.745 32.691 91.777 32.755 ;
		RECT	92.081 32.691 92.113 32.755 ;
		RECT	92.417 32.691 92.449 32.755 ;
		RECT	92.753 32.691 92.785 32.755 ;
		RECT	93.089 32.691 93.121 32.755 ;
		RECT	93.425 32.691 93.457 32.755 ;
		RECT	93.761 32.691 93.793 32.755 ;
		RECT	81.665 32.691 81.697 32.755 ;
		RECT	94.097 32.691 94.129 32.755 ;
		RECT	94.433 32.691 94.465 32.755 ;
		RECT	94.769 32.691 94.801 32.755 ;
		RECT	95.105 32.691 95.137 32.755 ;
		RECT	95.441 32.691 95.473 32.755 ;
		RECT	95.777 32.691 95.809 32.755 ;
		RECT	96.113 32.691 96.145 32.755 ;
		RECT	96.449 32.691 96.481 32.755 ;
		RECT	96.785 32.691 96.817 32.755 ;
		RECT	97.121 32.691 97.153 32.755 ;
		RECT	82.001 32.691 82.033 32.755 ;
		RECT	97.457 32.691 97.489 32.755 ;
		RECT	97.793 32.691 97.825 32.755 ;
		RECT	98.129 32.691 98.161 32.755 ;
		RECT	98.465 32.691 98.497 32.755 ;
		RECT	98.801 32.691 98.833 32.755 ;
		RECT	99.137 32.691 99.169 32.755 ;
		RECT	99.473 32.691 99.505 32.755 ;
		RECT	99.809 32.691 99.841 32.755 ;
		RECT	100.145 32.691 100.177 32.755 ;
		RECT	100.481 32.691 100.513 32.755 ;
		RECT	82.337 32.691 82.369 32.755 ;
		RECT	100.817 32.691 100.849 32.755 ;
		RECT	101.153 32.691 101.185 32.755 ;
		RECT	101.489 32.691 101.521 32.755 ;
		RECT	101.825 32.691 101.857 32.755 ;
		RECT	82.673 32.691 82.705 32.755 ;
		RECT	83.009 32.691 83.041 32.755 ;
		RECT	83.345 32.691 83.377 32.755 ;
		RECT	83.681 32.691 83.713 32.755 ;
		RECT	64.492 43.125 64.524 43.157 ;
		RECT	65.5 43.125 65.532 43.157 ;
		RECT	66.844 43.125 66.876 43.157 ;
		RECT	67.852 43.125 67.884 43.157 ;
		RECT	69.532 43.125 69.564 43.157 ;
		RECT	69.868 43.125 69.9 43.157 ;
		RECT	71.212 43.125 71.244 43.157 ;
		RECT	72.22 43.125 72.252 43.157 ;
		RECT	59.116 44.026 59.148 44.09 ;
		RECT	62.812 44.026 62.844 44.09 ;
		RECT	76.252 44.026 76.284 44.09 ;
		RECT	77.596 44.026 77.628 44.09 ;
		RECT	79.612 44.026 79.644 44.09 ;
		RECT	102.379 44.026 102.411 44.09 ;
		RECT	58.829 32.691 58.893 32.755 ;
		RECT	58.468 39.399 58.5 39.431 ;
		RECT	58.641 41.87 58.673 41.902 ;
		RECT	58.531 42.425 58.563 42.457 ;
		RECT	58.251 43.431 58.283 43.495 ;
		RECT	58.845 44.026 58.877 44.09 ;
		RECT	80.615 44.026 80.647 44.09 ;
		RECT	80.951 44.026 80.983 44.09 ;
		RECT	83.975 44.026 84.007 44.09 ;
		RECT	84.311 44.026 84.343 44.09 ;
		RECT	84.647 44.026 84.679 44.09 ;
		RECT	84.983 44.026 85.015 44.09 ;
		RECT	85.319 44.026 85.351 44.09 ;
		RECT	85.655 44.026 85.687 44.09 ;
		RECT	85.991 44.026 86.023 44.09 ;
		RECT	86.327 44.026 86.359 44.09 ;
		RECT	86.663 44.026 86.695 44.09 ;
		RECT	86.999 44.026 87.031 44.09 ;
		RECT	81.287 44.026 81.319 44.09 ;
		RECT	87.335 44.026 87.367 44.09 ;
		RECT	87.671 44.026 87.703 44.09 ;
		RECT	88.007 44.026 88.039 44.09 ;
		RECT	88.343 44.026 88.375 44.09 ;
		RECT	88.679 44.026 88.711 44.09 ;
		RECT	89.015 44.026 89.047 44.09 ;
		RECT	89.351 44.026 89.383 44.09 ;
		RECT	89.687 44.026 89.719 44.09 ;
		RECT	90.023 44.026 90.055 44.09 ;
		RECT	90.359 44.026 90.391 44.09 ;
		RECT	81.623 44.026 81.655 44.09 ;
		RECT	90.695 44.026 90.727 44.09 ;
		RECT	91.031 44.026 91.063 44.09 ;
		RECT	91.367 44.026 91.399 44.09 ;
		RECT	91.703 44.026 91.735 44.09 ;
		RECT	92.039 44.026 92.071 44.09 ;
		RECT	92.375 44.026 92.407 44.09 ;
		RECT	92.711 44.026 92.743 44.09 ;
		RECT	93.047 44.026 93.079 44.09 ;
		RECT	93.383 44.026 93.415 44.09 ;
		RECT	93.719 44.026 93.751 44.09 ;
		RECT	81.959 44.026 81.991 44.09 ;
		RECT	94.055 44.026 94.087 44.09 ;
		RECT	94.391 44.026 94.423 44.09 ;
		RECT	94.727 44.026 94.759 44.09 ;
		RECT	95.063 44.026 95.095 44.09 ;
		RECT	95.399 44.026 95.431 44.09 ;
		RECT	95.735 44.026 95.767 44.09 ;
		RECT	96.071 44.026 96.103 44.09 ;
		RECT	96.407 44.026 96.439 44.09 ;
		RECT	96.743 44.026 96.775 44.09 ;
		RECT	97.079 44.026 97.111 44.09 ;
		RECT	82.295 44.026 82.327 44.09 ;
		RECT	97.415 44.026 97.447 44.09 ;
		RECT	97.751 44.026 97.783 44.09 ;
		RECT	98.087 44.026 98.119 44.09 ;
		RECT	98.423 44.026 98.455 44.09 ;
		RECT	98.759 44.026 98.791 44.09 ;
		RECT	99.095 44.026 99.127 44.09 ;
		RECT	99.431 44.026 99.463 44.09 ;
		RECT	99.767 44.026 99.799 44.09 ;
		RECT	100.103 44.026 100.135 44.09 ;
		RECT	100.439 44.026 100.471 44.09 ;
		RECT	82.631 44.026 82.663 44.09 ;
		RECT	100.775 44.026 100.807 44.09 ;
		RECT	101.111 44.026 101.143 44.09 ;
		RECT	101.447 44.026 101.479 44.09 ;
		RECT	82.967 44.026 82.999 44.09 ;
		RECT	83.303 44.026 83.335 44.09 ;
		RECT	83.639 44.026 83.671 44.09 ;
		RECT	59.405 33.488 59.437 33.552 ;
		RECT	79.901 33.488 79.933 33.552 ;
		RECT	59.069 33.65 59.101 33.714 ;
		RECT	80.237 33.65 80.269 33.714 ;
		RECT	60.077 33.896 60.109 33.928 ;
		RECT	59.405 34.641 59.437 34.673 ;
		RECT	79.901 34.641 79.933 34.673 ;
		RECT	59.069 34.721 59.101 34.753 ;
		RECT	80.237 34.721 80.269 34.753 ;
		RECT	63.82 39.158 63.852 39.19 ;
		RECT	69.196 39.158 69.228 39.19 ;
		RECT	72.556 39.158 72.588 39.19 ;
		RECT	74.572 39.158 74.604 39.19 ;
		RECT	79.948 39.158 79.98 39.19 ;
		RECT	59.081 39.187 59.113 39.251 ;
		RECT	59.62 39.187 59.684 39.251 ;
		RECT	59.788 39.187 59.82 39.251 ;
		RECT	61.132 39.187 61.164 39.251 ;
		RECT	61.804 39.187 61.836 39.251 ;
		RECT	63.148 39.258 63.18 39.29 ;
		RECT	68.86 39.258 68.892 39.29 ;
		RECT	71.884 39.258 71.916 39.29 ;
		RECT	74.236 39.258 74.268 39.29 ;
		RECT	79.276 39.258 79.308 39.29 ;
		RECT	62.476 39.358 62.508 39.39 ;
		RECT	71.548 39.358 71.58 39.39 ;
		RECT	73.228 39.358 73.26 39.39 ;
		RECT	78.604 39.358 78.636 39.39 ;
		RECT	59.081 39.413 59.113 39.477 ;
		RECT	59.62 39.413 59.684 39.477 ;
		RECT	59.788 39.413 59.82 39.477 ;
		RECT	61.804 39.458 61.836 39.49 ;
		RECT	71.212 39.458 71.244 39.49 ;
		RECT	72.556 39.458 72.588 39.49 ;
		RECT	77.932 39.458 77.964 39.49 ;
		RECT	61.132 39.558 61.164 39.59 ;
		RECT	66.508 39.558 66.54 39.59 ;
		RECT	68.188 39.558 68.22 39.59 ;
		RECT	71.884 39.558 71.916 39.59 ;
		RECT	77.26 39.558 77.292 39.59 ;
		RECT	60.796 39.658 60.828 39.69 ;
		RECT	66.172 39.658 66.204 39.69 ;
		RECT	67.852 39.658 67.884 39.69 ;
		RECT	71.212 39.658 71.244 39.69 ;
		RECT	76.588 39.658 76.62 39.69 ;
		RECT	59.788 39.758 59.82 39.79 ;
		RECT	65.164 39.758 65.196 39.79 ;
		RECT	67.516 39.758 67.548 39.79 ;
		RECT	70.54 39.758 70.572 39.79 ;
		RECT	75.916 39.758 75.948 39.79 ;
		RECT	59.081 39.858 59.113 39.89 ;
		RECT	64.492 39.858 64.524 39.89 ;
		RECT	67.18 39.858 67.212 39.89 ;
		RECT	70.204 39.858 70.236 39.89 ;
		RECT	75.244 39.858 75.276 39.89 ;
		RECT	59.788 41.87 59.82 41.902 ;
		RECT	61.132 42.425 61.164 42.457 ;
		RECT	66.508 42.425 66.54 42.457 ;
		RECT	59.62 42.454 59.684 42.518 ;
		RECT	67.516 42.525 67.548 42.557 ;
		RECT	68.188 42.625 68.22 42.657 ;
		RECT	72.892 42.625 72.924 42.657 ;
		RECT	64.492 42.649 64.524 42.713 ;
		RECT	65.5 42.649 65.532 42.713 ;
		RECT	66.844 42.649 66.876 42.713 ;
		RECT	59.62 42.659 59.684 42.723 ;
		RECT	61.132 42.659 61.164 42.723 ;
		RECT	62.14 42.659 62.172 42.723 ;
		RECT	68.86 42.725 68.892 42.757 ;
		RECT	75.58 42.725 75.612 42.757 ;
		RECT	70.208 42.825 70.24 42.857 ;
		RECT	64.492 42.854 64.524 42.918 ;
		RECT	65.5 42.854 65.532 42.918 ;
		RECT	66.844 42.854 66.876 42.918 ;
		RECT	67.852 42.854 67.884 42.918 ;
		RECT	69.532 42.859 69.564 42.923 ;
		RECT	69.868 42.859 69.9 42.923 ;
		RECT	59.62 42.864 59.684 42.928 ;
		RECT	61.132 42.864 61.164 42.928 ;
		RECT	62.14 42.864 62.172 42.928 ;
		RECT	70.544 42.925 70.576 42.957 ;
		RECT	63.148 43.025 63.18 43.057 ;
		RECT	63.82 43.025 63.852 43.057 ;
		RECT	64.828 43.025 64.86 43.057 ;
		RECT	65.164 43.025 65.196 43.057 ;
		RECT	65.836 43.025 65.868 43.057 ;
		RECT	66.172 43.025 66.204 43.057 ;
		RECT	67.18 43.025 67.212 43.057 ;
		RECT	68.524 43.025 68.556 43.057 ;
		RECT	69.196 43.025 69.228 43.057 ;
		RECT	71.548 43.025 71.58 43.057 ;
		RECT	71.888 43.025 71.92 43.057 ;
		RECT	59.636 43.069 59.668 43.133 ;
		RECT	61.132 43.069 61.164 43.133 ;
		RECT	62.14 43.069 62.172 43.133 ;
		RECT	62.812 43.125 62.844 43.157 ;
		RECT	63.484 43.125 63.516 43.157 ;
		RECT	64.156 43.125 64.188 43.157 ;
		RECT	70.876 43.125 70.908 43.157 ;
		RECT	72.556 43.125 72.588 43.157 ;
		RECT	72.896 43.125 72.928 43.157 ;
		RECT	59.636 44.026 59.668 44.09 ;
		RECT	61.132 44.026 61.164 44.09 ;
		RECT	62.14 44.026 62.172 44.09 ;
		RECT	64.492 44.026 64.524 44.09 ;
		RECT	65.5 44.026 65.532 44.09 ;
		RECT	66.844 44.026 66.876 44.09 ;
		RECT	67.852 44.026 67.884 44.09 ;
		RECT	68.524 44.026 68.556 44.09 ;
		RECT	69.532 44.026 69.564 44.09 ;
		RECT	69.868 44.026 69.9 44.09 ;
		RECT	70.876 44.026 70.908 44.09 ;
		RECT	71.212 44.026 71.244 44.09 ;
		RECT	72.22 44.026 72.252 44.09 ;
		RECT	72.556 44.026 72.588 44.09 ;
		RECT	73.564 44.026 73.596 44.09 ;
		RECT	73.9 44.026 73.932 44.09 ;
		RECT	75.58 44.026 75.612 44.09 ;
		RECT	76.588 44.026 76.62 44.09 ;
		RECT	77.26 44.026 77.292 44.09 ;
		RECT	77.932 44.026 77.964 44.09 ;
		RECT	78.268 44.026 78.3 44.09 ;
		RECT	78.604 44.026 78.636 44.09 ;
		RECT	78.94 44.026 78.972 44.09 ;
		RECT	80.284 44.026 80.316 44.09 ;
		RECT	102.383 43.431 102.415 43.495 ;
		RECT	101.783 44.026 101.815 44.09 ;
		RECT	150.001 33.796 150.033 33.828 ;
		RECT	150.122 32.691 150.154 32.755 ;
		RECT	150.576 32.691 150.608 32.755 ;
		RECT	150.966 32.691 151.03 32.755 ;
		RECT	152.249 32.691 152.281 32.755 ;
		RECT	153.56 32.691 153.624 32.755 ;
		RECT	153.801 32.691 153.833 32.755 ;
		RECT	152.957 32.876 152.989 32.94 ;
		RECT	148.328 33.437 148.36 33.469 ;
		RECT	155.929 33.437 155.961 33.469 ;
		RECT	150.076 33.701 150.108 33.733 ;
		RECT	152.961 33.701 152.993 33.733 ;
		RECT	152.277 34.641 152.309 34.673 ;
		RECT	153.456 34.721 153.488 34.753 ;
		RECT	151.243 34.801 151.275 34.833 ;
		RECT	150.452 34.896 150.484 34.928 ;
		RECT	148.586 35.948 148.618 35.98 ;
		RECT	150.289 36.454 150.321 36.486 ;
		RECT	152.357 36.454 152.389 36.486 ;
		RECT	155.836 36.454 155.868 36.486 ;
		RECT	151.103 37.589 151.135 37.621 ;
		RECT	149.884 37.689 149.916 37.721 ;
		RECT	150.148 38.361 150.18 38.393 ;
		RECT	151.102 38.651 151.134 38.683 ;
		RECT	149.918 39.191 149.95 39.255 ;
		RECT	148.415 39.192 148.479 39.256 ;
		RECT	149.272 39.192 149.304 39.256 ;
		RECT	151.908 39.192 151.94 39.256 ;
		RECT	152.361 39.192 152.425 39.256 ;
		RECT	152.81 39.192 152.842 39.256 ;
		RECT	153.206 39.192 153.27 39.256 ;
		RECT	153.56 39.192 153.624 39.256 ;
		RECT	153.967 39.192 154.031 39.256 ;
		RECT	155.361 39.192 155.393 39.256 ;
		RECT	154.142 39.193 154.174 39.257 ;
		RECT	153.033 39.399 153.065 39.431 ;
		RECT	150.966 39.672 151.03 39.736 ;
		RECT	153.526 39.672 153.59 39.736 ;
		RECT	154.662 39.672 154.694 39.736 ;
		RECT	155.507 39.672 155.571 39.736 ;
		RECT	152.135 39.853 152.167 39.885 ;
		RECT	155.508 39.853 155.54 39.885 ;
		RECT	150.148 40.363 150.18 40.395 ;
		RECT	148.328 40.458 148.36 40.49 ;
		RECT	150.219 40.538 150.251 40.57 ;
		RECT	153.874 40.618 153.906 40.65 ;
		RECT	150.148 40.903 150.18 40.935 ;
		RECT	152.063 41.53 152.095 41.562 ;
		RECT	153.808 41.53 153.84 41.562 ;
		RECT	150.076 41.87 150.108 41.902 ;
		RECT	152.063 41.87 152.095 41.902 ;
		RECT	151.102 41.97 151.134 42.002 ;
		RECT	148.66 42.425 148.692 42.457 ;
		RECT	150.289 42.425 150.321 42.457 ;
		RECT	150.452 42.425 150.484 42.457 ;
		RECT	152.357 42.425 152.389 42.457 ;
		RECT	153.808 42.425 153.84 42.457 ;
		RECT	150.219 42.52 150.251 42.552 ;
		RECT	155.251 42.52 155.283 42.552 ;
		RECT	148.656 42.659 148.688 42.723 ;
		RECT	150.966 42.675 151.03 42.707 ;
		RECT	152.249 42.675 152.281 42.707 ;
		RECT	153.56 42.675 153.624 42.707 ;
		RECT	148.656 42.864 148.688 42.928 ;
		RECT	150.966 42.864 151.03 42.928 ;
		RECT	152.249 42.864 152.281 42.928 ;
		RECT	153.56 42.864 153.624 42.928 ;
		RECT	148.656 43.069 148.688 43.133 ;
		RECT	152.249 43.069 152.281 43.133 ;
		RECT	150.966 43.085 151.03 43.117 ;
		RECT	153.56 43.085 153.624 43.117 ;
		RECT	150.452 43.467 150.484 43.499 ;
		RECT	150.024 44.026 150.056 44.09 ;
		RECT	152.249 44.026 152.281 44.09 ;
		RECT	153.84 44.026 153.872 44.09 ;
		RECT	150.966 44.042 151.03 44.074 ;
		RECT	153.56 44.042 153.624 44.074 ;
		RECT	150.128 44.199 150.16 44.231 ;
		RECT	151.102 44.469 151.134 44.501 ;
		RECT	151.102 44.759 151.134 44.791 ;
		RECT	148.656 45.197 148.688 45.229 ;
		RECT	151.243 45.197 151.275 45.229 ;
		RECT	151.092 46.057 151.124 46.089 ;
		RECT	151.093 46.632 151.125 46.664 ;
		RECT	148.555 47.367 148.587 47.399 ;
		RECT	150.275 47.467 150.307 47.499 ;
		RECT	152.357 47.467 152.389 47.499 ;
		RECT	150.452 48.217 150.484 48.249 ;
		RECT	148.33 48.317 148.362 48.349 ;
		RECT	150.045 49.263 150.077 49.327 ;
		RECT	152.733 50.027 152.765 50.059 ;
		RECT	151.995 34.896 152.027 34.928 ;
		RECT	155.367 43.467 155.399 43.499 ;
		RECT	150.148 37.474 150.18 37.506 ;
		RECT	153.46 47.367 153.492 47.399 ;
		RECT	151.102 41.004 151.134 41.036 ;
		RECT	153.526 36.238 153.558 36.27 ;
		RECT	150.148 39.192 150.18 39.256 ;
		RECT	150.452 39.192 150.484 39.256 ;
		RECT	150.966 39.192 151.03 39.256 ;
		RECT	154.662 39.192 154.694 39.256 ;
		RECT	148.415 39.672 148.479 39.736 ;
		RECT	149.272 39.672 149.304 39.736 ;
		RECT	149.918 39.672 149.95 39.736 ;
		RECT	151.892 39.672 151.924 39.736 ;
		RECT	152.361 39.672 152.425 39.736 ;
		RECT	152.802 39.672 152.834 39.736 ;
		RECT	153.967 39.672 154.031 39.736 ;
		RECT	154.142 39.672 154.174 39.736 ;
		RECT	155.361 39.672 155.393 39.736 ;
		RECT	149.918 42.659 149.95 42.723 ;
		RECT	151.908 42.659 151.94 42.723 ;
		RECT	152.81 42.659 152.842 42.723 ;
		RECT	153.967 42.675 154.031 42.707 ;
		RECT	149.918 42.864 149.95 42.928 ;
		RECT	151.908 42.864 151.94 42.928 ;
		RECT	152.81 42.864 152.842 42.928 ;
		RECT	153.967 42.864 154.031 42.928 ;
		RECT	149.918 43.069 149.95 43.133 ;
		RECT	151.908 43.069 151.94 43.133 ;
		RECT	152.81 43.069 152.842 43.133 ;
		RECT	153.967 43.085 154.031 43.117 ;
		RECT	152.655 44.026 152.687 44.09 ;
		RECT	152.807 44.026 152.839 44.09 ;
		RECT	153.206 44.042 153.27 44.074 ;
		RECT	149.965 2.939 149.997 2.971 ;
		RECT	151.908 3.044 151.94 3.076 ;
		RECT	148.377 3.374 148.441 3.406 ;
		RECT	149.272 3.374 149.304 3.406 ;
		RECT	149.792 3.374 149.824 3.406 ;
		RECT	151.705 3.374 151.737 3.406 ;
		RECT	153.214 3.374 153.278 3.406 ;
		RECT	154.142 3.374 154.174 3.406 ;
		RECT	154.662 3.374 154.694 3.406 ;
		RECT	155.529 3.374 155.593 3.406 ;
		RECT	150.034 3.479 150.066 3.511 ;
		RECT	153.568 3.613 153.6 3.677 ;
		RECT	150.122 3.629 150.154 3.661 ;
		RECT	150.575 3.629 150.607 3.661 ;
		RECT	151.146 3.629 151.178 3.661 ;
		RECT	152.244 3.629 152.276 3.661 ;
		RECT	153.805 3.629 153.837 3.661 ;
		RECT	149.965 20.219 149.997 20.251 ;
		RECT	151.908 20.324 151.94 20.356 ;
		RECT	148.377 20.654 148.441 20.686 ;
		RECT	149.272 20.654 149.304 20.686 ;
		RECT	149.792 20.654 149.824 20.686 ;
		RECT	151.705 20.654 151.737 20.686 ;
		RECT	153.214 20.654 153.278 20.686 ;
		RECT	154.142 20.654 154.174 20.686 ;
		RECT	154.662 20.654 154.694 20.686 ;
		RECT	155.529 20.654 155.593 20.686 ;
		RECT	150.034 20.759 150.066 20.791 ;
		RECT	153.568 20.893 153.6 20.957 ;
		RECT	150.122 20.909 150.154 20.941 ;
		RECT	150.575 20.909 150.607 20.941 ;
		RECT	151.146 20.909 151.178 20.941 ;
		RECT	152.244 20.909 152.276 20.941 ;
		RECT	153.805 20.909 153.837 20.941 ;
		RECT	149.965 22.139 149.997 22.171 ;
		RECT	151.908 22.244 151.94 22.276 ;
		RECT	148.377 22.574 148.441 22.606 ;
		RECT	149.272 22.574 149.304 22.606 ;
		RECT	149.792 22.574 149.824 22.606 ;
		RECT	151.705 22.574 151.737 22.606 ;
		RECT	153.214 22.574 153.278 22.606 ;
		RECT	154.142 22.574 154.174 22.606 ;
		RECT	154.662 22.574 154.694 22.606 ;
		RECT	155.529 22.574 155.593 22.606 ;
		RECT	150.034 22.679 150.066 22.711 ;
		RECT	153.568 22.813 153.6 22.877 ;
		RECT	150.122 22.829 150.154 22.861 ;
		RECT	150.575 22.829 150.607 22.861 ;
		RECT	151.146 22.829 151.178 22.861 ;
		RECT	152.244 22.829 152.276 22.861 ;
		RECT	153.805 22.829 153.837 22.861 ;
		RECT	149.965 24.059 149.997 24.091 ;
		RECT	151.908 24.164 151.94 24.196 ;
		RECT	148.377 24.494 148.441 24.526 ;
		RECT	149.272 24.494 149.304 24.526 ;
		RECT	149.792 24.494 149.824 24.526 ;
		RECT	151.705 24.494 151.737 24.526 ;
		RECT	153.214 24.494 153.278 24.526 ;
		RECT	154.142 24.494 154.174 24.526 ;
		RECT	154.662 24.494 154.694 24.526 ;
		RECT	155.529 24.494 155.593 24.526 ;
		RECT	150.034 24.599 150.066 24.631 ;
		RECT	153.568 24.733 153.6 24.797 ;
		RECT	150.122 24.749 150.154 24.781 ;
		RECT	150.575 24.749 150.607 24.781 ;
		RECT	151.146 24.749 151.178 24.781 ;
		RECT	152.244 24.749 152.276 24.781 ;
		RECT	153.805 24.749 153.837 24.781 ;
		RECT	149.965 25.979 149.997 26.011 ;
		RECT	151.908 26.084 151.94 26.116 ;
		RECT	148.377 26.414 148.441 26.446 ;
		RECT	149.272 26.414 149.304 26.446 ;
		RECT	149.792 26.414 149.824 26.446 ;
		RECT	151.705 26.414 151.737 26.446 ;
		RECT	153.214 26.414 153.278 26.446 ;
		RECT	154.142 26.414 154.174 26.446 ;
		RECT	154.662 26.414 154.694 26.446 ;
		RECT	155.529 26.414 155.593 26.446 ;
		RECT	150.034 26.519 150.066 26.551 ;
		RECT	153.568 26.653 153.6 26.717 ;
		RECT	150.122 26.669 150.154 26.701 ;
		RECT	150.575 26.669 150.607 26.701 ;
		RECT	151.146 26.669 151.178 26.701 ;
		RECT	152.244 26.669 152.276 26.701 ;
		RECT	153.805 26.669 153.837 26.701 ;
		RECT	149.965 27.899 149.997 27.931 ;
		RECT	151.908 28.004 151.94 28.036 ;
		RECT	148.377 28.334 148.441 28.366 ;
		RECT	149.272 28.334 149.304 28.366 ;
		RECT	149.792 28.334 149.824 28.366 ;
		RECT	151.705 28.334 151.737 28.366 ;
		RECT	153.214 28.334 153.278 28.366 ;
		RECT	154.142 28.334 154.174 28.366 ;
		RECT	154.662 28.334 154.694 28.366 ;
		RECT	155.529 28.334 155.593 28.366 ;
		RECT	150.034 28.439 150.066 28.471 ;
		RECT	153.568 28.573 153.6 28.637 ;
		RECT	150.122 28.589 150.154 28.621 ;
		RECT	150.575 28.589 150.607 28.621 ;
		RECT	151.146 28.589 151.178 28.621 ;
		RECT	152.244 28.589 152.276 28.621 ;
		RECT	153.805 28.589 153.837 28.621 ;
		RECT	149.965 4.859 149.997 4.891 ;
		RECT	151.908 4.964 151.94 4.996 ;
		RECT	148.377 5.294 148.441 5.326 ;
		RECT	149.272 5.294 149.304 5.326 ;
		RECT	149.792 5.294 149.824 5.326 ;
		RECT	151.705 5.294 151.737 5.326 ;
		RECT	153.214 5.294 153.278 5.326 ;
		RECT	154.142 5.294 154.174 5.326 ;
		RECT	154.662 5.294 154.694 5.326 ;
		RECT	155.529 5.294 155.593 5.326 ;
		RECT	150.034 5.399 150.066 5.431 ;
		RECT	153.568 5.533 153.6 5.597 ;
		RECT	150.122 5.549 150.154 5.581 ;
		RECT	150.575 5.549 150.607 5.581 ;
		RECT	151.146 5.549 151.178 5.581 ;
		RECT	152.244 5.549 152.276 5.581 ;
		RECT	153.805 5.549 153.837 5.581 ;
		RECT	149.965 6.779 149.997 6.811 ;
		RECT	151.908 6.884 151.94 6.916 ;
		RECT	148.377 7.214 148.441 7.246 ;
		RECT	149.272 7.214 149.304 7.246 ;
		RECT	149.792 7.214 149.824 7.246 ;
		RECT	151.705 7.214 151.737 7.246 ;
		RECT	153.214 7.214 153.278 7.246 ;
		RECT	154.142 7.214 154.174 7.246 ;
		RECT	154.662 7.214 154.694 7.246 ;
		RECT	155.529 7.214 155.593 7.246 ;
		RECT	150.034 7.319 150.066 7.351 ;
		RECT	153.568 7.453 153.6 7.517 ;
		RECT	150.122 7.469 150.154 7.501 ;
		RECT	150.575 7.469 150.607 7.501 ;
		RECT	151.146 7.469 151.178 7.501 ;
		RECT	152.244 7.469 152.276 7.501 ;
		RECT	153.805 7.469 153.837 7.501 ;
		RECT	149.965 8.699 149.997 8.731 ;
		RECT	151.908 8.804 151.94 8.836 ;
		RECT	148.377 9.134 148.441 9.166 ;
		RECT	149.272 9.134 149.304 9.166 ;
		RECT	149.792 9.134 149.824 9.166 ;
		RECT	151.705 9.134 151.737 9.166 ;
		RECT	153.214 9.134 153.278 9.166 ;
		RECT	154.142 9.134 154.174 9.166 ;
		RECT	154.662 9.134 154.694 9.166 ;
		RECT	155.529 9.134 155.593 9.166 ;
		RECT	150.034 9.239 150.066 9.271 ;
		RECT	153.568 9.373 153.6 9.437 ;
		RECT	150.122 9.389 150.154 9.421 ;
		RECT	150.575 9.389 150.607 9.421 ;
		RECT	151.146 9.389 151.178 9.421 ;
		RECT	152.244 9.389 152.276 9.421 ;
		RECT	153.805 9.389 153.837 9.421 ;
		RECT	149.965 10.619 149.997 10.651 ;
		RECT	151.908 10.724 151.94 10.756 ;
		RECT	148.377 11.054 148.441 11.086 ;
		RECT	149.272 11.054 149.304 11.086 ;
		RECT	149.792 11.054 149.824 11.086 ;
		RECT	151.705 11.054 151.737 11.086 ;
		RECT	153.214 11.054 153.278 11.086 ;
		RECT	154.142 11.054 154.174 11.086 ;
		RECT	154.662 11.054 154.694 11.086 ;
		RECT	155.529 11.054 155.593 11.086 ;
		RECT	150.034 11.159 150.066 11.191 ;
		RECT	153.568 11.293 153.6 11.357 ;
		RECT	150.122 11.309 150.154 11.341 ;
		RECT	150.575 11.309 150.607 11.341 ;
		RECT	151.146 11.309 151.178 11.341 ;
		RECT	152.244 11.309 152.276 11.341 ;
		RECT	153.805 11.309 153.837 11.341 ;
		RECT	149.965 12.539 149.997 12.571 ;
		RECT	151.908 12.644 151.94 12.676 ;
		RECT	148.377 12.974 148.441 13.006 ;
		RECT	149.272 12.974 149.304 13.006 ;
		RECT	149.792 12.974 149.824 13.006 ;
		RECT	151.705 12.974 151.737 13.006 ;
		RECT	153.214 12.974 153.278 13.006 ;
		RECT	154.142 12.974 154.174 13.006 ;
		RECT	154.662 12.974 154.694 13.006 ;
		RECT	155.529 12.974 155.593 13.006 ;
		RECT	150.034 13.079 150.066 13.111 ;
		RECT	153.568 13.213 153.6 13.277 ;
		RECT	150.122 13.229 150.154 13.261 ;
		RECT	150.575 13.229 150.607 13.261 ;
		RECT	151.146 13.229 151.178 13.261 ;
		RECT	152.244 13.229 152.276 13.261 ;
		RECT	153.805 13.229 153.837 13.261 ;
		RECT	149.965 14.459 149.997 14.491 ;
		RECT	151.908 14.564 151.94 14.596 ;
		RECT	148.377 14.894 148.441 14.926 ;
		RECT	149.272 14.894 149.304 14.926 ;
		RECT	149.792 14.894 149.824 14.926 ;
		RECT	151.705 14.894 151.737 14.926 ;
		RECT	153.214 14.894 153.278 14.926 ;
		RECT	154.142 14.894 154.174 14.926 ;
		RECT	154.662 14.894 154.694 14.926 ;
		RECT	155.529 14.894 155.593 14.926 ;
		RECT	150.034 14.999 150.066 15.031 ;
		RECT	153.568 15.133 153.6 15.197 ;
		RECT	150.122 15.149 150.154 15.181 ;
		RECT	150.575 15.149 150.607 15.181 ;
		RECT	151.146 15.149 151.178 15.181 ;
		RECT	152.244 15.149 152.276 15.181 ;
		RECT	153.805 15.149 153.837 15.181 ;
		RECT	149.965 16.379 149.997 16.411 ;
		RECT	151.908 16.484 151.94 16.516 ;
		RECT	148.377 16.814 148.441 16.846 ;
		RECT	149.272 16.814 149.304 16.846 ;
		RECT	149.792 16.814 149.824 16.846 ;
		RECT	151.705 16.814 151.737 16.846 ;
		RECT	153.214 16.814 153.278 16.846 ;
		RECT	154.142 16.814 154.174 16.846 ;
		RECT	154.662 16.814 154.694 16.846 ;
		RECT	155.529 16.814 155.593 16.846 ;
		RECT	150.034 16.919 150.066 16.951 ;
		RECT	153.568 17.053 153.6 17.117 ;
		RECT	150.122 17.069 150.154 17.101 ;
		RECT	150.575 17.069 150.607 17.101 ;
		RECT	151.146 17.069 151.178 17.101 ;
		RECT	152.244 17.069 152.276 17.101 ;
		RECT	153.805 17.069 153.837 17.101 ;
		RECT	149.965 18.299 149.997 18.331 ;
		RECT	151.908 18.404 151.94 18.436 ;
		RECT	148.377 18.734 148.441 18.766 ;
		RECT	149.272 18.734 149.304 18.766 ;
		RECT	149.792 18.734 149.824 18.766 ;
		RECT	151.705 18.734 151.737 18.766 ;
		RECT	153.214 18.734 153.278 18.766 ;
		RECT	154.142 18.734 154.174 18.766 ;
		RECT	154.662 18.734 154.694 18.766 ;
		RECT	155.529 18.734 155.593 18.766 ;
		RECT	150.034 18.839 150.066 18.871 ;
		RECT	153.568 18.973 153.6 19.037 ;
		RECT	150.122 18.989 150.154 19.021 ;
		RECT	150.575 18.989 150.607 19.021 ;
		RECT	151.146 18.989 151.178 19.021 ;
		RECT	152.244 18.989 152.276 19.021 ;
		RECT	153.805 18.989 153.837 19.021 ;
		RECT	149.965 1.019 149.997 1.051 ;
		RECT	151.908 1.124 151.94 1.156 ;
		RECT	148.377 1.454 148.441 1.486 ;
		RECT	149.272 1.454 149.304 1.486 ;
		RECT	149.792 1.454 149.824 1.486 ;
		RECT	151.705 1.454 151.737 1.486 ;
		RECT	153.214 1.454 153.278 1.486 ;
		RECT	154.142 1.454 154.174 1.486 ;
		RECT	154.662 1.454 154.694 1.486 ;
		RECT	155.529 1.454 155.593 1.486 ;
		RECT	150.034 1.559 150.066 1.591 ;
		RECT	153.568 1.693 153.6 1.757 ;
		RECT	150.122 1.709 150.154 1.741 ;
		RECT	150.575 1.709 150.607 1.741 ;
		RECT	151.146 1.709 151.178 1.741 ;
		RECT	152.244 1.709 152.276 1.741 ;
		RECT	153.805 1.709 153.837 1.741 ;
		RECT	149.965 29.819 149.997 29.851 ;
		RECT	151.908 29.924 151.94 29.956 ;
		RECT	148.377 30.254 148.441 30.286 ;
		RECT	149.272 30.254 149.304 30.286 ;
		RECT	149.792 30.254 149.824 30.286 ;
		RECT	151.705 30.254 151.737 30.286 ;
		RECT	153.214 30.254 153.278 30.286 ;
		RECT	154.142 30.254 154.174 30.286 ;
		RECT	154.662 30.254 154.694 30.286 ;
		RECT	155.529 30.254 155.593 30.286 ;
		RECT	150.034 30.359 150.066 30.391 ;
		RECT	153.568 30.493 153.6 30.557 ;
		RECT	150.122 30.509 150.154 30.541 ;
		RECT	150.575 30.509 150.607 30.541 ;
		RECT	151.146 30.509 151.178 30.541 ;
		RECT	152.244 30.509 152.276 30.541 ;
		RECT	153.805 30.509 153.837 30.541 ;
		RECT	150.457 1.964 150.489 1.996 ;
		RECT	150.457 3.884 150.489 3.916 ;
		RECT	150.457 5.804 150.489 5.836 ;
		RECT	150.457 7.724 150.489 7.756 ;
		RECT	150.457 9.644 150.489 9.676 ;
		RECT	150.457 11.564 150.489 11.596 ;
		RECT	150.457 13.484 150.489 13.516 ;
		RECT	150.457 15.404 150.489 15.436 ;
		RECT	150.457 17.324 150.489 17.356 ;
		RECT	150.457 19.244 150.489 19.276 ;
		RECT	150.457 21.164 150.489 21.196 ;
		RECT	150.457 23.084 150.489 23.116 ;
		RECT	150.457 25.004 150.489 25.036 ;
		RECT	150.457 26.924 150.489 26.956 ;
		RECT	150.457 28.844 150.489 28.876 ;
		RECT	150.457 30.764 150.489 30.796 ;
		RECT	151.908 1.693 151.94 1.757 ;
		RECT	151.908 20.893 151.94 20.957 ;
		RECT	151.908 22.813 151.94 22.877 ;
		RECT	151.908 24.733 151.94 24.797 ;
		RECT	151.908 26.653 151.94 26.717 ;
		RECT	151.908 28.573 151.94 28.637 ;
		RECT	151.908 30.493 151.94 30.557 ;
		RECT	151.908 3.613 151.94 3.677 ;
		RECT	151.908 5.533 151.94 5.597 ;
		RECT	151.908 7.453 151.94 7.517 ;
		RECT	151.908 9.373 151.94 9.437 ;
		RECT	151.908 11.293 151.94 11.357 ;
		RECT	151.908 13.213 151.94 13.277 ;
		RECT	151.908 15.133 151.94 15.197 ;
		RECT	151.908 17.053 151.94 17.117 ;
		RECT	151.908 18.973 151.94 19.037 ;
		RECT	149.965 54.245 149.997 54.277 ;
		RECT	151.908 54.14 151.94 54.172 ;
		RECT	148.377 53.81 148.441 53.842 ;
		RECT	149.272 53.81 149.304 53.842 ;
		RECT	149.792 53.81 149.824 53.842 ;
		RECT	151.705 53.81 151.737 53.842 ;
		RECT	153.214 53.81 153.278 53.842 ;
		RECT	154.142 53.81 154.174 53.842 ;
		RECT	154.662 53.81 154.694 53.842 ;
		RECT	155.529 53.81 155.593 53.842 ;
		RECT	150.034 53.705 150.066 53.737 ;
		RECT	153.568 53.539 153.6 53.603 ;
		RECT	150.122 53.555 150.154 53.587 ;
		RECT	150.575 53.555 150.607 53.587 ;
		RECT	151.146 53.555 151.178 53.587 ;
		RECT	152.244 53.555 152.276 53.587 ;
		RECT	153.805 53.555 153.837 53.587 ;
		RECT	149.965 71.525 149.997 71.557 ;
		RECT	151.908 71.42 151.94 71.452 ;
		RECT	148.377 71.09 148.441 71.122 ;
		RECT	149.272 71.09 149.304 71.122 ;
		RECT	149.792 71.09 149.824 71.122 ;
		RECT	151.705 71.09 151.737 71.122 ;
		RECT	153.214 71.09 153.278 71.122 ;
		RECT	154.142 71.09 154.174 71.122 ;
		RECT	154.662 71.09 154.694 71.122 ;
		RECT	155.529 71.09 155.593 71.122 ;
		RECT	150.034 70.985 150.066 71.017 ;
		RECT	153.568 70.819 153.6 70.883 ;
		RECT	150.122 70.835 150.154 70.867 ;
		RECT	150.575 70.835 150.607 70.867 ;
		RECT	151.146 70.835 151.178 70.867 ;
		RECT	152.244 70.835 152.276 70.867 ;
		RECT	153.805 70.835 153.837 70.867 ;
		RECT	149.965 73.445 149.997 73.477 ;
		RECT	151.908 73.34 151.94 73.372 ;
		RECT	148.377 73.01 148.441 73.042 ;
		RECT	149.272 73.01 149.304 73.042 ;
		RECT	149.792 73.01 149.824 73.042 ;
		RECT	151.705 73.01 151.737 73.042 ;
		RECT	153.214 73.01 153.278 73.042 ;
		RECT	154.142 73.01 154.174 73.042 ;
		RECT	154.662 73.01 154.694 73.042 ;
		RECT	155.529 73.01 155.593 73.042 ;
		RECT	150.034 72.905 150.066 72.937 ;
		RECT	153.568 72.739 153.6 72.803 ;
		RECT	150.122 72.755 150.154 72.787 ;
		RECT	150.575 72.755 150.607 72.787 ;
		RECT	151.146 72.755 151.178 72.787 ;
		RECT	152.244 72.755 152.276 72.787 ;
		RECT	153.805 72.755 153.837 72.787 ;
		RECT	149.965 75.365 149.997 75.397 ;
		RECT	151.908 75.26 151.94 75.292 ;
		RECT	148.377 74.93 148.441 74.962 ;
		RECT	149.272 74.93 149.304 74.962 ;
		RECT	149.792 74.93 149.824 74.962 ;
		RECT	151.705 74.93 151.737 74.962 ;
		RECT	153.214 74.93 153.278 74.962 ;
		RECT	154.142 74.93 154.174 74.962 ;
		RECT	154.662 74.93 154.694 74.962 ;
		RECT	155.529 74.93 155.593 74.962 ;
		RECT	150.034 74.825 150.066 74.857 ;
		RECT	153.568 74.659 153.6 74.723 ;
		RECT	150.122 74.675 150.154 74.707 ;
		RECT	150.575 74.675 150.607 74.707 ;
		RECT	151.146 74.675 151.178 74.707 ;
		RECT	152.244 74.675 152.276 74.707 ;
		RECT	153.805 74.675 153.837 74.707 ;
		RECT	149.965 77.285 149.997 77.317 ;
		RECT	151.908 77.18 151.94 77.212 ;
		RECT	148.377 76.85 148.441 76.882 ;
		RECT	149.272 76.85 149.304 76.882 ;
		RECT	149.792 76.85 149.824 76.882 ;
		RECT	151.705 76.85 151.737 76.882 ;
		RECT	153.214 76.85 153.278 76.882 ;
		RECT	154.142 76.85 154.174 76.882 ;
		RECT	154.662 76.85 154.694 76.882 ;
		RECT	155.529 76.85 155.593 76.882 ;
		RECT	150.034 76.745 150.066 76.777 ;
		RECT	153.568 76.579 153.6 76.643 ;
		RECT	150.122 76.595 150.154 76.627 ;
		RECT	150.575 76.595 150.607 76.627 ;
		RECT	151.146 76.595 151.178 76.627 ;
		RECT	152.244 76.595 152.276 76.627 ;
		RECT	153.805 76.595 153.837 76.627 ;
		RECT	149.965 79.205 149.997 79.237 ;
		RECT	151.908 79.1 151.94 79.132 ;
		RECT	148.377 78.77 148.441 78.802 ;
		RECT	149.272 78.77 149.304 78.802 ;
		RECT	149.792 78.77 149.824 78.802 ;
		RECT	151.705 78.77 151.737 78.802 ;
		RECT	153.214 78.77 153.278 78.802 ;
		RECT	154.142 78.77 154.174 78.802 ;
		RECT	154.662 78.77 154.694 78.802 ;
		RECT	155.529 78.77 155.593 78.802 ;
		RECT	150.034 78.665 150.066 78.697 ;
		RECT	153.568 78.499 153.6 78.563 ;
		RECT	150.122 78.515 150.154 78.547 ;
		RECT	150.575 78.515 150.607 78.547 ;
		RECT	151.146 78.515 151.178 78.547 ;
		RECT	152.244 78.515 152.276 78.547 ;
		RECT	153.805 78.515 153.837 78.547 ;
		RECT	149.965 56.165 149.997 56.197 ;
		RECT	151.908 56.06 151.94 56.092 ;
		RECT	148.377 55.73 148.441 55.762 ;
		RECT	149.272 55.73 149.304 55.762 ;
		RECT	149.792 55.73 149.824 55.762 ;
		RECT	151.705 55.73 151.737 55.762 ;
		RECT	153.214 55.73 153.278 55.762 ;
		RECT	154.142 55.73 154.174 55.762 ;
		RECT	154.662 55.73 154.694 55.762 ;
		RECT	155.529 55.73 155.593 55.762 ;
		RECT	150.034 55.625 150.066 55.657 ;
		RECT	153.568 55.459 153.6 55.523 ;
		RECT	150.122 55.475 150.154 55.507 ;
		RECT	150.575 55.475 150.607 55.507 ;
		RECT	151.146 55.475 151.178 55.507 ;
		RECT	152.244 55.475 152.276 55.507 ;
		RECT	153.805 55.475 153.837 55.507 ;
		RECT	149.965 58.085 149.997 58.117 ;
		RECT	151.908 57.98 151.94 58.012 ;
		RECT	148.377 57.65 148.441 57.682 ;
		RECT	149.272 57.65 149.304 57.682 ;
		RECT	149.792 57.65 149.824 57.682 ;
		RECT	151.705 57.65 151.737 57.682 ;
		RECT	153.214 57.65 153.278 57.682 ;
		RECT	154.142 57.65 154.174 57.682 ;
		RECT	154.662 57.65 154.694 57.682 ;
		RECT	155.529 57.65 155.593 57.682 ;
		RECT	150.034 57.545 150.066 57.577 ;
		RECT	153.568 57.379 153.6 57.443 ;
		RECT	150.122 57.395 150.154 57.427 ;
		RECT	150.575 57.395 150.607 57.427 ;
		RECT	151.146 57.395 151.178 57.427 ;
		RECT	152.244 57.395 152.276 57.427 ;
		RECT	153.805 57.395 153.837 57.427 ;
		RECT	149.965 60.005 149.997 60.037 ;
		RECT	151.908 59.9 151.94 59.932 ;
		RECT	148.377 59.57 148.441 59.602 ;
		RECT	149.272 59.57 149.304 59.602 ;
		RECT	149.792 59.57 149.824 59.602 ;
		RECT	151.705 59.57 151.737 59.602 ;
		RECT	153.214 59.57 153.278 59.602 ;
		RECT	154.142 59.57 154.174 59.602 ;
		RECT	154.662 59.57 154.694 59.602 ;
		RECT	155.529 59.57 155.593 59.602 ;
		RECT	150.034 59.465 150.066 59.497 ;
		RECT	153.568 59.299 153.6 59.363 ;
		RECT	150.122 59.315 150.154 59.347 ;
		RECT	150.575 59.315 150.607 59.347 ;
		RECT	151.146 59.315 151.178 59.347 ;
		RECT	152.244 59.315 152.276 59.347 ;
		RECT	153.805 59.315 153.837 59.347 ;
		RECT	149.965 61.925 149.997 61.957 ;
		RECT	151.908 61.82 151.94 61.852 ;
		RECT	148.377 61.49 148.441 61.522 ;
		RECT	149.272 61.49 149.304 61.522 ;
		RECT	149.792 61.49 149.824 61.522 ;
		RECT	151.705 61.49 151.737 61.522 ;
		RECT	153.214 61.49 153.278 61.522 ;
		RECT	154.142 61.49 154.174 61.522 ;
		RECT	154.662 61.49 154.694 61.522 ;
		RECT	155.529 61.49 155.593 61.522 ;
		RECT	150.034 61.385 150.066 61.417 ;
		RECT	153.568 61.219 153.6 61.283 ;
		RECT	150.122 61.235 150.154 61.267 ;
		RECT	150.575 61.235 150.607 61.267 ;
		RECT	151.146 61.235 151.178 61.267 ;
		RECT	152.244 61.235 152.276 61.267 ;
		RECT	153.805 61.235 153.837 61.267 ;
		RECT	149.965 63.845 149.997 63.877 ;
		RECT	151.908 63.74 151.94 63.772 ;
		RECT	148.377 63.41 148.441 63.442 ;
		RECT	149.272 63.41 149.304 63.442 ;
		RECT	149.792 63.41 149.824 63.442 ;
		RECT	151.705 63.41 151.737 63.442 ;
		RECT	153.214 63.41 153.278 63.442 ;
		RECT	154.142 63.41 154.174 63.442 ;
		RECT	154.662 63.41 154.694 63.442 ;
		RECT	155.529 63.41 155.593 63.442 ;
		RECT	150.034 63.305 150.066 63.337 ;
		RECT	153.568 63.139 153.6 63.203 ;
		RECT	150.122 63.155 150.154 63.187 ;
		RECT	150.575 63.155 150.607 63.187 ;
		RECT	151.146 63.155 151.178 63.187 ;
		RECT	152.244 63.155 152.276 63.187 ;
		RECT	153.805 63.155 153.837 63.187 ;
		RECT	149.965 65.765 149.997 65.797 ;
		RECT	151.908 65.66 151.94 65.692 ;
		RECT	148.377 65.33 148.441 65.362 ;
		RECT	149.272 65.33 149.304 65.362 ;
		RECT	149.792 65.33 149.824 65.362 ;
		RECT	151.705 65.33 151.737 65.362 ;
		RECT	153.214 65.33 153.278 65.362 ;
		RECT	154.142 65.33 154.174 65.362 ;
		RECT	154.662 65.33 154.694 65.362 ;
		RECT	155.529 65.33 155.593 65.362 ;
		RECT	150.034 65.225 150.066 65.257 ;
		RECT	153.568 65.059 153.6 65.123 ;
		RECT	150.122 65.075 150.154 65.107 ;
		RECT	150.575 65.075 150.607 65.107 ;
		RECT	151.146 65.075 151.178 65.107 ;
		RECT	152.244 65.075 152.276 65.107 ;
		RECT	153.805 65.075 153.837 65.107 ;
		RECT	149.965 67.685 149.997 67.717 ;
		RECT	151.908 67.58 151.94 67.612 ;
		RECT	148.377 67.25 148.441 67.282 ;
		RECT	149.272 67.25 149.304 67.282 ;
		RECT	149.792 67.25 149.824 67.282 ;
		RECT	151.705 67.25 151.737 67.282 ;
		RECT	153.214 67.25 153.278 67.282 ;
		RECT	154.142 67.25 154.174 67.282 ;
		RECT	154.662 67.25 154.694 67.282 ;
		RECT	155.529 67.25 155.593 67.282 ;
		RECT	150.034 67.145 150.066 67.177 ;
		RECT	153.568 66.979 153.6 67.043 ;
		RECT	150.122 66.995 150.154 67.027 ;
		RECT	150.575 66.995 150.607 67.027 ;
		RECT	151.146 66.995 151.178 67.027 ;
		RECT	152.244 66.995 152.276 67.027 ;
		RECT	153.805 66.995 153.837 67.027 ;
		RECT	149.965 69.605 149.997 69.637 ;
		RECT	151.908 69.5 151.94 69.532 ;
		RECT	148.377 69.17 148.441 69.202 ;
		RECT	149.272 69.17 149.304 69.202 ;
		RECT	149.792 69.17 149.824 69.202 ;
		RECT	151.705 69.17 151.737 69.202 ;
		RECT	153.214 69.17 153.278 69.202 ;
		RECT	154.142 69.17 154.174 69.202 ;
		RECT	154.662 69.17 154.694 69.202 ;
		RECT	155.529 69.17 155.593 69.202 ;
		RECT	150.034 69.065 150.066 69.097 ;
		RECT	153.568 68.899 153.6 68.963 ;
		RECT	150.122 68.915 150.154 68.947 ;
		RECT	150.575 68.915 150.607 68.947 ;
		RECT	151.146 68.915 151.178 68.947 ;
		RECT	152.244 68.915 152.276 68.947 ;
		RECT	153.805 68.915 153.837 68.947 ;
		RECT	149.965 52.325 149.997 52.357 ;
		RECT	151.908 52.22 151.94 52.252 ;
		RECT	148.377 51.89 148.441 51.922 ;
		RECT	149.272 51.89 149.304 51.922 ;
		RECT	149.792 51.89 149.824 51.922 ;
		RECT	151.705 51.89 151.737 51.922 ;
		RECT	153.214 51.89 153.278 51.922 ;
		RECT	154.142 51.89 154.174 51.922 ;
		RECT	154.662 51.89 154.694 51.922 ;
		RECT	155.529 51.89 155.593 51.922 ;
		RECT	150.034 51.785 150.066 51.817 ;
		RECT	153.568 51.619 153.6 51.683 ;
		RECT	150.122 51.635 150.154 51.667 ;
		RECT	150.575 51.635 150.607 51.667 ;
		RECT	151.146 51.635 151.178 51.667 ;
		RECT	152.244 51.635 152.276 51.667 ;
		RECT	153.805 51.635 153.837 51.667 ;
		RECT	149.965 81.125 149.997 81.157 ;
		RECT	151.908 81.02 151.94 81.052 ;
		RECT	148.377 80.69 148.441 80.722 ;
		RECT	149.272 80.69 149.304 80.722 ;
		RECT	149.792 80.69 149.824 80.722 ;
		RECT	151.705 80.69 151.737 80.722 ;
		RECT	153.214 80.69 153.278 80.722 ;
		RECT	154.142 80.69 154.174 80.722 ;
		RECT	154.662 80.69 154.694 80.722 ;
		RECT	155.529 80.69 155.593 80.722 ;
		RECT	150.034 80.585 150.066 80.617 ;
		RECT	153.568 80.419 153.6 80.483 ;
		RECT	150.122 80.435 150.154 80.467 ;
		RECT	150.575 80.435 150.607 80.467 ;
		RECT	151.146 80.435 151.178 80.467 ;
		RECT	152.244 80.435 152.276 80.467 ;
		RECT	153.805 80.435 153.837 80.467 ;
		RECT	150.457 51.38 150.489 51.412 ;
		RECT	150.457 53.3 150.489 53.332 ;
		RECT	150.457 55.22 150.489 55.252 ;
		RECT	150.457 57.14 150.489 57.172 ;
		RECT	150.457 59.06 150.489 59.092 ;
		RECT	150.457 60.98 150.489 61.012 ;
		RECT	150.457 62.9 150.489 62.932 ;
		RECT	150.457 64.82 150.489 64.852 ;
		RECT	150.457 66.74 150.489 66.772 ;
		RECT	150.457 68.66 150.489 68.692 ;
		RECT	150.457 70.58 150.489 70.612 ;
		RECT	150.457 72.5 150.489 72.532 ;
		RECT	150.457 74.42 150.489 74.452 ;
		RECT	150.457 76.34 150.489 76.372 ;
		RECT	150.457 78.26 150.489 78.292 ;
		RECT	150.457 80.18 150.489 80.212 ;
		RECT	151.908 51.619 151.94 51.683 ;
		RECT	151.908 70.819 151.94 70.883 ;
		RECT	151.908 72.739 151.94 72.803 ;
		RECT	151.908 74.659 151.94 74.723 ;
		RECT	151.908 76.579 151.94 76.643 ;
		RECT	151.908 78.499 151.94 78.563 ;
		RECT	151.908 80.419 151.94 80.483 ;
		RECT	151.908 53.539 151.94 53.603 ;
		RECT	151.908 55.459 151.94 55.523 ;
		RECT	151.908 57.379 151.94 57.443 ;
		RECT	151.908 59.299 151.94 59.363 ;
		RECT	151.908 61.219 151.94 61.283 ;
		RECT	151.908 63.139 151.94 63.203 ;
		RECT	151.908 65.059 151.94 65.123 ;
		RECT	151.908 66.979 151.94 67.043 ;
		RECT	151.908 68.899 151.94 68.963 ;
		RECT	103.512 31.762 103.576 31.794 ;
		RECT	103.512 50.382 103.576 50.414 ;
		RECT	125.555 39.858 125.587 39.89 ;
		RECT	122.195 39.358 122.227 39.39 ;
		RECT	121.859 39.358 121.891 39.39 ;
		RECT	121.523 39.258 121.555 39.29 ;
		RECT	121.187 39.258 121.219 39.29 ;
		RECT	120.851 39.158 120.883 39.19 ;
		RECT	120.515 39.158 120.547 39.19 ;
		RECT	120.179 39.858 120.211 39.89 ;
		RECT	119.843 39.858 119.875 39.89 ;
		RECT	119.507 39.758 119.539 39.79 ;
		RECT	119.171 39.758 119.203 39.79 ;
		RECT	125.219 39.858 125.251 39.89 ;
		RECT	118.835 39.658 118.867 39.69 ;
		RECT	118.499 39.658 118.531 39.69 ;
		RECT	118.163 39.558 118.195 39.59 ;
		RECT	117.827 39.558 117.859 39.59 ;
		RECT	117.491 39.458 117.523 39.49 ;
		RECT	117.155 39.458 117.187 39.49 ;
		RECT	116.819 39.358 116.851 39.39 ;
		RECT	116.483 39.358 116.515 39.39 ;
		RECT	116.147 39.258 116.179 39.29 ;
		RECT	115.811 39.258 115.843 39.29 ;
		RECT	124.883 39.758 124.915 39.79 ;
		RECT	115.475 39.158 115.507 39.19 ;
		RECT	115.139 39.158 115.171 39.19 ;
		RECT	114.803 39.858 114.835 39.89 ;
		RECT	114.467 39.858 114.499 39.89 ;
		RECT	114.131 39.758 114.163 39.79 ;
		RECT	113.795 39.758 113.827 39.79 ;
		RECT	113.459 39.658 113.491 39.69 ;
		RECT	113.123 39.658 113.155 39.69 ;
		RECT	112.787 39.558 112.819 39.59 ;
		RECT	112.451 39.558 112.483 39.59 ;
		RECT	124.547 39.758 124.579 39.79 ;
		RECT	112.115 39.458 112.147 39.49 ;
		RECT	111.779 39.458 111.811 39.49 ;
		RECT	111.443 39.358 111.475 39.39 ;
		RECT	111.107 39.358 111.139 39.39 ;
		RECT	110.771 39.258 110.803 39.29 ;
		RECT	110.435 39.258 110.467 39.29 ;
		RECT	110.099 39.158 110.131 39.19 ;
		RECT	109.763 39.158 109.795 39.19 ;
		RECT	109.427 39.858 109.459 39.89 ;
		RECT	109.091 39.858 109.123 39.89 ;
		RECT	124.211 39.658 124.243 39.69 ;
		RECT	108.755 39.758 108.787 39.79 ;
		RECT	108.419 39.758 108.451 39.79 ;
		RECT	108.083 39.658 108.115 39.69 ;
		RECT	107.747 39.658 107.779 39.69 ;
		RECT	107.411 39.558 107.443 39.59 ;
		RECT	107.075 39.558 107.107 39.59 ;
		RECT	106.739 39.458 106.771 39.49 ;
		RECT	106.403 39.458 106.435 39.49 ;
		RECT	106.067 39.358 106.099 39.39 ;
		RECT	105.731 39.358 105.763 39.39 ;
		RECT	123.875 39.658 123.907 39.69 ;
		RECT	105.395 39.258 105.427 39.29 ;
		RECT	105.059 39.258 105.091 39.29 ;
		RECT	104.723 39.158 104.755 39.19 ;
		RECT	104.387 39.158 104.419 39.19 ;
		RECT	123.539 39.558 123.571 39.59 ;
		RECT	123.203 39.558 123.235 39.59 ;
		RECT	122.867 39.458 122.899 39.49 ;
		RECT	122.531 39.458 122.563 39.49 ;
		RECT	125.555 42.825 125.587 42.857 ;
		RECT	122.195 42.825 122.227 42.857 ;
		RECT	121.859 42.825 121.891 42.857 ;
		RECT	121.523 42.825 121.555 42.857 ;
		RECT	121.187 42.825 121.219 42.857 ;
		RECT	120.851 42.825 120.883 42.857 ;
		RECT	120.515 42.825 120.547 42.857 ;
		RECT	120.179 42.925 120.211 42.957 ;
		RECT	119.843 42.925 119.875 42.957 ;
		RECT	119.507 42.925 119.539 42.957 ;
		RECT	119.171 42.925 119.203 42.957 ;
		RECT	125.219 42.825 125.251 42.857 ;
		RECT	118.835 42.925 118.867 42.957 ;
		RECT	118.499 42.925 118.531 42.957 ;
		RECT	118.163 42.925 118.195 42.957 ;
		RECT	117.827 42.925 117.859 42.957 ;
		RECT	117.491 42.925 117.523 42.957 ;
		RECT	117.155 42.925 117.187 42.957 ;
		RECT	116.819 42.925 116.851 42.957 ;
		RECT	116.483 42.925 116.515 42.957 ;
		RECT	116.147 42.925 116.179 42.957 ;
		RECT	115.811 42.925 115.843 42.957 ;
		RECT	124.883 42.825 124.915 42.857 ;
		RECT	115.475 42.925 115.507 42.957 ;
		RECT	115.139 42.925 115.171 42.957 ;
		RECT	114.803 43.025 114.835 43.057 ;
		RECT	114.467 43.025 114.499 43.057 ;
		RECT	114.131 43.025 114.163 43.057 ;
		RECT	113.795 43.025 113.827 43.057 ;
		RECT	113.459 43.025 113.491 43.057 ;
		RECT	113.123 43.025 113.155 43.057 ;
		RECT	112.787 43.025 112.819 43.057 ;
		RECT	112.451 43.025 112.483 43.057 ;
		RECT	124.547 42.825 124.579 42.857 ;
		RECT	112.115 43.025 112.147 43.057 ;
		RECT	111.779 43.025 111.811 43.057 ;
		RECT	111.443 43.025 111.475 43.057 ;
		RECT	111.107 43.025 111.139 43.057 ;
		RECT	110.771 43.025 110.803 43.057 ;
		RECT	110.435 43.025 110.467 43.057 ;
		RECT	110.099 43.025 110.131 43.057 ;
		RECT	109.763 43.025 109.795 43.057 ;
		RECT	109.427 43.125 109.459 43.157 ;
		RECT	109.091 43.125 109.123 43.157 ;
		RECT	124.211 42.825 124.243 42.857 ;
		RECT	108.755 43.125 108.787 43.157 ;
		RECT	108.419 43.125 108.451 43.157 ;
		RECT	108.083 43.125 108.115 43.157 ;
		RECT	107.747 43.125 107.779 43.157 ;
		RECT	107.411 43.125 107.443 43.157 ;
		RECT	107.075 43.125 107.107 43.157 ;
		RECT	106.739 43.125 106.771 43.157 ;
		RECT	106.403 43.125 106.435 43.157 ;
		RECT	106.067 43.125 106.099 43.157 ;
		RECT	105.731 43.125 105.763 43.157 ;
		RECT	123.875 42.825 123.907 42.857 ;
		RECT	105.395 43.125 105.427 43.157 ;
		RECT	105.059 43.125 105.091 43.157 ;
		RECT	104.723 43.125 104.755 43.157 ;
		RECT	104.387 43.125 104.419 43.157 ;
		RECT	123.539 42.825 123.571 42.857 ;
		RECT	123.203 42.825 123.235 42.857 ;
		RECT	122.867 42.825 122.899 42.857 ;
		RECT	122.531 42.825 122.563 42.857 ;
		RECT	125.513 32.691 125.545 32.755 ;
		RECT	147.709 39.672 147.741 39.736 ;
		RECT	147.673 44.026 147.705 44.09 ;
		RECT	122.153 32.691 122.185 32.755 ;
		RECT	121.817 32.691 121.849 32.755 ;
		RECT	121.481 32.691 121.513 32.755 ;
		RECT	121.145 32.691 121.177 32.755 ;
		RECT	120.809 32.691 120.841 32.755 ;
		RECT	120.473 32.691 120.505 32.755 ;
		RECT	120.137 32.691 120.169 32.755 ;
		RECT	119.801 32.691 119.833 32.755 ;
		RECT	119.465 32.691 119.497 32.755 ;
		RECT	119.129 32.691 119.161 32.755 ;
		RECT	125.177 32.691 125.209 32.755 ;
		RECT	118.793 32.691 118.825 32.755 ;
		RECT	118.457 32.691 118.489 32.755 ;
		RECT	118.121 32.691 118.153 32.755 ;
		RECT	117.785 32.691 117.817 32.755 ;
		RECT	117.449 32.691 117.481 32.755 ;
		RECT	117.113 32.691 117.145 32.755 ;
		RECT	116.777 32.691 116.809 32.755 ;
		RECT	116.441 32.691 116.473 32.755 ;
		RECT	116.105 32.691 116.137 32.755 ;
		RECT	115.769 32.691 115.801 32.755 ;
		RECT	124.841 32.691 124.873 32.755 ;
		RECT	115.433 32.691 115.465 32.755 ;
		RECT	115.097 32.691 115.129 32.755 ;
		RECT	114.761 32.691 114.793 32.755 ;
		RECT	114.425 32.691 114.457 32.755 ;
		RECT	114.089 32.691 114.121 32.755 ;
		RECT	113.753 32.691 113.785 32.755 ;
		RECT	113.417 32.691 113.449 32.755 ;
		RECT	113.081 32.691 113.113 32.755 ;
		RECT	112.745 32.691 112.777 32.755 ;
		RECT	112.409 32.691 112.441 32.755 ;
		RECT	124.505 32.691 124.537 32.755 ;
		RECT	112.073 32.691 112.105 32.755 ;
		RECT	111.737 32.691 111.769 32.755 ;
		RECT	111.401 32.691 111.433 32.755 ;
		RECT	111.065 32.691 111.097 32.755 ;
		RECT	110.729 32.691 110.761 32.755 ;
		RECT	110.393 32.691 110.425 32.755 ;
		RECT	110.057 32.691 110.089 32.755 ;
		RECT	109.721 32.691 109.753 32.755 ;
		RECT	109.385 32.691 109.417 32.755 ;
		RECT	109.049 32.691 109.081 32.755 ;
		RECT	124.169 32.691 124.201 32.755 ;
		RECT	108.713 32.691 108.745 32.755 ;
		RECT	108.377 32.691 108.409 32.755 ;
		RECT	108.041 32.691 108.073 32.755 ;
		RECT	107.705 32.691 107.737 32.755 ;
		RECT	107.369 32.691 107.401 32.755 ;
		RECT	107.033 32.691 107.065 32.755 ;
		RECT	106.697 32.691 106.729 32.755 ;
		RECT	106.361 32.691 106.393 32.755 ;
		RECT	106.025 32.691 106.057 32.755 ;
		RECT	105.689 32.691 105.721 32.755 ;
		RECT	123.833 32.691 123.865 32.755 ;
		RECT	105.353 32.691 105.385 32.755 ;
		RECT	105.017 32.691 105.049 32.755 ;
		RECT	104.681 32.691 104.713 32.755 ;
		RECT	104.345 32.691 104.377 32.755 ;
		RECT	123.497 32.691 123.529 32.755 ;
		RECT	123.161 32.691 123.193 32.755 ;
		RECT	122.825 32.691 122.857 32.755 ;
		RECT	122.489 32.691 122.521 32.755 ;
		RECT	141.678 43.125 141.71 43.157 ;
		RECT	140.67 43.125 140.702 43.157 ;
		RECT	139.326 43.125 139.358 43.157 ;
		RECT	138.318 43.125 138.35 43.157 ;
		RECT	136.638 43.125 136.67 43.157 ;
		RECT	136.302 43.125 136.334 43.157 ;
		RECT	134.958 43.125 134.99 43.157 ;
		RECT	133.95 43.125 133.982 43.157 ;
		RECT	147.054 44.026 147.086 44.09 ;
		RECT	143.358 44.026 143.39 44.09 ;
		RECT	129.918 44.026 129.95 44.09 ;
		RECT	128.574 44.026 128.606 44.09 ;
		RECT	126.558 44.026 126.59 44.09 ;
		RECT	103.791 44.026 103.823 44.09 ;
		RECT	147.309 32.691 147.373 32.755 ;
		RECT	147.702 39.399 147.734 39.431 ;
		RECT	147.529 41.87 147.561 41.902 ;
		RECT	147.639 42.425 147.671 42.457 ;
		RECT	147.919 43.431 147.951 43.495 ;
		RECT	147.325 44.026 147.357 44.09 ;
		RECT	125.555 44.026 125.587 44.09 ;
		RECT	125.219 44.026 125.251 44.09 ;
		RECT	122.195 44.026 122.227 44.09 ;
		RECT	121.859 44.026 121.891 44.09 ;
		RECT	121.523 44.026 121.555 44.09 ;
		RECT	121.187 44.026 121.219 44.09 ;
		RECT	120.851 44.026 120.883 44.09 ;
		RECT	120.515 44.026 120.547 44.09 ;
		RECT	120.179 44.026 120.211 44.09 ;
		RECT	119.843 44.026 119.875 44.09 ;
		RECT	119.507 44.026 119.539 44.09 ;
		RECT	119.171 44.026 119.203 44.09 ;
		RECT	124.883 44.026 124.915 44.09 ;
		RECT	118.835 44.026 118.867 44.09 ;
		RECT	118.499 44.026 118.531 44.09 ;
		RECT	118.163 44.026 118.195 44.09 ;
		RECT	117.827 44.026 117.859 44.09 ;
		RECT	117.491 44.026 117.523 44.09 ;
		RECT	117.155 44.026 117.187 44.09 ;
		RECT	116.819 44.026 116.851 44.09 ;
		RECT	116.483 44.026 116.515 44.09 ;
		RECT	116.147 44.026 116.179 44.09 ;
		RECT	115.811 44.026 115.843 44.09 ;
		RECT	124.547 44.026 124.579 44.09 ;
		RECT	115.475 44.026 115.507 44.09 ;
		RECT	115.139 44.026 115.171 44.09 ;
		RECT	114.803 44.026 114.835 44.09 ;
		RECT	114.467 44.026 114.499 44.09 ;
		RECT	114.131 44.026 114.163 44.09 ;
		RECT	113.795 44.026 113.827 44.09 ;
		RECT	113.459 44.026 113.491 44.09 ;
		RECT	113.123 44.026 113.155 44.09 ;
		RECT	112.787 44.026 112.819 44.09 ;
		RECT	112.451 44.026 112.483 44.09 ;
		RECT	124.211 44.026 124.243 44.09 ;
		RECT	112.115 44.026 112.147 44.09 ;
		RECT	111.779 44.026 111.811 44.09 ;
		RECT	111.443 44.026 111.475 44.09 ;
		RECT	111.107 44.026 111.139 44.09 ;
		RECT	110.771 44.026 110.803 44.09 ;
		RECT	110.435 44.026 110.467 44.09 ;
		RECT	110.099 44.026 110.131 44.09 ;
		RECT	109.763 44.026 109.795 44.09 ;
		RECT	109.427 44.026 109.459 44.09 ;
		RECT	109.091 44.026 109.123 44.09 ;
		RECT	123.875 44.026 123.907 44.09 ;
		RECT	108.755 44.026 108.787 44.09 ;
		RECT	108.419 44.026 108.451 44.09 ;
		RECT	108.083 44.026 108.115 44.09 ;
		RECT	107.747 44.026 107.779 44.09 ;
		RECT	107.411 44.026 107.443 44.09 ;
		RECT	107.075 44.026 107.107 44.09 ;
		RECT	106.739 44.026 106.771 44.09 ;
		RECT	106.403 44.026 106.435 44.09 ;
		RECT	106.067 44.026 106.099 44.09 ;
		RECT	105.731 44.026 105.763 44.09 ;
		RECT	123.539 44.026 123.571 44.09 ;
		RECT	105.395 44.026 105.427 44.09 ;
		RECT	105.059 44.026 105.091 44.09 ;
		RECT	104.723 44.026 104.755 44.09 ;
		RECT	123.203 44.026 123.235 44.09 ;
		RECT	122.867 44.026 122.899 44.09 ;
		RECT	122.531 44.026 122.563 44.09 ;
		RECT	146.765 33.488 146.797 33.552 ;
		RECT	126.269 33.488 126.301 33.552 ;
		RECT	147.101 33.65 147.133 33.714 ;
		RECT	125.933 33.65 125.965 33.714 ;
		RECT	146.093 33.896 146.125 33.928 ;
		RECT	146.765 34.641 146.797 34.673 ;
		RECT	126.269 34.641 126.301 34.673 ;
		RECT	147.101 34.721 147.133 34.753 ;
		RECT	125.933 34.721 125.965 34.753 ;
		RECT	142.35 39.158 142.382 39.19 ;
		RECT	136.974 39.158 137.006 39.19 ;
		RECT	133.614 39.158 133.646 39.19 ;
		RECT	131.598 39.158 131.63 39.19 ;
		RECT	126.222 39.158 126.254 39.19 ;
		RECT	147.089 39.187 147.121 39.251 ;
		RECT	146.518 39.187 146.582 39.251 ;
		RECT	146.382 39.187 146.414 39.251 ;
		RECT	145.038 39.187 145.07 39.251 ;
		RECT	144.366 39.187 144.398 39.251 ;
		RECT	143.022 39.258 143.054 39.29 ;
		RECT	137.31 39.258 137.342 39.29 ;
		RECT	134.286 39.258 134.318 39.29 ;
		RECT	131.934 39.258 131.966 39.29 ;
		RECT	126.894 39.258 126.926 39.29 ;
		RECT	143.694 39.358 143.726 39.39 ;
		RECT	134.622 39.358 134.654 39.39 ;
		RECT	132.942 39.358 132.974 39.39 ;
		RECT	127.566 39.358 127.598 39.39 ;
		RECT	147.089 39.413 147.121 39.477 ;
		RECT	146.518 39.413 146.582 39.477 ;
		RECT	146.382 39.413 146.414 39.477 ;
		RECT	144.366 39.458 144.398 39.49 ;
		RECT	134.958 39.458 134.99 39.49 ;
		RECT	133.614 39.458 133.646 39.49 ;
		RECT	128.238 39.458 128.27 39.49 ;
		RECT	145.038 39.558 145.07 39.59 ;
		RECT	139.662 39.558 139.694 39.59 ;
		RECT	137.982 39.558 138.014 39.59 ;
		RECT	134.286 39.558 134.318 39.59 ;
		RECT	128.91 39.558 128.942 39.59 ;
		RECT	145.374 39.658 145.406 39.69 ;
		RECT	139.998 39.658 140.03 39.69 ;
		RECT	138.318 39.658 138.35 39.69 ;
		RECT	134.958 39.658 134.99 39.69 ;
		RECT	129.582 39.658 129.614 39.69 ;
		RECT	146.382 39.758 146.414 39.79 ;
		RECT	141.006 39.758 141.038 39.79 ;
		RECT	138.654 39.758 138.686 39.79 ;
		RECT	135.63 39.758 135.662 39.79 ;
		RECT	130.254 39.758 130.286 39.79 ;
		RECT	147.089 39.858 147.121 39.89 ;
		RECT	141.678 39.858 141.71 39.89 ;
		RECT	138.99 39.858 139.022 39.89 ;
		RECT	135.966 39.858 135.998 39.89 ;
		RECT	130.926 39.858 130.958 39.89 ;
		RECT	146.382 41.87 146.414 41.902 ;
		RECT	145.038 42.425 145.07 42.457 ;
		RECT	139.662 42.425 139.694 42.457 ;
		RECT	146.518 42.454 146.582 42.518 ;
		RECT	138.654 42.525 138.686 42.557 ;
		RECT	137.982 42.625 138.014 42.657 ;
		RECT	133.278 42.625 133.31 42.657 ;
		RECT	141.678 42.649 141.71 42.713 ;
		RECT	140.67 42.649 140.702 42.713 ;
		RECT	139.326 42.649 139.358 42.713 ;
		RECT	146.518 42.659 146.582 42.723 ;
		RECT	145.038 42.659 145.07 42.723 ;
		RECT	144.03 42.659 144.062 42.723 ;
		RECT	137.31 42.725 137.342 42.757 ;
		RECT	130.59 42.725 130.622 42.757 ;
		RECT	135.962 42.825 135.994 42.857 ;
		RECT	141.678 42.854 141.71 42.918 ;
		RECT	140.67 42.854 140.702 42.918 ;
		RECT	139.326 42.854 139.358 42.918 ;
		RECT	138.318 42.854 138.35 42.918 ;
		RECT	136.638 42.859 136.67 42.923 ;
		RECT	136.302 42.859 136.334 42.923 ;
		RECT	146.518 42.864 146.582 42.928 ;
		RECT	145.038 42.864 145.07 42.928 ;
		RECT	144.03 42.864 144.062 42.928 ;
		RECT	135.626 42.925 135.658 42.957 ;
		RECT	143.022 43.025 143.054 43.057 ;
		RECT	142.35 43.025 142.382 43.057 ;
		RECT	141.342 43.025 141.374 43.057 ;
		RECT	141.006 43.025 141.038 43.057 ;
		RECT	140.334 43.025 140.366 43.057 ;
		RECT	139.998 43.025 140.03 43.057 ;
		RECT	138.99 43.025 139.022 43.057 ;
		RECT	137.646 43.025 137.678 43.057 ;
		RECT	136.974 43.025 137.006 43.057 ;
		RECT	134.622 43.025 134.654 43.057 ;
		RECT	134.282 43.025 134.314 43.057 ;
		RECT	146.534 43.069 146.566 43.133 ;
		RECT	145.038 43.069 145.07 43.133 ;
		RECT	144.03 43.069 144.062 43.133 ;
		RECT	143.358 43.125 143.39 43.157 ;
		RECT	142.686 43.125 142.718 43.157 ;
		RECT	142.014 43.125 142.046 43.157 ;
		RECT	135.294 43.125 135.326 43.157 ;
		RECT	133.614 43.125 133.646 43.157 ;
		RECT	133.274 43.125 133.306 43.157 ;
		RECT	146.534 44.026 146.566 44.09 ;
		RECT	145.038 44.026 145.07 44.09 ;
		RECT	144.03 44.026 144.062 44.09 ;
		RECT	141.678 44.026 141.71 44.09 ;
		RECT	140.67 44.026 140.702 44.09 ;
		RECT	139.326 44.026 139.358 44.09 ;
		RECT	138.318 44.026 138.35 44.09 ;
		RECT	137.646 44.026 137.678 44.09 ;
		RECT	136.638 44.026 136.67 44.09 ;
		RECT	136.302 44.026 136.334 44.09 ;
		RECT	135.294 44.026 135.326 44.09 ;
		RECT	134.958 44.026 134.99 44.09 ;
		RECT	133.95 44.026 133.982 44.09 ;
		RECT	133.614 44.026 133.646 44.09 ;
		RECT	132.606 44.026 132.638 44.09 ;
		RECT	132.27 44.026 132.302 44.09 ;
		RECT	130.59 44.026 130.622 44.09 ;
		RECT	129.582 44.026 129.614 44.09 ;
		RECT	128.91 44.026 128.942 44.09 ;
		RECT	128.238 44.026 128.27 44.09 ;
		RECT	127.902 44.026 127.934 44.09 ;
		RECT	127.566 44.026 127.598 44.09 ;
		RECT	127.23 44.026 127.262 44.09 ;
		RECT	125.886 44.026 125.918 44.09 ;
		RECT	103.787 43.431 103.819 43.495 ;
		RECT	104.387 44.026 104.419 44.09 ;
		RECT	200.624 31.762 200.688 31.794 ;
		RECT	200.624 50.382 200.688 50.414 ;
		RECT	178.613 39.858 178.645 39.89 ;
		RECT	181.973 39.358 182.005 39.39 ;
		RECT	182.309 39.358 182.341 39.39 ;
		RECT	182.645 39.258 182.677 39.29 ;
		RECT	182.981 39.258 183.013 39.29 ;
		RECT	183.317 39.158 183.349 39.19 ;
		RECT	183.653 39.158 183.685 39.19 ;
		RECT	183.989 39.858 184.021 39.89 ;
		RECT	184.325 39.858 184.357 39.89 ;
		RECT	184.661 39.758 184.693 39.79 ;
		RECT	184.997 39.758 185.029 39.79 ;
		RECT	178.949 39.858 178.981 39.89 ;
		RECT	185.333 39.658 185.365 39.69 ;
		RECT	185.669 39.658 185.701 39.69 ;
		RECT	186.005 39.558 186.037 39.59 ;
		RECT	186.341 39.558 186.373 39.59 ;
		RECT	186.677 39.458 186.709 39.49 ;
		RECT	187.013 39.458 187.045 39.49 ;
		RECT	187.349 39.358 187.381 39.39 ;
		RECT	187.685 39.358 187.717 39.39 ;
		RECT	188.021 39.258 188.053 39.29 ;
		RECT	188.357 39.258 188.389 39.29 ;
		RECT	179.285 39.758 179.317 39.79 ;
		RECT	188.693 39.158 188.725 39.19 ;
		RECT	189.029 39.158 189.061 39.19 ;
		RECT	189.365 39.858 189.397 39.89 ;
		RECT	189.701 39.858 189.733 39.89 ;
		RECT	190.037 39.758 190.069 39.79 ;
		RECT	190.373 39.758 190.405 39.79 ;
		RECT	190.709 39.658 190.741 39.69 ;
		RECT	191.045 39.658 191.077 39.69 ;
		RECT	191.381 39.558 191.413 39.59 ;
		RECT	191.717 39.558 191.749 39.59 ;
		RECT	179.621 39.758 179.653 39.79 ;
		RECT	192.053 39.458 192.085 39.49 ;
		RECT	192.389 39.458 192.421 39.49 ;
		RECT	192.725 39.358 192.757 39.39 ;
		RECT	193.061 39.358 193.093 39.39 ;
		RECT	193.397 39.258 193.429 39.29 ;
		RECT	193.733 39.258 193.765 39.29 ;
		RECT	194.069 39.158 194.101 39.19 ;
		RECT	194.405 39.158 194.437 39.19 ;
		RECT	194.741 39.858 194.773 39.89 ;
		RECT	195.077 39.858 195.109 39.89 ;
		RECT	179.957 39.658 179.989 39.69 ;
		RECT	195.413 39.758 195.445 39.79 ;
		RECT	195.749 39.758 195.781 39.79 ;
		RECT	196.085 39.658 196.117 39.69 ;
		RECT	196.421 39.658 196.453 39.69 ;
		RECT	196.757 39.558 196.789 39.59 ;
		RECT	197.093 39.558 197.125 39.59 ;
		RECT	197.429 39.458 197.461 39.49 ;
		RECT	197.765 39.458 197.797 39.49 ;
		RECT	198.101 39.358 198.133 39.39 ;
		RECT	198.437 39.358 198.469 39.39 ;
		RECT	180.293 39.658 180.325 39.69 ;
		RECT	198.773 39.258 198.805 39.29 ;
		RECT	199.109 39.258 199.141 39.29 ;
		RECT	199.445 39.158 199.477 39.19 ;
		RECT	199.781 39.158 199.813 39.19 ;
		RECT	180.629 39.558 180.661 39.59 ;
		RECT	180.965 39.558 180.997 39.59 ;
		RECT	181.301 39.458 181.333 39.49 ;
		RECT	181.637 39.458 181.669 39.49 ;
		RECT	178.613 42.825 178.645 42.857 ;
		RECT	181.973 42.825 182.005 42.857 ;
		RECT	182.309 42.825 182.341 42.857 ;
		RECT	182.645 42.825 182.677 42.857 ;
		RECT	182.981 42.825 183.013 42.857 ;
		RECT	183.317 42.825 183.349 42.857 ;
		RECT	183.653 42.825 183.685 42.857 ;
		RECT	183.989 42.925 184.021 42.957 ;
		RECT	184.325 42.925 184.357 42.957 ;
		RECT	184.661 42.925 184.693 42.957 ;
		RECT	184.997 42.925 185.029 42.957 ;
		RECT	178.949 42.825 178.981 42.857 ;
		RECT	185.333 42.925 185.365 42.957 ;
		RECT	185.669 42.925 185.701 42.957 ;
		RECT	186.005 42.925 186.037 42.957 ;
		RECT	186.341 42.925 186.373 42.957 ;
		RECT	186.677 42.925 186.709 42.957 ;
		RECT	187.013 42.925 187.045 42.957 ;
		RECT	187.349 42.925 187.381 42.957 ;
		RECT	187.685 42.925 187.717 42.957 ;
		RECT	188.021 42.925 188.053 42.957 ;
		RECT	188.357 42.925 188.389 42.957 ;
		RECT	179.285 42.825 179.317 42.857 ;
		RECT	188.693 42.925 188.725 42.957 ;
		RECT	189.029 42.925 189.061 42.957 ;
		RECT	189.365 43.025 189.397 43.057 ;
		RECT	189.701 43.025 189.733 43.057 ;
		RECT	190.037 43.025 190.069 43.057 ;
		RECT	190.373 43.025 190.405 43.057 ;
		RECT	190.709 43.025 190.741 43.057 ;
		RECT	191.045 43.025 191.077 43.057 ;
		RECT	191.381 43.025 191.413 43.057 ;
		RECT	191.717 43.025 191.749 43.057 ;
		RECT	179.621 42.825 179.653 42.857 ;
		RECT	192.053 43.025 192.085 43.057 ;
		RECT	192.389 43.025 192.421 43.057 ;
		RECT	192.725 43.025 192.757 43.057 ;
		RECT	193.061 43.025 193.093 43.057 ;
		RECT	193.397 43.025 193.429 43.057 ;
		RECT	193.733 43.025 193.765 43.057 ;
		RECT	194.069 43.025 194.101 43.057 ;
		RECT	194.405 43.025 194.437 43.057 ;
		RECT	194.741 43.125 194.773 43.157 ;
		RECT	195.077 43.125 195.109 43.157 ;
		RECT	179.957 42.825 179.989 42.857 ;
		RECT	195.413 43.125 195.445 43.157 ;
		RECT	195.749 43.125 195.781 43.157 ;
		RECT	196.085 43.125 196.117 43.157 ;
		RECT	196.421 43.125 196.453 43.157 ;
		RECT	196.757 43.125 196.789 43.157 ;
		RECT	197.093 43.125 197.125 43.157 ;
		RECT	197.429 43.125 197.461 43.157 ;
		RECT	197.765 43.125 197.797 43.157 ;
		RECT	198.101 43.125 198.133 43.157 ;
		RECT	198.437 43.125 198.469 43.157 ;
		RECT	180.293 42.825 180.325 42.857 ;
		RECT	198.773 43.125 198.805 43.157 ;
		RECT	199.109 43.125 199.141 43.157 ;
		RECT	199.445 43.125 199.477 43.157 ;
		RECT	199.781 43.125 199.813 43.157 ;
		RECT	180.629 42.825 180.661 42.857 ;
		RECT	180.965 42.825 180.997 42.857 ;
		RECT	181.301 42.825 181.333 42.857 ;
		RECT	181.637 42.825 181.669 42.857 ;
		RECT	178.655 32.691 178.687 32.755 ;
		RECT	156.459 39.672 156.491 39.736 ;
		RECT	156.495 44.026 156.527 44.09 ;
		RECT	182.015 32.691 182.047 32.755 ;
		RECT	182.351 32.691 182.383 32.755 ;
		RECT	182.687 32.691 182.719 32.755 ;
		RECT	183.023 32.691 183.055 32.755 ;
		RECT	183.359 32.691 183.391 32.755 ;
		RECT	183.695 32.691 183.727 32.755 ;
		RECT	184.031 32.691 184.063 32.755 ;
		RECT	184.367 32.691 184.399 32.755 ;
		RECT	184.703 32.691 184.735 32.755 ;
		RECT	185.039 32.691 185.071 32.755 ;
		RECT	178.991 32.691 179.023 32.755 ;
		RECT	185.375 32.691 185.407 32.755 ;
		RECT	185.711 32.691 185.743 32.755 ;
		RECT	186.047 32.691 186.079 32.755 ;
		RECT	186.383 32.691 186.415 32.755 ;
		RECT	186.719 32.691 186.751 32.755 ;
		RECT	187.055 32.691 187.087 32.755 ;
		RECT	187.391 32.691 187.423 32.755 ;
		RECT	187.727 32.691 187.759 32.755 ;
		RECT	188.063 32.691 188.095 32.755 ;
		RECT	188.399 32.691 188.431 32.755 ;
		RECT	179.327 32.691 179.359 32.755 ;
		RECT	188.735 32.691 188.767 32.755 ;
		RECT	189.071 32.691 189.103 32.755 ;
		RECT	189.407 32.691 189.439 32.755 ;
		RECT	189.743 32.691 189.775 32.755 ;
		RECT	190.079 32.691 190.111 32.755 ;
		RECT	190.415 32.691 190.447 32.755 ;
		RECT	190.751 32.691 190.783 32.755 ;
		RECT	191.087 32.691 191.119 32.755 ;
		RECT	191.423 32.691 191.455 32.755 ;
		RECT	191.759 32.691 191.791 32.755 ;
		RECT	179.663 32.691 179.695 32.755 ;
		RECT	192.095 32.691 192.127 32.755 ;
		RECT	192.431 32.691 192.463 32.755 ;
		RECT	192.767 32.691 192.799 32.755 ;
		RECT	193.103 32.691 193.135 32.755 ;
		RECT	193.439 32.691 193.471 32.755 ;
		RECT	193.775 32.691 193.807 32.755 ;
		RECT	194.111 32.691 194.143 32.755 ;
		RECT	194.447 32.691 194.479 32.755 ;
		RECT	194.783 32.691 194.815 32.755 ;
		RECT	195.119 32.691 195.151 32.755 ;
		RECT	179.999 32.691 180.031 32.755 ;
		RECT	195.455 32.691 195.487 32.755 ;
		RECT	195.791 32.691 195.823 32.755 ;
		RECT	196.127 32.691 196.159 32.755 ;
		RECT	196.463 32.691 196.495 32.755 ;
		RECT	196.799 32.691 196.831 32.755 ;
		RECT	197.135 32.691 197.167 32.755 ;
		RECT	197.471 32.691 197.503 32.755 ;
		RECT	197.807 32.691 197.839 32.755 ;
		RECT	198.143 32.691 198.175 32.755 ;
		RECT	198.479 32.691 198.511 32.755 ;
		RECT	180.335 32.691 180.367 32.755 ;
		RECT	198.815 32.691 198.847 32.755 ;
		RECT	199.151 32.691 199.183 32.755 ;
		RECT	199.487 32.691 199.519 32.755 ;
		RECT	199.823 32.691 199.855 32.755 ;
		RECT	180.671 32.691 180.703 32.755 ;
		RECT	181.007 32.691 181.039 32.755 ;
		RECT	181.343 32.691 181.375 32.755 ;
		RECT	181.679 32.691 181.711 32.755 ;
		RECT	162.49 43.125 162.522 43.157 ;
		RECT	163.498 43.125 163.53 43.157 ;
		RECT	164.842 43.125 164.874 43.157 ;
		RECT	165.85 43.125 165.882 43.157 ;
		RECT	167.53 43.125 167.562 43.157 ;
		RECT	167.866 43.125 167.898 43.157 ;
		RECT	169.21 43.125 169.242 43.157 ;
		RECT	170.218 43.125 170.25 43.157 ;
		RECT	157.114 44.026 157.146 44.09 ;
		RECT	160.81 44.026 160.842 44.09 ;
		RECT	174.25 44.026 174.282 44.09 ;
		RECT	175.594 44.026 175.626 44.09 ;
		RECT	177.61 44.026 177.642 44.09 ;
		RECT	200.377 44.026 200.409 44.09 ;
		RECT	156.827 32.691 156.891 32.755 ;
		RECT	156.466 39.399 156.498 39.431 ;
		RECT	156.639 41.87 156.671 41.902 ;
		RECT	156.529 42.425 156.561 42.457 ;
		RECT	156.249 43.431 156.281 43.495 ;
		RECT	156.843 44.026 156.875 44.09 ;
		RECT	178.613 44.026 178.645 44.09 ;
		RECT	178.949 44.026 178.981 44.09 ;
		RECT	181.973 44.026 182.005 44.09 ;
		RECT	182.309 44.026 182.341 44.09 ;
		RECT	182.645 44.026 182.677 44.09 ;
		RECT	182.981 44.026 183.013 44.09 ;
		RECT	183.317 44.026 183.349 44.09 ;
		RECT	183.653 44.026 183.685 44.09 ;
		RECT	183.989 44.026 184.021 44.09 ;
		RECT	184.325 44.026 184.357 44.09 ;
		RECT	184.661 44.026 184.693 44.09 ;
		RECT	184.997 44.026 185.029 44.09 ;
		RECT	179.285 44.026 179.317 44.09 ;
		RECT	185.333 44.026 185.365 44.09 ;
		RECT	185.669 44.026 185.701 44.09 ;
		RECT	186.005 44.026 186.037 44.09 ;
		RECT	186.341 44.026 186.373 44.09 ;
		RECT	186.677 44.026 186.709 44.09 ;
		RECT	187.013 44.026 187.045 44.09 ;
		RECT	187.349 44.026 187.381 44.09 ;
		RECT	187.685 44.026 187.717 44.09 ;
		RECT	188.021 44.026 188.053 44.09 ;
		RECT	188.357 44.026 188.389 44.09 ;
		RECT	179.621 44.026 179.653 44.09 ;
		RECT	188.693 44.026 188.725 44.09 ;
		RECT	189.029 44.026 189.061 44.09 ;
		RECT	189.365 44.026 189.397 44.09 ;
		RECT	189.701 44.026 189.733 44.09 ;
		RECT	190.037 44.026 190.069 44.09 ;
		RECT	190.373 44.026 190.405 44.09 ;
		RECT	190.709 44.026 190.741 44.09 ;
		RECT	191.045 44.026 191.077 44.09 ;
		RECT	191.381 44.026 191.413 44.09 ;
		RECT	191.717 44.026 191.749 44.09 ;
		RECT	179.957 44.026 179.989 44.09 ;
		RECT	192.053 44.026 192.085 44.09 ;
		RECT	192.389 44.026 192.421 44.09 ;
		RECT	192.725 44.026 192.757 44.09 ;
		RECT	193.061 44.026 193.093 44.09 ;
		RECT	193.397 44.026 193.429 44.09 ;
		RECT	193.733 44.026 193.765 44.09 ;
		RECT	194.069 44.026 194.101 44.09 ;
		RECT	194.405 44.026 194.437 44.09 ;
		RECT	194.741 44.026 194.773 44.09 ;
		RECT	195.077 44.026 195.109 44.09 ;
		RECT	180.293 44.026 180.325 44.09 ;
		RECT	195.413 44.026 195.445 44.09 ;
		RECT	195.749 44.026 195.781 44.09 ;
		RECT	196.085 44.026 196.117 44.09 ;
		RECT	196.421 44.026 196.453 44.09 ;
		RECT	196.757 44.026 196.789 44.09 ;
		RECT	197.093 44.026 197.125 44.09 ;
		RECT	197.429 44.026 197.461 44.09 ;
		RECT	197.765 44.026 197.797 44.09 ;
		RECT	198.101 44.026 198.133 44.09 ;
		RECT	198.437 44.026 198.469 44.09 ;
		RECT	180.629 44.026 180.661 44.09 ;
		RECT	198.773 44.026 198.805 44.09 ;
		RECT	199.109 44.026 199.141 44.09 ;
		RECT	199.445 44.026 199.477 44.09 ;
		RECT	180.965 44.026 180.997 44.09 ;
		RECT	181.301 44.026 181.333 44.09 ;
		RECT	181.637 44.026 181.669 44.09 ;
		RECT	157.403 33.488 157.435 33.552 ;
		RECT	177.899 33.488 177.931 33.552 ;
		RECT	157.067 33.65 157.099 33.714 ;
		RECT	178.235 33.65 178.267 33.714 ;
		RECT	158.075 33.896 158.107 33.928 ;
		RECT	157.403 34.641 157.435 34.673 ;
		RECT	177.899 34.641 177.931 34.673 ;
		RECT	157.067 34.721 157.099 34.753 ;
		RECT	178.235 34.721 178.267 34.753 ;
		RECT	161.818 39.158 161.85 39.19 ;
		RECT	167.194 39.158 167.226 39.19 ;
		RECT	170.554 39.158 170.586 39.19 ;
		RECT	172.57 39.158 172.602 39.19 ;
		RECT	177.946 39.158 177.978 39.19 ;
		RECT	157.079 39.187 157.111 39.251 ;
		RECT	157.618 39.187 157.682 39.251 ;
		RECT	157.786 39.187 157.818 39.251 ;
		RECT	159.13 39.187 159.162 39.251 ;
		RECT	159.802 39.187 159.834 39.251 ;
		RECT	161.146 39.258 161.178 39.29 ;
		RECT	166.858 39.258 166.89 39.29 ;
		RECT	169.882 39.258 169.914 39.29 ;
		RECT	172.234 39.258 172.266 39.29 ;
		RECT	177.274 39.258 177.306 39.29 ;
		RECT	160.474 39.358 160.506 39.39 ;
		RECT	169.546 39.358 169.578 39.39 ;
		RECT	171.226 39.358 171.258 39.39 ;
		RECT	176.602 39.358 176.634 39.39 ;
		RECT	157.079 39.413 157.111 39.477 ;
		RECT	157.618 39.413 157.682 39.477 ;
		RECT	157.786 39.413 157.818 39.477 ;
		RECT	159.802 39.458 159.834 39.49 ;
		RECT	169.21 39.458 169.242 39.49 ;
		RECT	170.554 39.458 170.586 39.49 ;
		RECT	175.93 39.458 175.962 39.49 ;
		RECT	159.13 39.558 159.162 39.59 ;
		RECT	164.506 39.558 164.538 39.59 ;
		RECT	166.186 39.558 166.218 39.59 ;
		RECT	169.882 39.558 169.914 39.59 ;
		RECT	175.258 39.558 175.29 39.59 ;
		RECT	158.794 39.658 158.826 39.69 ;
		RECT	164.17 39.658 164.202 39.69 ;
		RECT	165.85 39.658 165.882 39.69 ;
		RECT	169.21 39.658 169.242 39.69 ;
		RECT	174.586 39.658 174.618 39.69 ;
		RECT	157.786 39.758 157.818 39.79 ;
		RECT	163.162 39.758 163.194 39.79 ;
		RECT	165.514 39.758 165.546 39.79 ;
		RECT	168.538 39.758 168.57 39.79 ;
		RECT	173.914 39.758 173.946 39.79 ;
		RECT	157.079 39.858 157.111 39.89 ;
		RECT	162.49 39.858 162.522 39.89 ;
		RECT	165.178 39.858 165.21 39.89 ;
		RECT	168.202 39.858 168.234 39.89 ;
		RECT	173.242 39.858 173.274 39.89 ;
		RECT	157.786 41.87 157.818 41.902 ;
		RECT	159.13 42.425 159.162 42.457 ;
		RECT	164.506 42.425 164.538 42.457 ;
		RECT	157.618 42.454 157.682 42.518 ;
		RECT	165.514 42.525 165.546 42.557 ;
		RECT	166.186 42.625 166.218 42.657 ;
		RECT	170.89 42.625 170.922 42.657 ;
		RECT	162.49 42.649 162.522 42.713 ;
		RECT	163.498 42.649 163.53 42.713 ;
		RECT	164.842 42.649 164.874 42.713 ;
		RECT	157.618 42.659 157.682 42.723 ;
		RECT	159.13 42.659 159.162 42.723 ;
		RECT	160.138 42.659 160.17 42.723 ;
		RECT	166.858 42.725 166.89 42.757 ;
		RECT	173.578 42.725 173.61 42.757 ;
		RECT	168.206 42.825 168.238 42.857 ;
		RECT	162.49 42.854 162.522 42.918 ;
		RECT	163.498 42.854 163.53 42.918 ;
		RECT	164.842 42.854 164.874 42.918 ;
		RECT	165.85 42.854 165.882 42.918 ;
		RECT	167.53 42.859 167.562 42.923 ;
		RECT	167.866 42.859 167.898 42.923 ;
		RECT	157.618 42.864 157.682 42.928 ;
		RECT	159.13 42.864 159.162 42.928 ;
		RECT	160.138 42.864 160.17 42.928 ;
		RECT	168.542 42.925 168.574 42.957 ;
		RECT	161.146 43.025 161.178 43.057 ;
		RECT	161.818 43.025 161.85 43.057 ;
		RECT	162.826 43.025 162.858 43.057 ;
		RECT	163.162 43.025 163.194 43.057 ;
		RECT	163.834 43.025 163.866 43.057 ;
		RECT	164.17 43.025 164.202 43.057 ;
		RECT	165.178 43.025 165.21 43.057 ;
		RECT	166.522 43.025 166.554 43.057 ;
		RECT	167.194 43.025 167.226 43.057 ;
		RECT	169.546 43.025 169.578 43.057 ;
		RECT	169.886 43.025 169.918 43.057 ;
		RECT	157.634 43.069 157.666 43.133 ;
		RECT	159.13 43.069 159.162 43.133 ;
		RECT	160.138 43.069 160.17 43.133 ;
		RECT	160.81 43.125 160.842 43.157 ;
		RECT	161.482 43.125 161.514 43.157 ;
		RECT	162.154 43.125 162.186 43.157 ;
		RECT	168.874 43.125 168.906 43.157 ;
		RECT	170.554 43.125 170.586 43.157 ;
		RECT	170.894 43.125 170.926 43.157 ;
		RECT	157.634 44.026 157.666 44.09 ;
		RECT	159.13 44.026 159.162 44.09 ;
		RECT	160.138 44.026 160.17 44.09 ;
		RECT	162.49 44.026 162.522 44.09 ;
		RECT	163.498 44.026 163.53 44.09 ;
		RECT	164.842 44.026 164.874 44.09 ;
		RECT	165.85 44.026 165.882 44.09 ;
		RECT	166.522 44.026 166.554 44.09 ;
		RECT	167.53 44.026 167.562 44.09 ;
		RECT	167.866 44.026 167.898 44.09 ;
		RECT	168.874 44.026 168.906 44.09 ;
		RECT	169.21 44.026 169.242 44.09 ;
		RECT	170.218 44.026 170.25 44.09 ;
		RECT	170.554 44.026 170.586 44.09 ;
		RECT	171.562 44.026 171.594 44.09 ;
		RECT	171.898 44.026 171.93 44.09 ;
		RECT	173.578 44.026 173.61 44.09 ;
		RECT	174.586 44.026 174.618 44.09 ;
		RECT	175.258 44.026 175.29 44.09 ;
		RECT	175.93 44.026 175.962 44.09 ;
		RECT	176.266 44.026 176.298 44.09 ;
		RECT	176.602 44.026 176.634 44.09 ;
		RECT	176.938 44.026 176.97 44.09 ;
		RECT	178.282 44.026 178.314 44.09 ;
		RECT	200.381 43.431 200.413 43.495 ;
		RECT	199.781 44.026 199.813 44.09 ;
		RECT	201.156 31.746 201.188 31.81 ;
		RECT	201.403 32.691 201.435 32.755 ;
		LAYER	M1 DESIGNRULEWIDTH 0.032 ;
		RECT	0.134 0.206 201.531 81.97 ;
		RECT	0 0 0.134 82.176 ;
		RECT	201.531 0 201.665 82.176 ;
		RECT	0.134 0 201.531 0.206 ;
		RECT	0.134 81.97 201.531 82.176 ;
		LAYER	M2 DESIGNRULEWIDTH 0.032 ;
		RECT	0.134 0.206 201.531 81.97 ;
		RECT	0 0 0.134 0.876 ;
		RECT	0 1.092 0.134 1.359 ;
		RECT	0 1.575 0.134 2.22 ;
		RECT	0 2.436 0.134 2.796 ;
		RECT	0 3.012 0.134 3.279 ;
		RECT	0 3.495 0.134 4.14 ;
		RECT	0 4.356 0.134 4.716 ;
		RECT	0 4.932 0.134 5.199 ;
		RECT	0 5.415 0.134 6.06 ;
		RECT	0 6.276 0.134 6.636 ;
		RECT	0 6.852 0.134 7.119 ;
		RECT	0 7.335 0.134 7.98 ;
		RECT	0 8.196 0.134 8.556 ;
		RECT	0 8.772 0.134 9.039 ;
		RECT	0 9.255 0.134 9.9 ;
		RECT	0 10.116 0.134 10.476 ;
		RECT	0 10.692 0.134 10.959 ;
		RECT	0 11.175 0.134 11.82 ;
		RECT	0 12.036 0.134 12.396 ;
		RECT	0 12.612 0.134 12.879 ;
		RECT	0 13.095 0.134 13.74 ;
		RECT	0 13.956 0.134 14.316 ;
		RECT	0 14.532 0.134 14.799 ;
		RECT	0 15.015 0.134 15.66 ;
		RECT	0 15.876 0.134 16.236 ;
		RECT	0 16.452 0.134 16.719 ;
		RECT	0 16.935 0.134 17.58 ;
		RECT	0 17.796 0.134 18.156 ;
		RECT	0 18.372 0.134 18.639 ;
		RECT	0 18.855 0.134 19.5 ;
		RECT	0 19.716 0.134 20.076 ;
		RECT	0 20.292 0.134 20.559 ;
		RECT	0 20.775 0.134 21.42 ;
		RECT	0 21.636 0.134 21.996 ;
		RECT	0 22.212 0.134 22.479 ;
		RECT	0 22.695 0.134 23.34 ;
		RECT	0 23.556 0.134 23.916 ;
		RECT	0 24.132 0.134 24.399 ;
		RECT	0 24.615 0.134 25.26 ;
		RECT	0 25.476 0.134 25.836 ;
		RECT	0 26.052 0.134 26.319 ;
		RECT	0 26.535 0.134 27.18 ;
		RECT	0 27.396 0.134 27.756 ;
		RECT	0 27.972 0.134 28.239 ;
		RECT	0 28.455 0.134 29.1 ;
		RECT	0 29.316 0.134 29.676 ;
		RECT	0 29.892 0.134 30.159 ;
		RECT	0 30.375 0.134 31.02 ;
		RECT	0 31.236 0.134 33.9 ;
		RECT	0 34.452 0.134 34.524 ;
		RECT	0 34.74 0.134 35.052 ;
		RECT	0 35.412 0.134 35.532 ;
		RECT	0 35.892 0.134 37.26 ;
		RECT	0 37.668 0.134 37.932 ;
		RECT	0 38.148 0.134 39.18 ;
		RECT	0 39.588 0.134 39.852 ;
		RECT	0 40.068 0.134 40.476 ;
		RECT	0 40.692 0.134 40.956 ;
		RECT	0 41.172 0.134 41.484 ;
		RECT	0 41.7 0.134 41.964 ;
		RECT	0 42.372 0.134 43.644 ;
		RECT	0 43.86 0.134 44.124 ;
		RECT	0 44.34 0.134 44.988 ;
		RECT	0 45.204 0.134 47.532 ;
		RECT	0 47.748 0.134 50.94 ;
		RECT	0 51.156 0.134 51.801 ;
		RECT	0 52.017 0.134 52.284 ;
		RECT	0 52.5 0.134 52.86 ;
		RECT	0 53.076 0.134 53.721 ;
		RECT	0 53.937 0.134 54.204 ;
		RECT	0 54.42 0.134 54.78 ;
		RECT	0 54.996 0.134 55.641 ;
		RECT	0 55.857 0.134 56.124 ;
		RECT	0 56.34 0.134 56.7 ;
		RECT	0 56.916 0.134 57.561 ;
		RECT	0 57.777 0.134 58.044 ;
		RECT	0 58.26 0.134 58.62 ;
		RECT	0 58.836 0.134 59.481 ;
		RECT	0 59.697 0.134 59.964 ;
		RECT	0 60.18 0.134 60.54 ;
		RECT	0 60.756 0.134 61.401 ;
		RECT	0 61.617 0.134 61.884 ;
		RECT	0 62.1 0.134 62.46 ;
		RECT	0 62.676 0.134 63.321 ;
		RECT	0 63.537 0.134 63.804 ;
		RECT	0 64.02 0.134 64.38 ;
		RECT	0 64.596 0.134 65.241 ;
		RECT	0 65.457 0.134 65.724 ;
		RECT	0 65.94 0.134 66.3 ;
		RECT	0 66.516 0.134 67.161 ;
		RECT	0 67.377 0.134 67.644 ;
		RECT	0 67.86 0.134 68.22 ;
		RECT	0 68.436 0.134 69.081 ;
		RECT	0 69.297 0.134 69.564 ;
		RECT	0 69.78 0.134 70.14 ;
		RECT	0 70.356 0.134 71.001 ;
		RECT	0 71.217 0.134 71.484 ;
		RECT	0 71.7 0.134 72.06 ;
		RECT	0 72.276 0.134 72.921 ;
		RECT	0 73.137 0.134 73.404 ;
		RECT	0 73.62 0.134 73.98 ;
		RECT	0 74.196 0.134 74.841 ;
		RECT	0 75.057 0.134 75.324 ;
		RECT	0 75.54 0.134 75.9 ;
		RECT	0 76.116 0.134 76.761 ;
		RECT	0 76.977 0.134 77.244 ;
		RECT	0 77.46 0.134 77.82 ;
		RECT	0 78.036 0.134 78.681 ;
		RECT	0 78.897 0.134 79.164 ;
		RECT	0 79.38 0.134 79.74 ;
		RECT	0 79.956 0.134 80.601 ;
		RECT	0 80.817 0.134 81.084 ;
		RECT	0 81.3 0.134 82.176 ;
		RECT	201.531 0 201.665 82.176 ;
		RECT	0.134 0 201.531 0.206 ;
		RECT	0.134 81.97 201.531 82.176 ;
		LAYER	M3 DESIGNRULEWIDTH 0.032 ;
		RECT	0.134 0.206 201.531 81.97 ;
		RECT	0 0 0.134 0.876 ;
		RECT	0 1.092 0.134 1.359 ;
		RECT	0 1.575 0.134 2.22 ;
		RECT	0 2.436 0.134 2.796 ;
		RECT	0 3.012 0.134 3.279 ;
		RECT	0 3.495 0.134 4.14 ;
		RECT	0 4.356 0.134 4.716 ;
		RECT	0 4.932 0.134 5.199 ;
		RECT	0 5.415 0.134 6.06 ;
		RECT	0 6.276 0.134 6.636 ;
		RECT	0 6.852 0.134 7.119 ;
		RECT	0 7.335 0.134 7.98 ;
		RECT	0 8.196 0.134 8.556 ;
		RECT	0 8.772 0.134 9.039 ;
		RECT	0 9.255 0.134 9.9 ;
		RECT	0 10.116 0.134 10.476 ;
		RECT	0 10.692 0.134 10.959 ;
		RECT	0 11.175 0.134 11.82 ;
		RECT	0 12.036 0.134 12.396 ;
		RECT	0 12.612 0.134 12.879 ;
		RECT	0 13.095 0.134 13.74 ;
		RECT	0 13.956 0.134 14.316 ;
		RECT	0 14.532 0.134 14.799 ;
		RECT	0 15.015 0.134 15.66 ;
		RECT	0 15.876 0.134 16.236 ;
		RECT	0 16.452 0.134 16.719 ;
		RECT	0 16.935 0.134 17.58 ;
		RECT	0 17.796 0.134 18.156 ;
		RECT	0 18.372 0.134 18.639 ;
		RECT	0 18.855 0.134 19.5 ;
		RECT	0 19.716 0.134 20.076 ;
		RECT	0 20.292 0.134 20.559 ;
		RECT	0 20.775 0.134 21.42 ;
		RECT	0 21.636 0.134 21.996 ;
		RECT	0 22.212 0.134 22.479 ;
		RECT	0 22.695 0.134 23.34 ;
		RECT	0 23.556 0.134 23.916 ;
		RECT	0 24.132 0.134 24.399 ;
		RECT	0 24.615 0.134 25.26 ;
		RECT	0 25.476 0.134 25.836 ;
		RECT	0 26.052 0.134 26.319 ;
		RECT	0 26.535 0.134 27.18 ;
		RECT	0 27.396 0.134 27.756 ;
		RECT	0 27.972 0.134 28.239 ;
		RECT	0 28.455 0.134 29.1 ;
		RECT	0 29.316 0.134 29.676 ;
		RECT	0 29.892 0.134 30.159 ;
		RECT	0 30.375 0.134 31.02 ;
		RECT	0 31.236 0.134 33.9 ;
		RECT	0 34.452 0.134 34.524 ;
		RECT	0 34.74 0.134 35.052 ;
		RECT	0 35.412 0.134 35.532 ;
		RECT	0 35.892 0.134 37.26 ;
		RECT	0 37.668 0.134 37.932 ;
		RECT	0 38.148 0.134 39.18 ;
		RECT	0 39.588 0.134 39.852 ;
		RECT	0 40.068 0.134 40.476 ;
		RECT	0 40.692 0.134 40.956 ;
		RECT	0 41.172 0.134 41.484 ;
		RECT	0 41.7 0.134 41.964 ;
		RECT	0 42.372 0.134 43.644 ;
		RECT	0 43.86 0.134 44.124 ;
		RECT	0 44.34 0.134 44.988 ;
		RECT	0 45.204 0.134 47.532 ;
		RECT	0 47.748 0.134 50.94 ;
		RECT	0 51.156 0.134 51.801 ;
		RECT	0 52.017 0.134 52.284 ;
		RECT	0 52.5 0.134 52.86 ;
		RECT	0 53.076 0.134 53.721 ;
		RECT	0 53.937 0.134 54.204 ;
		RECT	0 54.42 0.134 54.78 ;
		RECT	0 54.996 0.134 55.641 ;
		RECT	0 55.857 0.134 56.124 ;
		RECT	0 56.34 0.134 56.7 ;
		RECT	0 56.916 0.134 57.561 ;
		RECT	0 57.777 0.134 58.044 ;
		RECT	0 58.26 0.134 58.62 ;
		RECT	0 58.836 0.134 59.481 ;
		RECT	0 59.697 0.134 59.964 ;
		RECT	0 60.18 0.134 60.54 ;
		RECT	0 60.756 0.134 61.401 ;
		RECT	0 61.617 0.134 61.884 ;
		RECT	0 62.1 0.134 62.46 ;
		RECT	0 62.676 0.134 63.321 ;
		RECT	0 63.537 0.134 63.804 ;
		RECT	0 64.02 0.134 64.38 ;
		RECT	0 64.596 0.134 65.241 ;
		RECT	0 65.457 0.134 65.724 ;
		RECT	0 65.94 0.134 66.3 ;
		RECT	0 66.516 0.134 67.161 ;
		RECT	0 67.377 0.134 67.644 ;
		RECT	0 67.86 0.134 68.22 ;
		RECT	0 68.436 0.134 69.081 ;
		RECT	0 69.297 0.134 69.564 ;
		RECT	0 69.78 0.134 70.14 ;
		RECT	0 70.356 0.134 71.001 ;
		RECT	0 71.217 0.134 71.484 ;
		RECT	0 71.7 0.134 72.06 ;
		RECT	0 72.276 0.134 72.921 ;
		RECT	0 73.137 0.134 73.404 ;
		RECT	0 73.62 0.134 73.98 ;
		RECT	0 74.196 0.134 74.841 ;
		RECT	0 75.057 0.134 75.324 ;
		RECT	0 75.54 0.134 75.9 ;
		RECT	0 76.116 0.134 76.761 ;
		RECT	0 76.977 0.134 77.244 ;
		RECT	0 77.46 0.134 77.82 ;
		RECT	0 78.036 0.134 78.681 ;
		RECT	0 78.897 0.134 79.164 ;
		RECT	0 79.38 0.134 79.74 ;
		RECT	0 79.956 0.134 80.601 ;
		RECT	0 80.817 0.134 81.084 ;
		RECT	0 81.3 0.134 82.176 ;
		RECT	201.531 0 201.665 82.176 ;
		RECT	0.134 0 201.531 0.206 ;
		RECT	0.134 81.97 201.531 82.176 ;
		LAYER	V1 DESIGNRULEWIDTH 0 ;
		RECT	0 0 201.665 82.176 ;
		LAYER	V2 DESIGNRULEWIDTH 0 ;
		RECT	0 0 201.665 82.176 ;
	END

END gf12lp_1rw_lg12_w32_bit

END LIBRARY

