##
## LEF for PtnCells ;
## created by Innovus v18.10-p002_1 on Mon Oct 26 17:19:57 2020
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO temp_hd_inv8_header3
  CLASS BLOCK ;
  SIZE 100.280000 BY 100.300000 ;
  FOREIGN temp_hd_inv8_header3 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK_REF
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.637 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.8956 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.384 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 25.841 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 127.983 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.160000 99.815000 0.300000 100.300000 ;
    END
  END CLK_REF
  PIN RESET_COUNTERn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.4281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 117.975 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 11.844 LAYER met2  ;
    ANTENNAMAXAREACAR 13.7206 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 60.5698 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 9.820000 99.815000 9.960000 100.300000 ;
    END
  END RESET_COUNTERn
  PIN SEL_CONV_TIME[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4231 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8895 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 7.23293 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.2747 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.162222 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 30.060000 99.815000 30.200000 100.300000 ;
    END
  END SEL_CONV_TIME[3]
  PIN SEL_CONV_TIME[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.604 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.8328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.912 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met3  ;
    ANTENNAMAXAREACAR 12.0329 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 58.0975 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.248081 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 39.720000 99.815000 39.860000 100.300000 ;
    END
  END SEL_CONV_TIME[2]
  PIN SEL_CONV_TIME[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3375 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.3535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 6.3401 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.6588 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 49.840000 99.815000 49.980000 100.300000 ;
    END
  END SEL_CONV_TIME[1]
  PIN SEL_CONV_TIME[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7299 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.5415 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.81 LAYER met2  ;
    ANTENNAMAXAREACAR 6.06024 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.5974 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.144545 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 59.960000 99.815000 60.100000 100.300000 ;
    END
  END SEL_CONV_TIME[0]
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.765 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.664 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.9028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.952 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 69.6681 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 356.226 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 69.620000 99.815000 69.760000 100.300000 ;
    END
  END en
  PIN DOUT[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1583 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.6835 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.980000 0.000000 100.120000 0.485000 ;
    END
  END DOUT[23]
  PIN DOUT[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0159 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.9715 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 95.840000 0.000000 95.980000 0.485000 ;
    END
  END DOUT[22]
  PIN DOUT[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8283 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0335 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 91.700000 0.000000 91.840000 0.485000 ;
    END
  END DOUT[21]
  PIN DOUT[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0675 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 87.100000 0.000000 87.240000 0.485000 ;
    END
  END DOUT[20]
  PIN DOUT[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0675 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 82.960000 0.000000 83.100000 0.485000 ;
    END
  END DOUT[19]
  PIN DOUT[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0675 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 78.360000 0.000000 78.500000 0.485000 ;
    END
  END DOUT[18]
  PIN DOUT[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0675 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 74.220000 0.000000 74.360000 0.485000 ;
    END
  END DOUT[17]
  PIN DOUT[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0675 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 69.620000 0.000000 69.760000 0.485000 ;
    END
  END DOUT[16]
  PIN DOUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0675 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 65.480000 0.000000 65.620000 0.485000 ;
    END
  END DOUT[15]
  PIN DOUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0675 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 61.340000 0.000000 61.480000 0.485000 ;
    END
  END DOUT[14]
  PIN DOUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0159 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.9715 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 56.740000 0.000000 56.880000 0.485000 ;
    END
  END DOUT[13]
  PIN DOUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0159 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.9715 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 52.600000 0.000000 52.740000 0.485000 ;
    END
  END DOUT[12]
  PIN DOUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0675 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 48.000000 0.000000 48.140000 0.485000 ;
    END
  END DOUT[11]
  PIN DOUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0159 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.9715 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 43.860000 0.000000 44.000000 0.485000 ;
    END
  END DOUT[10]
  PIN DOUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1111 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4475 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 39.260000 0.000000 39.400000 0.485000 ;
    END
  END DOUT[9]
  PIN DOUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5391 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.5875 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 35.120000 0.000000 35.260000 0.485000 ;
    END
  END DOUT[8]
  PIN DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.2747 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.2655 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 30.980000 0.000000 31.120000 0.485000 ;
    END
  END DOUT[7]
  PIN DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.0815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.2995 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 26.380000 0.000000 26.520000 0.485000 ;
    END
  END DOUT[6]
  PIN DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.8239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.0115 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 22.240000 0.000000 22.380000 0.485000 ;
    END
  END DOUT[5]
  PIN DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.8239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.0115 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 17.640000 0.000000 17.780000 0.485000 ;
    END
  END DOUT[4]
  PIN DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3391 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.5875 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 13.500000 0.000000 13.640000 0.485000 ;
    END
  END DOUT[3]
  PIN DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3335 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.5595 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 8.900000 0.000000 9.040000 0.485000 ;
    END
  END DOUT[2]
  PIN DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.0935 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.2415 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 4.760000 0.000000 4.900000 0.485000 ;
    END
  END DOUT[1]
  PIN DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4355 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.4903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.3435 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.160000 0.000000 0.300000 0.485000 ;
    END
  END DOUT[0]
  PIN DONE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0742 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.21 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.517 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.4648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.315 LAYER met3  ;
    ANTENNAMAXAREACAR 16.9838 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 85.0254 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.290159 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 79.740000 99.815000 79.880000 100.300000 ;
    END
  END DONE
  PIN out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5904 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.791 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.9548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.896 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 89.860000 99.815000 90.000000 100.300000 ;
    END
  END out
  PIN outb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4654 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.166 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.0087 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.512 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 99.520000 99.815000 99.660000 100.300000 ;
    END
  END outb
  PIN lc_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5303 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.4355 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 26.0869 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 120.274 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 19.940000 99.815000 20.080000 100.300000 ;
    END
  END lc_out
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 98.680000 8.020000 100.280000 9.620000 ;
    END
    PORT
      LAYER met4 ;
        RECT 90.840000 98.700000 92.440000 100.300000 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.840000 98.700000 9.440000 100.300000 ;
    END
    PORT
      LAYER met5 ;
        RECT 98.680000 88.980000 100.280000 90.580000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 88.980000 1.600000 90.580000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 8.020000 1.600000 9.620000 ;
    END
    PORT
      LAYER met4 ;
        RECT 90.840000 0.000000 92.440000 1.600000 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.840000 0.000000 9.440000 1.600000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 90.840000 0.000000 92.440000 100.300000 ;
        RECT 7.840000 0.000000 9.440000 100.300000 ;
      LAYER met5 ;
        RECT 0.000000 8.020000 100.280000 9.620000 ;
        RECT 0.000000 88.980000 100.280000 90.580000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 98.680000 4.820000 100.280000 6.420000 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.040000 98.700000 95.640000 100.300000 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.640000 98.700000 6.240000 100.300000 ;
    END
    PORT
      LAYER met5 ;
        RECT 98.680000 92.180000 100.280000 93.780000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 92.180000 1.600000 93.780000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 4.820000 1.600000 6.420000 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.040000 0.000000 95.640000 1.600000 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.640000 0.000000 6.240000 1.600000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 94.040000 0.000000 95.640000 100.300000 ;
        RECT 4.640000 0.000000 6.240000 100.300000 ;
      LAYER met5 ;
        RECT 0.000000 4.820000 100.280000 6.420000 ;
        RECT 0.000000 92.180000 100.280000 93.780000 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 100.280000 100.300000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 100.280000 100.300000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 100.280000 100.300000 ;
    LAYER met3 ;
      RECT 0.000000 0.000000 100.280000 100.300000 ;
    LAYER met4 ;
      RECT 0.000000 0.000000 100.280000 100.300000 ;
    LAYER met5 ;
      RECT 0.000000 0.000000 100.280000 100.300000 ;
  END
END temp_hd_inv8_header3

END LIBRARY
